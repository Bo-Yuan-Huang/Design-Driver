
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [6:0] \oc8051_golden_model_1.n0988 ;
  wire \oc8051_golden_model_1.n0989 ;
  wire \oc8051_golden_model_1.n0990 ;
  wire \oc8051_golden_model_1.n0991 ;
  wire \oc8051_golden_model_1.n0992 ;
  wire \oc8051_golden_model_1.n0993 ;
  wire \oc8051_golden_model_1.n0994 ;
  wire \oc8051_golden_model_1.n0995 ;
  wire \oc8051_golden_model_1.n0996 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire [7:0] \oc8051_golden_model_1.n1004 ;
  wire [7:0] \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire \oc8051_golden_model_1.n1018 ;
  wire \oc8051_golden_model_1.n1019 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire [7:0] \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1043 ;
  wire [7:0] \oc8051_golden_model_1.n1044 ;
  wire [3:0] \oc8051_golden_model_1.n1137 ;
  wire [3:0] \oc8051_golden_model_1.n1139 ;
  wire [3:0] \oc8051_golden_model_1.n1141 ;
  wire [3:0] \oc8051_golden_model_1.n1142 ;
  wire [3:0] \oc8051_golden_model_1.n1143 ;
  wire [3:0] \oc8051_golden_model_1.n1144 ;
  wire [3:0] \oc8051_golden_model_1.n1145 ;
  wire [3:0] \oc8051_golden_model_1.n1146 ;
  wire [3:0] \oc8051_golden_model_1.n1147 ;
  wire \oc8051_golden_model_1.n1194 ;
  wire \oc8051_golden_model_1.n1239 ;
  wire [8:0] \oc8051_golden_model_1.n1240 ;
  wire [8:0] \oc8051_golden_model_1.n1241 ;
  wire [7:0] \oc8051_golden_model_1.n1242 ;
  wire \oc8051_golden_model_1.n1243 ;
  wire [2:0] \oc8051_golden_model_1.n1244 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [1:0] \oc8051_golden_model_1.n1246 ;
  wire [7:0] \oc8051_golden_model_1.n1247 ;
  wire [6:0] \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1251 ;
  wire \oc8051_golden_model_1.n1252 ;
  wire \oc8051_golden_model_1.n1253 ;
  wire \oc8051_golden_model_1.n1254 ;
  wire \oc8051_golden_model_1.n1255 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [7:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1280 ;
  wire [7:0] \oc8051_golden_model_1.n1281 ;
  wire [15:0] \oc8051_golden_model_1.n1323 ;
  wire [7:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1328 ;
  wire \oc8051_golden_model_1.n1329 ;
  wire \oc8051_golden_model_1.n1330 ;
  wire \oc8051_golden_model_1.n1331 ;
  wire \oc8051_golden_model_1.n1332 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire \oc8051_golden_model_1.n1340 ;
  wire [7:0] \oc8051_golden_model_1.n1341 ;
  wire [8:0] \oc8051_golden_model_1.n1343 ;
  wire [8:0] \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire [3:0] \oc8051_golden_model_1.n1349 ;
  wire [4:0] \oc8051_golden_model_1.n1350 ;
  wire [4:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [8:0] \oc8051_golden_model_1.n1356 ;
  wire \oc8051_golden_model_1.n1364 ;
  wire [7:0] \oc8051_golden_model_1.n1365 ;
  wire [6:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1381 ;
  wire [7:0] \oc8051_golden_model_1.n1382 ;
  wire [8:0] \oc8051_golden_model_1.n1404 ;
  wire \oc8051_golden_model_1.n1405 ;
  wire [4:0] \oc8051_golden_model_1.n1410 ;
  wire \oc8051_golden_model_1.n1411 ;
  wire \oc8051_golden_model_1.n1419 ;
  wire [7:0] \oc8051_golden_model_1.n1420 ;
  wire [6:0] \oc8051_golden_model_1.n1421 ;
  wire \oc8051_golden_model_1.n1436 ;
  wire [7:0] \oc8051_golden_model_1.n1437 ;
  wire [8:0] \oc8051_golden_model_1.n1439 ;
  wire [8:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1442 ;
  wire [3:0] \oc8051_golden_model_1.n1443 ;
  wire [4:0] \oc8051_golden_model_1.n1444 ;
  wire [4:0] \oc8051_golden_model_1.n1446 ;
  wire \oc8051_golden_model_1.n1447 ;
  wire [8:0] \oc8051_golden_model_1.n1448 ;
  wire \oc8051_golden_model_1.n1455 ;
  wire [7:0] \oc8051_golden_model_1.n1456 ;
  wire [6:0] \oc8051_golden_model_1.n1457 ;
  wire \oc8051_golden_model_1.n1472 ;
  wire [7:0] \oc8051_golden_model_1.n1473 ;
  wire [8:0] \oc8051_golden_model_1.n1476 ;
  wire \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1484 ;
  wire [7:0] \oc8051_golden_model_1.n1485 ;
  wire [6:0] \oc8051_golden_model_1.n1486 ;
  wire [7:0] \oc8051_golden_model_1.n1487 ;
  wire [8:0] \oc8051_golden_model_1.n1489 ;
  wire [8:0] \oc8051_golden_model_1.n1491 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [4:0] \oc8051_golden_model_1.n1493 ;
  wire [4:0] \oc8051_golden_model_1.n1495 ;
  wire \oc8051_golden_model_1.n1496 ;
  wire [8:0] \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire [4:0] \oc8051_golden_model_1.n1524 ;
  wire \oc8051_golden_model_1.n1525 ;
  wire [7:0] \oc8051_golden_model_1.n1526 ;
  wire [6:0] \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [8:0] \oc8051_golden_model_1.n1530 ;
  wire \oc8051_golden_model_1.n1531 ;
  wire \oc8051_golden_model_1.n1538 ;
  wire [7:0] \oc8051_golden_model_1.n1539 ;
  wire [6:0] \oc8051_golden_model_1.n1540 ;
  wire [7:0] \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [6:0] \oc8051_golden_model_1.n1543 ;
  wire [7:0] \oc8051_golden_model_1.n1544 ;
  wire [8:0] \oc8051_golden_model_1.n1547 ;
  wire [8:0] \oc8051_golden_model_1.n1548 ;
  wire [7:0] \oc8051_golden_model_1.n1549 ;
  wire [7:0] \oc8051_golden_model_1.n1550 ;
  wire [6:0] \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1552 ;
  wire \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire \oc8051_golden_model_1.n1555 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1559 ;
  wire \oc8051_golden_model_1.n1566 ;
  wire [7:0] \oc8051_golden_model_1.n1567 ;
  wire [7:0] \oc8051_golden_model_1.n1568 ;
  wire [8:0] \oc8051_golden_model_1.n1571 ;
  wire [8:0] \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire [4:0] \oc8051_golden_model_1.n1575 ;
  wire [4:0] \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1585 ;
  wire [7:0] \oc8051_golden_model_1.n1586 ;
  wire [6:0] \oc8051_golden_model_1.n1587 ;
  wire \oc8051_golden_model_1.n1602 ;
  wire [7:0] \oc8051_golden_model_1.n1603 ;
  wire [8:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1608 ;
  wire [4:0] \oc8051_golden_model_1.n1610 ;
  wire \oc8051_golden_model_1.n1611 ;
  wire \oc8051_golden_model_1.n1618 ;
  wire [7:0] \oc8051_golden_model_1.n1619 ;
  wire [6:0] \oc8051_golden_model_1.n1620 ;
  wire \oc8051_golden_model_1.n1635 ;
  wire [7:0] \oc8051_golden_model_1.n1636 ;
  wire [8:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1641 ;
  wire [4:0] \oc8051_golden_model_1.n1643 ;
  wire \oc8051_golden_model_1.n1644 ;
  wire \oc8051_golden_model_1.n1651 ;
  wire [7:0] \oc8051_golden_model_1.n1652 ;
  wire [6:0] \oc8051_golden_model_1.n1653 ;
  wire \oc8051_golden_model_1.n1668 ;
  wire [7:0] \oc8051_golden_model_1.n1669 ;
  wire [8:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1674 ;
  wire [4:0] \oc8051_golden_model_1.n1676 ;
  wire \oc8051_golden_model_1.n1677 ;
  wire \oc8051_golden_model_1.n1684 ;
  wire [7:0] \oc8051_golden_model_1.n1685 ;
  wire [6:0] \oc8051_golden_model_1.n1686 ;
  wire \oc8051_golden_model_1.n1701 ;
  wire [7:0] \oc8051_golden_model_1.n1702 ;
  wire [7:0] \oc8051_golden_model_1.n1727 ;
  wire [6:0] \oc8051_golden_model_1.n1728 ;
  wire [7:0] \oc8051_golden_model_1.n1729 ;
  wire \oc8051_golden_model_1.n1784 ;
  wire [7:0] \oc8051_golden_model_1.n1785 ;
  wire \oc8051_golden_model_1.n1801 ;
  wire [7:0] \oc8051_golden_model_1.n1802 ;
  wire \oc8051_golden_model_1.n1818 ;
  wire [7:0] \oc8051_golden_model_1.n1819 ;
  wire \oc8051_golden_model_1.n1835 ;
  wire [7:0] \oc8051_golden_model_1.n1836 ;
  wire [7:0] \oc8051_golden_model_1.n1859 ;
  wire [6:0] \oc8051_golden_model_1.n1860 ;
  wire [7:0] \oc8051_golden_model_1.n1861 ;
  wire \oc8051_golden_model_1.n1916 ;
  wire [7:0] \oc8051_golden_model_1.n1917 ;
  wire \oc8051_golden_model_1.n1933 ;
  wire [7:0] \oc8051_golden_model_1.n1934 ;
  wire \oc8051_golden_model_1.n1950 ;
  wire [7:0] \oc8051_golden_model_1.n1951 ;
  wire \oc8051_golden_model_1.n1967 ;
  wire [7:0] \oc8051_golden_model_1.n1968 ;
  wire \oc8051_golden_model_1.n2065 ;
  wire [7:0] \oc8051_golden_model_1.n2066 ;
  wire \oc8051_golden_model_1.n2082 ;
  wire [7:0] \oc8051_golden_model_1.n2083 ;
  wire \oc8051_golden_model_1.n2099 ;
  wire [7:0] \oc8051_golden_model_1.n2100 ;
  wire \oc8051_golden_model_1.n2116 ;
  wire [7:0] \oc8051_golden_model_1.n2117 ;
  wire \oc8051_golden_model_1.n2121 ;
  wire [6:0] \oc8051_golden_model_1.n2122 ;
  wire [7:0] \oc8051_golden_model_1.n2123 ;
  wire [6:0] \oc8051_golden_model_1.n2124 ;
  wire [7:0] \oc8051_golden_model_1.n2125 ;
  wire \oc8051_golden_model_1.n2140 ;
  wire [7:0] \oc8051_golden_model_1.n2141 ;
  wire \oc8051_golden_model_1.n2180 ;
  wire [7:0] \oc8051_golden_model_1.n2181 ;
  wire [6:0] \oc8051_golden_model_1.n2182 ;
  wire [7:0] \oc8051_golden_model_1.n2183 ;
  wire [3:0] \oc8051_golden_model_1.n2190 ;
  wire \oc8051_golden_model_1.n2191 ;
  wire [7:0] \oc8051_golden_model_1.n2192 ;
  wire [6:0] \oc8051_golden_model_1.n2193 ;
  wire \oc8051_golden_model_1.n2208 ;
  wire [7:0] \oc8051_golden_model_1.n2209 ;
  wire [7:0] \oc8051_golden_model_1.n2421 ;
  wire \oc8051_golden_model_1.n2424 ;
  wire \oc8051_golden_model_1.n2426 ;
  wire \oc8051_golden_model_1.n2432 ;
  wire [7:0] \oc8051_golden_model_1.n2433 ;
  wire [6:0] \oc8051_golden_model_1.n2434 ;
  wire \oc8051_golden_model_1.n2449 ;
  wire [7:0] \oc8051_golden_model_1.n2450 ;
  wire \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2456 ;
  wire \oc8051_golden_model_1.n2462 ;
  wire [7:0] \oc8051_golden_model_1.n2463 ;
  wire [6:0] \oc8051_golden_model_1.n2464 ;
  wire \oc8051_golden_model_1.n2479 ;
  wire [7:0] \oc8051_golden_model_1.n2480 ;
  wire \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2486 ;
  wire \oc8051_golden_model_1.n2492 ;
  wire [7:0] \oc8051_golden_model_1.n2493 ;
  wire [6:0] \oc8051_golden_model_1.n2494 ;
  wire \oc8051_golden_model_1.n2509 ;
  wire [7:0] \oc8051_golden_model_1.n2510 ;
  wire \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2516 ;
  wire \oc8051_golden_model_1.n2522 ;
  wire [7:0] \oc8051_golden_model_1.n2523 ;
  wire [6:0] \oc8051_golden_model_1.n2524 ;
  wire \oc8051_golden_model_1.n2539 ;
  wire [7:0] \oc8051_golden_model_1.n2540 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire [7:0] \oc8051_golden_model_1.n2545 ;
  wire [7:0] \oc8051_golden_model_1.n2546 ;
  wire [6:0] \oc8051_golden_model_1.n2547 ;
  wire [7:0] \oc8051_golden_model_1.n2548 ;
  wire [15:0] \oc8051_golden_model_1.n2552 ;
  wire \oc8051_golden_model_1.n2558 ;
  wire [7:0] \oc8051_golden_model_1.n2559 ;
  wire [6:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2575 ;
  wire [7:0] \oc8051_golden_model_1.n2576 ;
  wire \oc8051_golden_model_1.n2579 ;
  wire [7:0] \oc8051_golden_model_1.n2580 ;
  wire [6:0] \oc8051_golden_model_1.n2581 ;
  wire [7:0] \oc8051_golden_model_1.n2582 ;
  wire \oc8051_golden_model_1.n2614 ;
  wire [7:0] \oc8051_golden_model_1.n2615 ;
  wire [6:0] \oc8051_golden_model_1.n2616 ;
  wire [7:0] \oc8051_golden_model_1.n2617 ;
  wire \oc8051_golden_model_1.n2622 ;
  wire [7:0] \oc8051_golden_model_1.n2623 ;
  wire [6:0] \oc8051_golden_model_1.n2624 ;
  wire [7:0] \oc8051_golden_model_1.n2625 ;
  wire \oc8051_golden_model_1.n2630 ;
  wire [7:0] \oc8051_golden_model_1.n2631 ;
  wire [6:0] \oc8051_golden_model_1.n2632 ;
  wire [7:0] \oc8051_golden_model_1.n2633 ;
  wire \oc8051_golden_model_1.n2638 ;
  wire [7:0] \oc8051_golden_model_1.n2639 ;
  wire [6:0] \oc8051_golden_model_1.n2640 ;
  wire [7:0] \oc8051_golden_model_1.n2641 ;
  wire \oc8051_golden_model_1.n2646 ;
  wire [7:0] \oc8051_golden_model_1.n2647 ;
  wire [6:0] \oc8051_golden_model_1.n2648 ;
  wire [7:0] \oc8051_golden_model_1.n2649 ;
  wire [7:0] \oc8051_golden_model_1.n2674 ;
  wire [6:0] \oc8051_golden_model_1.n2675 ;
  wire [7:0] \oc8051_golden_model_1.n2676 ;
  wire [3:0] \oc8051_golden_model_1.n2677 ;
  wire [7:0] \oc8051_golden_model_1.n2678 ;
  wire \oc8051_golden_model_1.n2679 ;
  wire \oc8051_golden_model_1.n2680 ;
  wire \oc8051_golden_model_1.n2681 ;
  wire \oc8051_golden_model_1.n2682 ;
  wire \oc8051_golden_model_1.n2683 ;
  wire \oc8051_golden_model_1.n2684 ;
  wire \oc8051_golden_model_1.n2685 ;
  wire \oc8051_golden_model_1.n2686 ;
  wire \oc8051_golden_model_1.n2693 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [6:0] \oc8051_golden_model_1.n2715 ;
  wire [7:0] \oc8051_golden_model_1.n2731 ;
  wire \oc8051_golden_model_1.n2732 ;
  wire \oc8051_golden_model_1.n2733 ;
  wire \oc8051_golden_model_1.n2734 ;
  wire \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2736 ;
  wire \oc8051_golden_model_1.n2737 ;
  wire \oc8051_golden_model_1.n2738 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire \oc8051_golden_model_1.n2746 ;
  wire [7:0] \oc8051_golden_model_1.n2747 ;
  wire \oc8051_golden_model_1.n2748 ;
  wire \oc8051_golden_model_1.n2749 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2762 ;
  wire [7:0] \oc8051_golden_model_1.n2763 ;
  wire [7:0] \oc8051_golden_model_1.n2795 ;
  wire [6:0] \oc8051_golden_model_1.n2796 ;
  wire [7:0] \oc8051_golden_model_1.n2797 ;
  wire \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire [6:0] \oc8051_golden_model_1.n2818 ;
  wire \oc8051_golden_model_1.n2833 ;
  wire [7:0] \oc8051_golden_model_1.n2834 ;
  wire [7:0] \oc8051_golden_model_1.n2838 ;
  wire [3:0] \oc8051_golden_model_1.n2839 ;
  wire [7:0] \oc8051_golden_model_1.n2840 ;
  wire \oc8051_golden_model_1.n2841 ;
  wire \oc8051_golden_model_1.n2842 ;
  wire \oc8051_golden_model_1.n2843 ;
  wire \oc8051_golden_model_1.n2844 ;
  wire \oc8051_golden_model_1.n2845 ;
  wire \oc8051_golden_model_1.n2846 ;
  wire \oc8051_golden_model_1.n2847 ;
  wire \oc8051_golden_model_1.n2848 ;
  wire \oc8051_golden_model_1.n2855 ;
  wire [7:0] \oc8051_golden_model_1.n2856 ;
  wire \oc8051_golden_model_1.n2874 ;
  wire [7:0] \oc8051_golden_model_1.n2875 ;
  wire \oc8051_golden_model_1.n2891 ;
  wire [7:0] \oc8051_golden_model_1.n2892 ;
  wire [7:0] \oc8051_golden_model_1.n2893 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  wire property_invalid_psw_1_r;
  output property_invalid_sp;
  wire property_invalid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not _44061_ (_41806_, rst);
  not _44062_ (_15625_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _44063_ (_15636_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _44064_ (_15647_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15636_);
  and _44065_ (_15658_, _15647_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44066_ (_15669_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15636_);
  and _44067_ (_15680_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _15636_);
  nor _44068_ (_15691_, _15680_, _15669_);
  and _44069_ (_15702_, _15691_, _15658_);
  nor _44070_ (_15713_, _15702_, _15625_);
  and _44071_ (_15724_, _15625_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44072_ (_15735_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _44073_ (_15746_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _15735_);
  nor _44074_ (_15757_, _15746_, _15724_);
  not _44075_ (_15768_, _15757_);
  and _44076_ (_15779_, _15768_, _15702_);
  or _44077_ (_15790_, _15779_, _15713_);
  and _44078_ (_22434_, _15790_, _41806_);
  nor _44079_ (_15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44080_ (_15821_, _15810_);
  and _44081_ (_15832_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _44082_ (_15843_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _44083_ (_15854_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _44084_ (_15865_, _15854_);
  not _44085_ (_15876_, _15746_);
  nor _44086_ (_15887_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _44087_ (_15898_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _44088_ (_15909_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _15898_);
  nor _44089_ (_15920_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not _44090_ (_15931_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor _44091_ (_15942_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _15931_);
  nor _44092_ (_15953_, _15942_, _15920_);
  nor _44093_ (_15964_, _15953_, _15909_);
  not _44094_ (_15975_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _44095_ (_15986_, _15909_, _15975_);
  nor _44096_ (_15997_, _15986_, _15964_);
  and _44097_ (_16008_, _15997_, _15887_);
  not _44098_ (_16019_, _16008_);
  and _44099_ (_16030_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44100_ (_16041_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _44101_ (_16052_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44102_ (_16063_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _16052_);
  and _44103_ (_16074_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _44104_ (_16085_, _16074_, _16041_);
  and _44105_ (_16096_, _16085_, _16019_);
  nor _44106_ (_16107_, _16096_, _15876_);
  not _44107_ (_16118_, _15724_);
  nor _44108_ (_16128_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor _44109_ (_16139_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _15931_);
  nor _44110_ (_16150_, _16139_, _16128_);
  nor _44111_ (_16161_, _16150_, _15909_);
  not _44112_ (_16172_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _44113_ (_16183_, _15909_, _16172_);
  nor _44114_ (_16194_, _16183_, _16161_);
  and _44115_ (_16205_, _16194_, _15887_);
  not _44116_ (_16216_, _16205_);
  and _44117_ (_16227_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _44118_ (_16238_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _44119_ (_16249_, _16238_, _16227_);
  and _44120_ (_16260_, _16249_, _16216_);
  nor _44121_ (_16271_, _16260_, _16118_);
  nor _44122_ (_16282_, _16271_, _16107_);
  nor _44123_ (_16293_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor _44124_ (_16304_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _15931_);
  nor _44125_ (_16315_, _16304_, _16293_);
  nor _44126_ (_16326_, _16315_, _15909_);
  not _44127_ (_16337_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _44128_ (_16348_, _15909_, _16337_);
  nor _44129_ (_16359_, _16348_, _16326_);
  and _44130_ (_16370_, _16359_, _15887_);
  not _44131_ (_16381_, _16370_);
  and _44132_ (_16392_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _44133_ (_16403_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _44134_ (_16414_, _16403_, _16392_);
  and _44135_ (_16425_, _16414_, _16381_);
  nor _44136_ (_16436_, _16425_, _15768_);
  nor _44137_ (_16446_, _16436_, _15810_);
  and _44138_ (_16457_, _16446_, _16282_);
  nor _44139_ (_16468_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor _44140_ (_16479_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _15931_);
  nor _44141_ (_16490_, _16479_, _16468_);
  nor _44142_ (_16501_, _16490_, _15909_);
  not _44143_ (_16512_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _44144_ (_16523_, _15909_, _16512_);
  nor _44145_ (_16534_, _16523_, _16501_);
  and _44146_ (_16556_, _16534_, _15887_);
  not _44147_ (_16557_, _16556_);
  and _44148_ (_16568_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _44149_ (_16579_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _44150_ (_16590_, _16579_, _16568_);
  and _44151_ (_16601_, _16590_, _16557_);
  and _44152_ (_16612_, _16601_, _15810_);
  nor _44153_ (_16623_, _16612_, _16457_);
  not _44154_ (_16634_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44155_ (_16645_, _16634_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44156_ (_16656_, _16645_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44157_ (_16667_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _44158_ (_16678_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44159_ (_16689_, _16678_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44160_ (_16700_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _44161_ (_16711_, _16700_, _16667_);
  nor _44162_ (_16722_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44163_ (_16733_, _16722_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44164_ (_16744_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _44165_ (_16755_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44166_ (_16766_, _16645_, _16755_);
  and _44167_ (_16776_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _44168_ (_16787_, _16776_, _16744_);
  and _44169_ (_16798_, _16787_, _16711_);
  and _44170_ (_16809_, _16722_, _16634_);
  and _44171_ (_16820_, _16809_, _16534_);
  and _44172_ (_16831_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44173_ (_16842_, _16831_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44174_ (_16853_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _44175_ (_16864_, _16831_, _16755_);
  and _44176_ (_16875_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _44177_ (_16886_, _16875_, _16853_);
  not _44178_ (_16897_, _16886_);
  nor _44179_ (_16908_, _16897_, _16820_);
  and _44180_ (_16919_, _16908_, _16798_);
  not _44181_ (_16930_, _16919_);
  and _44182_ (_16941_, _16930_, _16623_);
  not _44183_ (_16952_, _16941_);
  nor _44184_ (_16963_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor _44185_ (_16974_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _15931_);
  nor _44186_ (_16985_, _16974_, _16963_);
  nor _44187_ (_16996_, _16985_, _15909_);
  not _44188_ (_17007_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _44189_ (_17018_, _15909_, _17007_);
  nor _44190_ (_17029_, _17018_, _16996_);
  and _44191_ (_17040_, _17029_, _15887_);
  not _44192_ (_17051_, _17040_);
  and _44193_ (_17062_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _44194_ (_17073_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _44195_ (_17084_, _17073_, _17062_);
  and _44196_ (_17094_, _17084_, _17051_);
  nor _44197_ (_17105_, _17094_, _15876_);
  nor _44198_ (_17116_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor _44199_ (_17127_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _15931_);
  nor _44200_ (_17138_, _17127_, _17116_);
  nor _44201_ (_17149_, _17138_, _15909_);
  not _44202_ (_17160_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _44203_ (_17171_, _15909_, _17160_);
  nor _44204_ (_17181_, _17171_, _17149_);
  and _44205_ (_17192_, _17181_, _15887_);
  not _44206_ (_17203_, _17192_);
  and _44207_ (_17214_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _44208_ (_17225_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44209_ (_17236_, _17225_, _17214_);
  and _44210_ (_17247_, _17236_, _17203_);
  nor _44211_ (_17258_, _17247_, _16118_);
  nor _44212_ (_17278_, _17258_, _17105_);
  nor _44213_ (_17279_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor _44214_ (_17300_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _15931_);
  nor _44215_ (_17301_, _17300_, _17279_);
  nor _44216_ (_17312_, _17301_, _15909_);
  not _44217_ (_17323_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _44218_ (_17334_, _15909_, _17323_);
  nor _44219_ (_17345_, _17334_, _17312_);
  and _44220_ (_17356_, _17345_, _15887_);
  not _44221_ (_17366_, _17356_);
  and _44222_ (_17377_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _44223_ (_17388_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44224_ (_17399_, _17388_, _17377_);
  and _44225_ (_17410_, _17399_, _17366_);
  nor _44226_ (_17421_, _17410_, _15768_);
  nor _44227_ (_17432_, _17421_, _15810_);
  and _44228_ (_17443_, _17432_, _17278_);
  nor _44229_ (_17454_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor _44230_ (_17464_, _15931_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor _44231_ (_17475_, _17464_, _17454_);
  nor _44232_ (_17486_, _17475_, _15909_);
  not _44233_ (_17497_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _44234_ (_17508_, _15909_, _17497_);
  nor _44235_ (_17519_, _17508_, _17486_);
  and _44236_ (_17530_, _17519_, _15887_);
  not _44237_ (_17541_, _17530_);
  and _44238_ (_17552_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _44239_ (_17562_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _44240_ (_17573_, _17562_, _17552_);
  and _44241_ (_17584_, _17573_, _17541_);
  and _44242_ (_17595_, _17584_, _15810_);
  or _44243_ (_17606_, _17595_, _17443_);
  and _44244_ (_17617_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _44245_ (_17628_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _44246_ (_17639_, _17628_, _17617_);
  and _44247_ (_17649_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _44248_ (_17660_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _44249_ (_17671_, _17660_, _17649_);
  and _44250_ (_17682_, _17671_, _17639_);
  and _44251_ (_17693_, _17519_, _16809_);
  and _44252_ (_17704_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _44253_ (_17715_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _44254_ (_17726_, _17715_, _17704_);
  not _44255_ (_17737_, _17726_);
  nor _44256_ (_17747_, _17737_, _17693_);
  and _44257_ (_17758_, _17747_, _17682_);
  nor _44258_ (_17769_, _17758_, _17606_);
  and _44259_ (_17780_, _17769_, _16952_);
  not _44260_ (_17791_, _17780_);
  and _44261_ (_17802_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _44262_ (_17813_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _44263_ (_17824_, _17813_, _17802_);
  and _44264_ (_17834_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _44265_ (_17845_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _44266_ (_17856_, _17845_, _17834_);
  and _44267_ (_17867_, _17856_, _17824_);
  and _44268_ (_17878_, _17181_, _16809_);
  and _44269_ (_17889_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _44270_ (_17900_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44271_ (_17911_, _17900_, _17889_);
  not _44272_ (_17922_, _17911_);
  nor _44273_ (_17932_, _17922_, _17878_);
  and _44274_ (_17943_, _17932_, _17867_);
  nor _44275_ (_17954_, _17943_, _17606_);
  and _44276_ (_17965_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _44277_ (_17976_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _44278_ (_17987_, _17976_, _17965_);
  and _44279_ (_17998_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _44280_ (_18009_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _44281_ (_18019_, _18009_, _17998_);
  and _44282_ (_18030_, _18019_, _17987_);
  and _44283_ (_18041_, _16809_, _16194_);
  and _44284_ (_18052_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _44285_ (_18063_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _44286_ (_18074_, _18063_, _18052_);
  not _44287_ (_18085_, _18074_);
  nor _44288_ (_18096_, _18085_, _18041_);
  and _44289_ (_18107_, _18096_, _18030_);
  not _44290_ (_18117_, _18107_);
  and _44291_ (_18128_, _18117_, _16623_);
  and _44292_ (_18139_, _17954_, _18128_);
  and _44293_ (_18150_, _16930_, _18139_);
  nor _44294_ (_18161_, _16941_, _18139_);
  nor _44295_ (_18172_, _18161_, _18150_);
  and _44296_ (_18183_, _18172_, _17954_);
  and _44297_ (_18194_, _17769_, _16941_);
  nor _44298_ (_18204_, _16919_, _17606_);
  not _44299_ (_18215_, _17758_);
  and _44300_ (_18226_, _18215_, _16623_);
  nor _44301_ (_18237_, _18226_, _18204_);
  nor _44302_ (_18248_, _18237_, _18194_);
  and _44303_ (_18259_, _18248_, _18183_);
  nor _44304_ (_18270_, _18248_, _18183_);
  nor _44305_ (_18281_, _18270_, _18259_);
  and _44306_ (_18292_, _18281_, _18150_);
  nor _44307_ (_18302_, _18292_, _18259_);
  nor _44308_ (_18313_, _18302_, _17791_);
  nor _44309_ (_18324_, _17606_, _18107_);
  and _44310_ (_18335_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _44311_ (_18346_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _44312_ (_18357_, _18346_, _18335_);
  and _44313_ (_18368_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _44314_ (_18379_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _44315_ (_18390_, _18379_, _18368_);
  and _44316_ (_18400_, _18390_, _18357_);
  and _44317_ (_18411_, _17029_, _16809_);
  and _44318_ (_18422_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _44319_ (_18433_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor _44320_ (_18444_, _18433_, _18422_);
  not _44321_ (_18455_, _18444_);
  nor _44322_ (_18466_, _18455_, _18411_);
  and _44323_ (_18477_, _18466_, _18400_);
  not _44324_ (_18488_, _18477_);
  and _44325_ (_18498_, _18488_, _16623_);
  and _44326_ (_18509_, _18498_, _18324_);
  not _44327_ (_18520_, _17943_);
  and _44328_ (_18531_, _18520_, _16623_);
  nor _44329_ (_18542_, _18531_, _18324_);
  nor _44330_ (_18553_, _18542_, _18139_);
  and _44331_ (_18564_, _18553_, _18509_);
  nor _44332_ (_18575_, _16941_, _17954_);
  nor _44333_ (_18586_, _18575_, _18183_);
  and _44334_ (_18597_, _18586_, _18564_);
  nor _44335_ (_18608_, _18281_, _18150_);
  nor _44336_ (_18618_, _18608_, _18292_);
  and _44337_ (_18629_, _18618_, _18597_);
  nor _44338_ (_18640_, _18618_, _18597_);
  nor _44339_ (_18651_, _18640_, _18629_);
  not _44340_ (_18662_, _18651_);
  and _44341_ (_18673_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _44342_ (_18684_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _44343_ (_18695_, _18684_, _18673_);
  and _44344_ (_18706_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _44345_ (_18717_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor _44346_ (_18727_, _18717_, _18706_);
  and _44347_ (_18738_, _18727_, _18695_);
  and _44348_ (_18749_, _17345_, _16809_);
  and _44349_ (_18760_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _44350_ (_18771_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44351_ (_18782_, _18771_, _18760_);
  not _44352_ (_18793_, _18782_);
  nor _44353_ (_18804_, _18793_, _18749_);
  and _44354_ (_18815_, _18804_, _18738_);
  nor _44355_ (_18826_, _18815_, _17606_);
  and _44356_ (_18837_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _44357_ (_18847_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _44358_ (_18858_, _18847_, _18837_);
  and _44359_ (_18869_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _44360_ (_18880_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor _44361_ (_18891_, _18880_, _18869_);
  and _44362_ (_18902_, _18891_, _18858_);
  and _44363_ (_18913_, _16809_, _15997_);
  and _44364_ (_18924_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _44365_ (_18935_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor _44366_ (_18946_, _18935_, _18924_);
  not _44367_ (_18957_, _18946_);
  nor _44368_ (_18967_, _18957_, _18913_);
  and _44369_ (_18978_, _18967_, _18902_);
  not _44370_ (_18989_, _18978_);
  and _44371_ (_19000_, _18989_, _16623_);
  and _44372_ (_19011_, _19000_, _18826_);
  not _44373_ (_19022_, _18815_);
  and _44374_ (_19033_, _19022_, _16623_);
  not _44375_ (_19044_, _19033_);
  nor _44376_ (_19055_, _18978_, _17606_);
  and _44377_ (_19066_, _19055_, _19044_);
  and _44378_ (_19076_, _19066_, _18498_);
  nor _44379_ (_19087_, _19076_, _19011_);
  nor _44380_ (_19098_, _18477_, _17606_);
  nor _44381_ (_19109_, _19098_, _18128_);
  nor _44382_ (_19120_, _19109_, _18509_);
  not _44383_ (_19131_, _19120_);
  nor _44384_ (_19142_, _19131_, _19087_);
  nor _44385_ (_19153_, _18553_, _18509_);
  nor _44386_ (_19164_, _19153_, _18564_);
  and _44387_ (_19175_, _19164_, _19142_);
  nor _44388_ (_19186_, _18586_, _18564_);
  nor _44389_ (_19196_, _19186_, _18597_);
  and _44390_ (_19207_, _19196_, _19175_);
  and _44391_ (_19218_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _44392_ (_19229_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _44393_ (_19240_, _19229_, _19218_);
  and _44394_ (_19251_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _44395_ (_19262_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _44396_ (_19273_, _19262_, _19251_);
  and _44397_ (_19284_, _19273_, _19240_);
  and _44398_ (_19294_, _16809_, _16359_);
  and _44399_ (_19305_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _44400_ (_19316_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor _44401_ (_19327_, _19316_, _19305_);
  not _44402_ (_19338_, _19327_);
  nor _44403_ (_19349_, _19338_, _19294_);
  and _44404_ (_19360_, _19349_, _19284_);
  nor _44405_ (_19371_, _19360_, _17606_);
  and _44406_ (_19382_, _19371_, _19033_);
  nor _44407_ (_19393_, _19000_, _18826_);
  nor _44408_ (_19404_, _19393_, _19011_);
  and _44409_ (_19414_, _19404_, _19382_);
  nor _44410_ (_19425_, _19066_, _18498_);
  nor _44411_ (_19436_, _19425_, _19076_);
  and _44412_ (_19447_, _19436_, _19414_);
  and _44413_ (_19458_, _19131_, _19087_);
  nor _44414_ (_19469_, _19458_, _19142_);
  and _44415_ (_19480_, _19469_, _19447_);
  nor _44416_ (_19491_, _19164_, _19142_);
  nor _44417_ (_19502_, _19491_, _19175_);
  and _44418_ (_19513_, _19502_, _19480_);
  nor _44419_ (_19523_, _19196_, _19175_);
  nor _44420_ (_19534_, _19523_, _19207_);
  and _44421_ (_19545_, _19534_, _19513_);
  nor _44422_ (_19556_, _19545_, _19207_);
  nor _44423_ (_19567_, _19556_, _18662_);
  nor _44424_ (_19578_, _19567_, _18629_);
  and _44425_ (_19589_, _18302_, _17791_);
  nor _44426_ (_19600_, _19589_, _18313_);
  not _44427_ (_19611_, _19600_);
  nor _44428_ (_19622_, _19611_, _19578_);
  or _44429_ (_19633_, _19622_, _18194_);
  nor _44430_ (_19643_, _19633_, _18313_);
  nor _44431_ (_19654_, _19643_, _15865_);
  and _44432_ (_19665_, _19643_, _15865_);
  nor _44433_ (_19676_, _19665_, _19654_);
  not _44434_ (_19687_, _19676_);
  and _44435_ (_19698_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _44436_ (_19709_, _19611_, _19578_);
  nor _44437_ (_19720_, _19709_, _19622_);
  and _44438_ (_19731_, _19720_, _19698_);
  and _44439_ (_19742_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and _44440_ (_19753_, _19556_, _18662_);
  nor _44441_ (_19763_, _19753_, _19567_);
  and _44442_ (_19774_, _19763_, _19742_);
  nor _44443_ (_19785_, _19763_, _19742_);
  nor _44444_ (_19796_, _19785_, _19774_);
  not _44445_ (_19807_, _19796_);
  and _44446_ (_19818_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor _44447_ (_19829_, _19534_, _19513_);
  nor _44448_ (_19840_, _19829_, _19545_);
  and _44449_ (_19851_, _19840_, _19818_);
  nor _44450_ (_19862_, _19840_, _19818_);
  nor _44451_ (_19872_, _19862_, _19851_);
  not _44452_ (_19883_, _19872_);
  and _44453_ (_19894_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor _44454_ (_19905_, _19502_, _19480_);
  nor _44455_ (_19916_, _19905_, _19513_);
  and _44456_ (_19927_, _19916_, _19894_);
  nor _44457_ (_19938_, _19916_, _19894_);
  nor _44458_ (_19949_, _19938_, _19927_);
  not _44459_ (_19960_, _19949_);
  and _44460_ (_19971_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor _44461_ (_19981_, _19469_, _19447_);
  nor _44462_ (_19992_, _19981_, _19480_);
  and _44463_ (_20003_, _19992_, _19971_);
  and _44464_ (_20014_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor _44465_ (_20025_, _19436_, _19414_);
  nor _44466_ (_20036_, _20025_, _19447_);
  and _44467_ (_20047_, _20036_, _20014_);
  and _44468_ (_20058_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor _44469_ (_20069_, _19404_, _19382_);
  nor _44470_ (_20080_, _20069_, _19414_);
  and _44471_ (_20091_, _20080_, _20058_);
  nor _44472_ (_20101_, _20036_, _20014_);
  nor _44473_ (_20112_, _20101_, _20047_);
  and _44474_ (_20123_, _20112_, _20091_);
  nor _44475_ (_20134_, _20123_, _20047_);
  not _44476_ (_20145_, _20134_);
  nor _44477_ (_20156_, _19992_, _19971_);
  nor _44478_ (_20167_, _20156_, _20003_);
  and _44479_ (_20178_, _20167_, _20145_);
  nor _44480_ (_20189_, _20178_, _20003_);
  nor _44481_ (_20200_, _20189_, _19960_);
  nor _44482_ (_20211_, _20200_, _19927_);
  nor _44483_ (_20222_, _20211_, _19883_);
  nor _44484_ (_20232_, _20222_, _19851_);
  nor _44485_ (_20243_, _20232_, _19807_);
  nor _44486_ (_20254_, _20243_, _19774_);
  nor _44487_ (_20265_, _19720_, _19698_);
  nor _44488_ (_20276_, _20265_, _19731_);
  not _44489_ (_20287_, _20276_);
  nor _44490_ (_20298_, _20287_, _20254_);
  nor _44491_ (_20309_, _20298_, _19731_);
  nor _44492_ (_20320_, _20309_, _19687_);
  nor _44493_ (_20331_, _20320_, _19654_);
  not _44494_ (_20342_, _20331_);
  and _44495_ (_20352_, _20342_, _15843_);
  and _44496_ (_20363_, _20352_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _44497_ (_20374_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _44498_ (_20385_, _20374_, _20363_);
  and _44499_ (_20396_, _20385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _44500_ (_20407_, _20396_, _15832_);
  and _44501_ (_20418_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _44502_ (_20429_, _20418_, _20407_);
  and _44503_ (_20440_, _20407_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _44504_ (_20451_, _20440_, _20429_);
  and _44505_ (_24620_, _20451_, _41806_);
  nor _44506_ (_20471_, _15702_, _15735_);
  and _44507_ (_20482_, _15702_, _15735_);
  or _44508_ (_20493_, _20482_, _20471_);
  and _44509_ (_02465_, _20493_, _41806_);
  not _44510_ (_20514_, _19360_);
  and _44511_ (_20525_, _20514_, _16623_);
  and _44512_ (_02660_, _20525_, _41806_);
  nor _44513_ (_20546_, _19371_, _19033_);
  nor _44514_ (_20557_, _20546_, _19382_);
  and _44515_ (_02854_, _20557_, _41806_);
  nor _44516_ (_20578_, _20080_, _20058_);
  nor _44517_ (_20589_, _20578_, _20091_);
  and _44518_ (_03057_, _20589_, _41806_);
  nor _44519_ (_20609_, _20112_, _20091_);
  nor _44520_ (_20620_, _20609_, _20123_);
  and _44521_ (_03268_, _20620_, _41806_);
  nor _44522_ (_20641_, _20167_, _20145_);
  nor _44523_ (_20652_, _20641_, _20178_);
  and _44524_ (_03469_, _20652_, _41806_);
  and _44525_ (_20673_, _20189_, _19960_);
  nor _44526_ (_20684_, _20673_, _20200_);
  and _44527_ (_03670_, _20684_, _41806_);
  and _44528_ (_20705_, _20211_, _19883_);
  nor _44529_ (_20715_, _20705_, _20222_);
  and _44530_ (_03871_, _20715_, _41806_);
  and _44531_ (_20736_, _20232_, _19807_);
  nor _44532_ (_20747_, _20736_, _20243_);
  and _44533_ (_04072_, _20747_, _41806_);
  and _44534_ (_20768_, _20287_, _20254_);
  nor _44535_ (_20779_, _20768_, _20298_);
  and _44536_ (_04173_, _20779_, _41806_);
  and _44537_ (_20800_, _20309_, _19687_);
  nor _44538_ (_20811_, _20800_, _20320_);
  and _44539_ (_04274_, _20811_, _41806_);
  nor _44540_ (_20832_, _20342_, _15843_);
  nor _44541_ (_20842_, _20832_, _20352_);
  and _44542_ (_04375_, _20842_, _41806_);
  and _44543_ (_20863_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor _44544_ (_20874_, _20863_, _20352_);
  nor _44545_ (_20885_, _20874_, _20363_);
  and _44546_ (_04476_, _20885_, _41806_);
  nor _44547_ (_20906_, _20374_, _20363_);
  nor _44548_ (_20917_, _20906_, _20385_);
  and _44549_ (_04577_, _20917_, _41806_);
  and _44550_ (_20937_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _44551_ (_20948_, _20937_, _20385_);
  nor _44552_ (_20959_, _20948_, _20396_);
  and _44553_ (_04678_, _20959_, _41806_);
  nor _44554_ (_20980_, _20396_, _15832_);
  nor _44555_ (_20991_, _20980_, _20407_);
  and _44556_ (_04779_, _20991_, _41806_);
  and _44557_ (_21012_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15636_);
  nor _44558_ (_21023_, _21012_, _15647_);
  not _44559_ (_21034_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _44560_ (_21044_, _15669_, _21034_);
  and _44561_ (_21055_, _21044_, _21023_);
  and _44562_ (_21066_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _44563_ (_21077_, _21066_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44564_ (_21088_, _21066_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44565_ (_21099_, _21088_, _21077_);
  and _44566_ (_00862_, _21099_, _41806_);
  and _44567_ (_00893_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _41806_);
  not _44568_ (_21130_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _44569_ (_21141_, _17410_, _21130_);
  and _44570_ (_21152_, _17094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44571_ (_21162_, _21152_, _21141_);
  nor _44572_ (_21173_, _21162_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44573_ (_21184_, _17247_, _21130_);
  and _44574_ (_21195_, _17584_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _44575_ (_21206_, _21195_, _21184_);
  and _44576_ (_21217_, _21206_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44577_ (_21228_, _21217_, _21173_);
  nor _44578_ (_21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _44579_ (_21250_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and _44580_ (_21261_, _21239_, _17758_);
  nor _44581_ (_21271_, _21261_, _21250_);
  not _44582_ (_21282_, _21271_);
  and _44583_ (_21293_, _16425_, _21130_);
  and _44584_ (_21304_, _16096_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44585_ (_21315_, _21304_, _21293_);
  nor _44586_ (_21326_, _21315_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44587_ (_21337_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44588_ (_21348_, _16260_, _21130_);
  and _44589_ (_21359_, _16601_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44590_ (_21370_, _21359_, _21348_);
  nor _44591_ (_21380_, _21370_, _21337_);
  nor _44592_ (_21391_, _21380_, _21326_);
  nor _44593_ (_21402_, _21391_, _21282_);
  and _44594_ (_21413_, _21391_, _21282_);
  nor _44595_ (_21424_, _21413_, _21402_);
  nor _44596_ (_21435_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and _44597_ (_21446_, _21239_, _16919_);
  nor _44598_ (_21457_, _21446_, _21435_);
  not _44599_ (_21468_, _21457_);
  nor _44600_ (_21489_, _17410_, _21130_);
  nor _44601_ (_21501_, _21489_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44602_ (_21513_, _17094_, _21130_);
  and _44603_ (_21525_, _17247_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44604_ (_21537_, _21525_, _21513_);
  nor _44605_ (_21549_, _21537_, _21337_);
  nor _44606_ (_21550_, _21549_, _21501_);
  nor _44607_ (_21561_, _21550_, _21468_);
  and _44608_ (_21572_, _21550_, _21468_);
  nor _44609_ (_21583_, _21572_, _21561_);
  not _44610_ (_21594_, _21583_);
  nor _44611_ (_21604_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and _44612_ (_21615_, _21239_, _17943_);
  nor _44613_ (_21626_, _21615_, _21604_);
  not _44614_ (_21637_, _21626_);
  nor _44615_ (_21648_, _16425_, _21130_);
  nor _44616_ (_21659_, _21648_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44617_ (_21670_, _16096_, _21130_);
  and _44618_ (_21681_, _16260_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44619_ (_21692_, _21681_, _21670_);
  nor _44620_ (_21703_, _21692_, _21337_);
  nor _44621_ (_21713_, _21703_, _21659_);
  nor _44622_ (_21724_, _21713_, _21637_);
  and _44623_ (_21735_, _21713_, _21637_);
  nor _44624_ (_21746_, _21735_, _21724_);
  not _44625_ (_21757_, _21746_);
  and _44626_ (_21768_, _21162_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44627_ (_21779_, _21768_);
  nor _44628_ (_21790_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and _44629_ (_21801_, _21239_, _18107_);
  nor _44630_ (_21812_, _21801_, _21790_);
  and _44631_ (_21822_, _21812_, _21779_);
  and _44632_ (_21833_, _21315_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44633_ (_21844_, _21833_);
  and _44634_ (_21855_, _21239_, _18477_);
  nor _44635_ (_21866_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor _44636_ (_21877_, _21866_, _21855_);
  and _44637_ (_21888_, _21877_, _21844_);
  nor _44638_ (_21899_, _21877_, _21844_);
  nor _44639_ (_21910_, _21899_, _21888_);
  not _44640_ (_21921_, _21910_);
  and _44641_ (_21931_, _21489_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44642_ (_21942_, _21931_);
  and _44643_ (_21953_, _21239_, _18978_);
  nor _44644_ (_21964_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor _44645_ (_21975_, _21964_, _21953_);
  and _44646_ (_21986_, _21975_, _21942_);
  and _44647_ (_21997_, _21648_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44648_ (_22008_, _21997_);
  nor _44649_ (_22019_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and _44650_ (_22030_, _21239_, _18815_);
  nor _44651_ (_22040_, _22030_, _22019_);
  nor _44652_ (_22061_, _22040_, _22008_);
  not _44653_ (_22062_, _22061_);
  nor _44654_ (_22073_, _21975_, _21942_);
  nor _44655_ (_22084_, _22073_, _21986_);
  and _44656_ (_22095_, _22084_, _22062_);
  nor _44657_ (_22106_, _22095_, _21986_);
  nor _44658_ (_22117_, _22106_, _21921_);
  nor _44659_ (_22128_, _22117_, _21888_);
  nor _44660_ (_22139_, _21812_, _21779_);
  nor _44661_ (_22150_, _22139_, _21822_);
  not _44662_ (_22160_, _22150_);
  nor _44663_ (_22171_, _22160_, _22128_);
  nor _44664_ (_22182_, _22171_, _21822_);
  nor _44665_ (_22193_, _22182_, _21757_);
  nor _44666_ (_22204_, _22193_, _21724_);
  nor _44667_ (_22215_, _22204_, _21594_);
  nor _44668_ (_22226_, _22215_, _21561_);
  not _44669_ (_22237_, _22226_);
  and _44670_ (_22248_, _22237_, _21424_);
  or _44671_ (_22259_, _22248_, _21402_);
  and _44672_ (_22269_, _17584_, _16601_);
  or _44673_ (_22280_, _22269_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _44674_ (_22291_, _21370_);
  and _44675_ (_22302_, _21206_, _22291_);
  nor _44676_ (_22324_, _21692_, _21537_);
  and _44677_ (_22325_, _22324_, _22302_);
  or _44678_ (_22336_, _22325_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44679_ (_22347_, _22336_, _22280_);
  and _44680_ (_22358_, _22347_, _22259_);
  and _44681_ (_22369_, _22358_, _21228_);
  nor _44682_ (_22379_, _22237_, _21424_);
  or _44683_ (_22390_, _22379_, _22248_);
  and _44684_ (_22401_, _22390_, _22369_);
  nor _44685_ (_22412_, _22369_, _21271_);
  nor _44686_ (_22423_, _22412_, _22401_);
  not _44687_ (_22435_, _22423_);
  and _44688_ (_22446_, _22423_, _21228_);
  not _44689_ (_22457_, _21391_);
  and _44690_ (_22468_, _22204_, _21594_);
  or _44691_ (_22478_, _22468_, _22215_);
  and _44692_ (_22489_, _22478_, _22369_);
  nor _44693_ (_22500_, _22369_, _21457_);
  nor _44694_ (_22511_, _22500_, _22489_);
  and _44695_ (_22522_, _22511_, _22457_);
  nor _44696_ (_22533_, _22511_, _22457_);
  nor _44697_ (_22544_, _22533_, _22522_);
  not _44698_ (_22555_, _22544_);
  not _44699_ (_22566_, _21550_);
  nor _44700_ (_22577_, _22369_, _21637_);
  and _44701_ (_22588_, _22182_, _21757_);
  nor _44702_ (_22598_, _22588_, _22193_);
  and _44703_ (_22609_, _22598_, _22369_);
  or _44704_ (_22620_, _22609_, _22577_);
  and _44705_ (_22631_, _22620_, _22566_);
  nor _44706_ (_22642_, _22620_, _22566_);
  nor _44707_ (_22653_, _22642_, _22631_);
  not _44708_ (_22664_, _22653_);
  not _44709_ (_22675_, _21713_);
  and _44710_ (_22686_, _22160_, _22128_);
  or _44711_ (_22697_, _22686_, _22171_);
  and _44712_ (_22707_, _22697_, _22369_);
  nor _44713_ (_22718_, _22369_, _21812_);
  nor _44714_ (_22729_, _22718_, _22707_);
  and _44715_ (_22740_, _22729_, _22675_);
  and _44716_ (_22751_, _22106_, _21921_);
  nor _44717_ (_22762_, _22751_, _22117_);
  not _44718_ (_22773_, _22762_);
  and _44719_ (_22784_, _22773_, _22369_);
  nor _44720_ (_22795_, _22369_, _21877_);
  nor _44721_ (_22806_, _22795_, _22784_);
  and _44722_ (_22816_, _22806_, _21779_);
  nor _44723_ (_22827_, _22806_, _21779_);
  nor _44724_ (_22838_, _22827_, _22816_);
  not _44725_ (_22849_, _22838_);
  nor _44726_ (_22860_, _22084_, _22062_);
  nor _44727_ (_22871_, _22860_, _22095_);
  not _44728_ (_22882_, _22871_);
  and _44729_ (_22893_, _22882_, _22369_);
  nor _44730_ (_22904_, _22369_, _21975_);
  nor _44731_ (_22915_, _22904_, _22893_);
  and _44732_ (_22925_, _22915_, _21844_);
  not _44733_ (_22936_, _22040_);
  and _44734_ (_22947_, _22369_, _21997_);
  or _44735_ (_22958_, _22947_, _22936_);
  nand _44736_ (_22969_, _22369_, _21997_);
  or _44737_ (_22980_, _22969_, _22040_);
  and _44738_ (_23001_, _22980_, _22958_);
  nor _44739_ (_23002_, _23001_, _21931_);
  and _44740_ (_23013_, _23001_, _21931_);
  nor _44741_ (_23033_, _23013_, _23002_);
  and _44742_ (_23034_, _21239_, _19360_);
  nor _44743_ (_23045_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _44744_ (_23066_, _23045_, _23034_);
  nor _44745_ (_23067_, _23066_, _22008_);
  not _44746_ (_23078_, _23067_);
  and _44747_ (_23099_, _23078_, _23033_);
  nor _44748_ (_23100_, _23099_, _23002_);
  nor _44749_ (_23111_, _22915_, _21844_);
  nor _44750_ (_23132_, _23111_, _22925_);
  not _44751_ (_23133_, _23132_);
  nor _44752_ (_23143_, _23133_, _23100_);
  nor _44753_ (_23164_, _23143_, _22925_);
  nor _44754_ (_23165_, _23164_, _22849_);
  nor _44755_ (_23176_, _23165_, _22816_);
  nor _44756_ (_23197_, _22729_, _22675_);
  nor _44757_ (_23198_, _23197_, _22740_);
  not _44758_ (_23209_, _23198_);
  nor _44759_ (_23220_, _23209_, _23176_);
  nor _44760_ (_23231_, _23220_, _22740_);
  nor _44761_ (_23242_, _23231_, _22664_);
  nor _44762_ (_23253_, _23242_, _22631_);
  nor _44763_ (_23264_, _23253_, _22555_);
  or _44764_ (_23275_, _23264_, _22522_);
  or _44765_ (_23286_, _23275_, _22446_);
  and _44766_ (_23297_, _23286_, _22347_);
  nor _44767_ (_23308_, _23297_, _22435_);
  and _44768_ (_23319_, _22446_, _22347_);
  and _44769_ (_23330_, _23319_, _23275_);
  or _44770_ (_23341_, _23330_, _23308_);
  and _44771_ (_00914_, _23341_, _41806_);
  or _44772_ (_23362_, _22423_, _21228_);
  and _44773_ (_23373_, _23362_, _23297_);
  and _44774_ (_03014_, _23373_, _41806_);
  and _44775_ (_03025_, _22369_, _41806_);
  and _44776_ (_03046_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _41806_);
  and _44777_ (_03068_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _41806_);
  and _44778_ (_03089_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _41806_);
  or _44779_ (_23434_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44780_ (_23445_, _21066_, rst);
  and _44781_ (_03100_, _23445_, _23434_);
  and _44782_ (_23466_, _23373_, _21997_);
  or _44783_ (_23477_, _23466_, _23066_);
  nand _44784_ (_23488_, _23466_, _23066_);
  and _44785_ (_23499_, _23488_, _23477_);
  and _44786_ (_03111_, _23499_, _41806_);
  nor _44787_ (_23520_, _23373_, _23001_);
  nor _44788_ (_23531_, _23078_, _23033_);
  nor _44789_ (_23542_, _23531_, _23099_);
  and _44790_ (_23553_, _23542_, _23373_);
  or _44791_ (_23564_, _23553_, _23520_);
  and _44792_ (_03122_, _23564_, _41806_);
  and _44793_ (_23585_, _23133_, _23100_);
  or _44794_ (_23596_, _23585_, _23143_);
  nand _44795_ (_23607_, _23596_, _23373_);
  or _44796_ (_23618_, _23373_, _22915_);
  and _44797_ (_23629_, _23618_, _23607_);
  and _44798_ (_03133_, _23629_, _41806_);
  and _44799_ (_23650_, _23164_, _22849_);
  or _44800_ (_23661_, _23650_, _23165_);
  nand _44801_ (_23672_, _23661_, _23373_);
  or _44802_ (_23683_, _23373_, _22806_);
  and _44803_ (_23694_, _23683_, _23672_);
  and _44804_ (_03144_, _23694_, _41806_);
  and _44805_ (_23715_, _23209_, _23176_);
  or _44806_ (_23726_, _23715_, _23220_);
  nand _44807_ (_23737_, _23726_, _23373_);
  or _44808_ (_23748_, _23373_, _22729_);
  and _44809_ (_23759_, _23748_, _23737_);
  and _44810_ (_03155_, _23759_, _41806_);
  and _44811_ (_23780_, _23231_, _22664_);
  or _44812_ (_23791_, _23780_, _23242_);
  nand _44813_ (_23802_, _23791_, _23373_);
  or _44814_ (_23813_, _23373_, _22620_);
  and _44815_ (_23824_, _23813_, _23802_);
  and _44816_ (_03166_, _23824_, _41806_);
  and _44817_ (_23845_, _23253_, _22555_);
  or _44818_ (_23856_, _23845_, _23264_);
  nand _44819_ (_23867_, _23856_, _23373_);
  or _44820_ (_23878_, _23373_, _22511_);
  and _44821_ (_23889_, _23878_, _23867_);
  and _44822_ (_03177_, _23889_, _41806_);
  not _44823_ (_23910_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44824_ (_23921_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15636_);
  and _44825_ (_23932_, _23921_, _23910_);
  and _44826_ (_23943_, _23932_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _44827_ (_23954_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44828_ (_23965_, _23954_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44829_ (_23976_, _23954_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44830_ (_23987_, _23976_, _23965_);
  and _44831_ (_23998_, _23987_, _23943_);
  nor _44832_ (_24009_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44833_ (_24020_, _24009_, _23921_);
  and _44834_ (_24031_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _44835_ (_24042_, _24031_, _23998_);
  not _44836_ (_24053_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _44837_ (_24064_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15636_);
  and _44838_ (_24075_, _24064_, _24053_);
  and _44839_ (_24086_, _24075_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44840_ (_24097_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _44841_ (_24108_, _24075_, _23910_);
  and _44842_ (_24119_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  nor _44843_ (_24130_, _24009_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _44844_ (_24141_, _24130_, _23921_);
  and _44845_ (_24152_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _44846_ (_24163_, _24152_, _24119_);
  nor _44847_ (_24185_, _24163_, _24097_);
  and _44848_ (_24197_, _24185_, _24042_);
  and _44849_ (_24209_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor _44850_ (_24221_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _44851_ (_24233_, _24221_, _23954_);
  and _44852_ (_24245_, _24233_, _23943_);
  nor _44853_ (_24257_, _24245_, _24209_);
  and _44854_ (_24258_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and _44855_ (_24269_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _44856_ (_24280_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or _44857_ (_24291_, _24280_, _24269_);
  nor _44858_ (_24302_, _24291_, _24258_);
  and _44859_ (_24313_, _24302_, _24257_);
  and _44860_ (_24324_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and _44861_ (_24335_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor _44862_ (_24346_, _24335_, _24324_);
  and _44863_ (_24357_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not _44864_ (_24368_, _24357_);
  not _44865_ (_24379_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44866_ (_24390_, _23943_, _24379_);
  and _44867_ (_24401_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _44868_ (_24412_, _24401_, _24390_);
  and _44869_ (_24423_, _24412_, _24368_);
  and _44870_ (_24434_, _24423_, _24346_);
  and _44871_ (_24445_, _24434_, _24313_);
  and _44872_ (_24456_, _24445_, _24197_);
  and _44873_ (_24467_, _23965_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _44874_ (_24478_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _44875_ (_24489_, _24478_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _44876_ (_24500_, _24489_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _44877_ (_24511_, _24500_);
  not _44878_ (_24522_, _23943_);
  nor _44879_ (_24533_, _24489_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _44880_ (_24544_, _24533_, _24522_);
  and _44881_ (_24555_, _24544_, _24511_);
  not _44882_ (_24566_, _24555_);
  and _44883_ (_24577_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44884_ (_24587_, _24577_, _23921_);
  and _44885_ (_24598_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _44886_ (_24609_, _24598_, _24587_);
  and _44887_ (_24621_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _44888_ (_24632_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _44889_ (_24643_, _24632_, _24621_);
  and _44890_ (_24654_, _24643_, _24609_);
  and _44891_ (_24665_, _24654_, _24566_);
  nor _44892_ (_24676_, _24478_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _44893_ (_24687_, _24676_);
  nor _44894_ (_24697_, _24489_, _24522_);
  and _44895_ (_24708_, _24697_, _24687_);
  not _44896_ (_24719_, _24708_);
  and _44897_ (_24730_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _44898_ (_24741_, _24730_, _24587_);
  and _44899_ (_24752_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _44900_ (_24763_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _44901_ (_24774_, _24763_, _24752_);
  and _44902_ (_24785_, _24774_, _24741_);
  and _44903_ (_24796_, _24785_, _24719_);
  nor _44904_ (_24807_, _24796_, _24665_);
  not _44905_ (_24818_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _44906_ (_24829_, _24500_, _24818_);
  and _44907_ (_24840_, _24500_, _24818_);
  nor _44908_ (_24851_, _24840_, _24829_);
  nor _44909_ (_24862_, _24851_, _24522_);
  not _44910_ (_24873_, _24862_);
  and _44911_ (_24884_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor _44912_ (_24895_, _24884_, _24587_);
  and _44913_ (_24906_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _44914_ (_24917_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor _44915_ (_24928_, _24917_, _24906_);
  and _44916_ (_24938_, _24928_, _24895_);
  and _44917_ (_24949_, _24938_, _24873_);
  not _44918_ (_24960_, _24949_);
  not _44919_ (_24971_, _24467_);
  nor _44920_ (_24982_, _23965_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _44921_ (_24993_, _24982_, _24522_);
  and _44922_ (_25004_, _24993_, _24971_);
  not _44923_ (_25015_, _25004_);
  and _44924_ (_25026_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and _44925_ (_25037_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _44926_ (_25048_, _25037_, _25026_);
  and _44927_ (_25058_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _44928_ (_25069_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor _44929_ (_25080_, _25069_, _25058_);
  and _44930_ (_25091_, _25080_, _25048_);
  and _44931_ (_25112_, _25091_, _25015_);
  not _44932_ (_25113_, _25112_);
  nor _44933_ (_25124_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or _44934_ (_25135_, _25124_, _24522_);
  nor _44935_ (_25156_, _25135_, _24478_);
  and _44936_ (_25157_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor _44937_ (_25168_, _25157_, _25156_);
  and _44938_ (_25188_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and _44939_ (_25189_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor _44940_ (_25200_, _25189_, _25188_);
  and _44941_ (_25211_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _44942_ (_25222_, _25211_, _24587_);
  and _44943_ (_25243_, _25222_, _25200_);
  and _44944_ (_25244_, _25243_, _25168_);
  nor _44945_ (_25255_, _25244_, _25113_);
  and _44946_ (_25266_, _25255_, _24960_);
  and _44947_ (_25277_, _25266_, _24807_);
  nand _44948_ (_25287_, _25277_, _24456_);
  and _44949_ (_25298_, _23341_, _21055_);
  not _44950_ (_25309_, _25298_);
  and _44951_ (_25320_, _20451_, _15702_);
  not _44952_ (_25331_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44953_ (_25342_, _15647_, _25331_);
  and _44954_ (_25353_, _25342_, _15691_);
  not _44955_ (_25374_, _25353_);
  nor _44956_ (_25375_, _17758_, _17584_);
  and _44957_ (_25386_, _17758_, _17584_);
  nor _44958_ (_25397_, _25386_, _25375_);
  not _44959_ (_25408_, _16601_);
  nor _44960_ (_25419_, _16919_, _25408_);
  nor _44961_ (_25430_, _16919_, _16601_);
  and _44962_ (_25441_, _16919_, _16601_);
  nor _44963_ (_25452_, _25441_, _25430_);
  not _44964_ (_25462_, _17247_);
  nor _44965_ (_25473_, _17943_, _25462_);
  nor _44966_ (_25484_, _17943_, _17247_);
  and _44967_ (_25495_, _17943_, _17247_);
  nor _44968_ (_25506_, _25495_, _25484_);
  not _44969_ (_25517_, _16260_);
  and _44970_ (_25528_, _18107_, _25517_);
  nor _44971_ (_25548_, _25528_, _25506_);
  nor _44972_ (_25549_, _25548_, _25473_);
  nor _44973_ (_25560_, _25549_, _25452_);
  nor _44974_ (_25571_, _25560_, _25419_);
  and _44975_ (_25582_, _25549_, _25452_);
  nor _44976_ (_25593_, _25582_, _25560_);
  not _44977_ (_25604_, _25593_);
  and _44978_ (_25615_, _25528_, _25506_);
  nor _44979_ (_25626_, _25615_, _25548_);
  not _44980_ (_25636_, _25626_);
  nor _44981_ (_25647_, _18107_, _16260_);
  and _44982_ (_25658_, _18107_, _16260_);
  nor _44983_ (_25669_, _25658_, _25647_);
  not _44984_ (_25680_, _25669_);
  and _44985_ (_25691_, _18477_, _17094_);
  nor _44986_ (_25702_, _18477_, _17094_);
  nor _44987_ (_25713_, _25702_, _25691_);
  nor _44988_ (_25723_, _18978_, _16096_);
  and _44989_ (_25744_, _18978_, _16096_);
  nor _44990_ (_25745_, _25744_, _25723_);
  nor _44991_ (_25756_, _18815_, _17410_);
  and _44992_ (_25767_, _18815_, _17410_);
  nor _44993_ (_25778_, _25767_, _25756_);
  not _44994_ (_25789_, _16425_);
  and _44995_ (_25800_, _19360_, _25789_);
  nor _44996_ (_25810_, _25800_, _25778_);
  not _44997_ (_25821_, _17410_);
  nor _44998_ (_25832_, _18815_, _25821_);
  nor _44999_ (_25843_, _25832_, _25810_);
  nor _45000_ (_25854_, _25843_, _25745_);
  not _45001_ (_25865_, _16096_);
  nor _45002_ (_25876_, _18978_, _25865_);
  nor _45003_ (_25887_, _25876_, _25854_);
  nor _45004_ (_25897_, _25887_, _25713_);
  and _45005_ (_25908_, _25887_, _25713_);
  nor _45006_ (_25919_, _25908_, _25897_);
  not _45007_ (_25930_, _25919_);
  and _45008_ (_25941_, _25843_, _25745_);
  nor _45009_ (_25952_, _25941_, _25854_);
  not _45010_ (_25963_, _25952_);
  and _45011_ (_25974_, _25800_, _25778_);
  nor _45012_ (_25984_, _25974_, _25810_);
  not _45013_ (_25995_, _25984_);
  nor _45014_ (_26006_, _19360_, _16425_);
  and _45015_ (_26017_, _19360_, _16425_);
  nor _45016_ (_26028_, _26017_, _26006_);
  not _45017_ (_26039_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _45018_ (_26050_, _15909_, _26039_);
  not _45019_ (_26061_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _45020_ (_26071_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45021_ (_26092_, _26071_, _17475_);
  nor _45022_ (_26093_, _26092_, _26061_);
  nor _45023_ (_26104_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45024_ (_26115_, _26104_, _16150_);
  not _45025_ (_26126_, _26115_);
  not _45026_ (_26137_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _45027_ (_26147_, _26137_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45028_ (_26158_, _26147_, _16490_);
  not _45029_ (_26169_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45030_ (_26180_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _26169_);
  and _45031_ (_26201_, _26180_, _17138_);
  nor _45032_ (_26202_, _26201_, _26158_);
  and _45033_ (_26213_, _26202_, _26126_);
  and _45034_ (_26224_, _26213_, _26093_);
  and _45035_ (_26234_, _26071_, _16985_);
  nor _45036_ (_26245_, _26234_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _45037_ (_26256_, _26180_, _17301_);
  not _45038_ (_26267_, _26256_);
  and _45039_ (_26278_, _26147_, _15953_);
  and _45040_ (_26289_, _26104_, _16315_);
  nor _45041_ (_26300_, _26289_, _26278_);
  and _45042_ (_26311_, _26300_, _26267_);
  and _45043_ (_26321_, _26311_, _26245_);
  nor _45044_ (_26332_, _26321_, _26224_);
  nor _45045_ (_26343_, _26332_, _15909_);
  nor _45046_ (_26354_, _26343_, _26050_);
  and _45047_ (_26365_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _45048_ (_26376_, _26365_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _45049_ (_26387_, _26376_);
  and _45050_ (_26398_, _26387_, _26354_);
  and _45051_ (_26408_, _26387_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _45052_ (_26419_, _26408_, _26398_);
  nor _45053_ (_26430_, _26419_, _26028_);
  and _45054_ (_26441_, _26430_, _25995_);
  and _45055_ (_26452_, _26441_, _25963_);
  and _45056_ (_26463_, _26452_, _25930_);
  not _45057_ (_26474_, _17094_);
  or _45058_ (_26485_, _18477_, _26474_);
  and _45059_ (_26496_, _18477_, _26474_);
  or _45060_ (_26506_, _25887_, _26496_);
  and _45061_ (_26517_, _26506_, _26485_);
  or _45062_ (_26528_, _26517_, _26463_);
  and _45063_ (_26539_, _26528_, _25680_);
  and _45064_ (_26550_, _26539_, _25636_);
  and _45065_ (_26561_, _26550_, _25604_);
  nor _45066_ (_26572_, _26561_, _25571_);
  nor _45067_ (_26583_, _26572_, _25397_);
  and _45068_ (_26593_, _26572_, _25397_);
  nor _45069_ (_26604_, _26593_, _26583_);
  nor _45070_ (_26615_, _26604_, _25374_);
  not _45071_ (_26626_, _26615_);
  not _45072_ (_26647_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _45073_ (_26648_, _21012_, _26647_);
  and _45074_ (_26659_, _26648_, _15691_);
  not _45075_ (_26670_, _25452_);
  and _45076_ (_26680_, _25647_, _25506_);
  nor _45077_ (_26691_, _26680_, _25484_);
  nor _45078_ (_26702_, _26691_, _26670_);
  not _45079_ (_26713_, _25745_);
  and _45080_ (_26724_, _26006_, _25778_);
  nor _45081_ (_26735_, _26724_, _25756_);
  nor _45082_ (_26746_, _26735_, _26713_);
  nor _45083_ (_26757_, _26746_, _25723_);
  nor _45084_ (_26768_, _26757_, _25713_);
  and _45085_ (_26778_, _26757_, _25713_);
  nor _45086_ (_26789_, _26778_, _26768_);
  not _45087_ (_26800_, _26028_);
  nor _45088_ (_26811_, _26419_, _26800_);
  and _45089_ (_26822_, _26811_, _25778_);
  and _45090_ (_26833_, _26735_, _26713_);
  nor _45091_ (_26844_, _26833_, _26746_);
  and _45092_ (_26855_, _26844_, _26822_);
  not _45093_ (_26866_, _26855_);
  nor _45094_ (_26877_, _26866_, _26789_);
  nor _45095_ (_26888_, _26757_, _25691_);
  or _45096_ (_26898_, _26888_, _25702_);
  or _45097_ (_26909_, _26898_, _26877_);
  and _45098_ (_26920_, _26909_, _25669_);
  nor _45099_ (_26941_, _25647_, _25506_);
  nor _45100_ (_26942_, _26941_, _26680_);
  and _45101_ (_26953_, _26942_, _26920_);
  and _45102_ (_26964_, _26691_, _26670_);
  nor _45103_ (_26975_, _26964_, _26702_);
  and _45104_ (_26986_, _26975_, _26953_);
  or _45105_ (_26997_, _26986_, _26702_);
  nor _45106_ (_27007_, _26997_, _25430_);
  and _45107_ (_27018_, _27007_, _25397_);
  nor _45108_ (_27029_, _27007_, _25397_);
  or _45109_ (_27050_, _27029_, _27018_);
  and _45110_ (_27051_, _27050_, _26659_);
  and _45111_ (_27062_, _15680_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45112_ (_27073_, _27062_, _25342_);
  nor _45113_ (_27084_, _19360_, _18815_);
  and _45114_ (_27095_, _27084_, _18989_);
  and _45115_ (_27106_, _27095_, _18488_);
  and _45116_ (_27117_, _27106_, _18117_);
  and _45117_ (_27127_, _27117_, _18520_);
  and _45118_ (_27138_, _27127_, _16930_);
  and _45119_ (_27149_, _27138_, _26419_);
  not _45120_ (_27160_, _26419_);
  and _45121_ (_27171_, _16919_, _17943_);
  and _45122_ (_27182_, _19360_, _18815_);
  and _45123_ (_27193_, _27182_, _18978_);
  and _45124_ (_27204_, _27193_, _18477_);
  and _45125_ (_27215_, _27204_, _18107_);
  and _45126_ (_27226_, _27215_, _27171_);
  and _45127_ (_27237_, _27226_, _27160_);
  nor _45128_ (_27247_, _27237_, _27149_);
  and _45129_ (_27268_, _27247_, _17758_);
  nor _45130_ (_27269_, _27247_, _17758_);
  nor _45131_ (_27280_, _27269_, _27268_);
  and _45132_ (_27291_, _27280_, _27073_);
  not _45133_ (_27302_, _17584_);
  nor _45134_ (_27313_, _26419_, _27302_);
  not _45135_ (_27324_, _27313_);
  and _45136_ (_27335_, _26419_, _17758_);
  and _45137_ (_27346_, _27062_, _15658_);
  not _45138_ (_27356_, _27346_);
  nor _45139_ (_27367_, _27356_, _27335_);
  and _45140_ (_27378_, _27367_, _27324_);
  nor _45141_ (_27389_, _27378_, _27291_);
  and _45142_ (_27400_, _26648_, _21044_);
  not _45143_ (_27411_, _27400_);
  and _45144_ (_27422_, _18978_, _18815_);
  nor _45145_ (_27433_, _27422_, _18477_);
  and _45146_ (_27444_, _27433_, _27400_);
  and _45147_ (_27455_, _27444_, _18117_);
  nor _45148_ (_27466_, _27455_, _18520_);
  and _45149_ (_27476_, _27466_, _16919_);
  nor _45150_ (_27487_, _27171_, _17758_);
  nor _45151_ (_27498_, _27487_, _27444_);
  and _45152_ (_27509_, _27498_, _26419_);
  nor _45153_ (_27530_, _27509_, _27476_);
  nor _45154_ (_27531_, _27530_, _17758_);
  and _45155_ (_27542_, _27530_, _17758_);
  nor _45156_ (_27552_, _27542_, _27531_);
  nor _45157_ (_27563_, _27552_, _27411_);
  not _45158_ (_27574_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45159_ (_27585_, _15680_, _27574_);
  and _45160_ (_27596_, _27585_, _21023_);
  and _45161_ (_27607_, _27596_, _25397_);
  and _45162_ (_27618_, _21044_, _15658_);
  and _45163_ (_27629_, _27618_, _25375_);
  and _45164_ (_27640_, _27585_, _26648_);
  not _45165_ (_27651_, _27640_);
  nor _45166_ (_27662_, _27651_, _25386_);
  and _45167_ (_27672_, _25342_, _21044_);
  and _45168_ (_27683_, _27672_, _17758_);
  or _45169_ (_27694_, _27683_, _27662_);
  or _45170_ (_27705_, _27694_, _27629_);
  nor _45171_ (_27716_, _27705_, _27607_);
  and _45172_ (_27727_, _27062_, _26648_);
  not _45173_ (_27738_, _27727_);
  nor _45174_ (_27749_, _27738_, _26419_);
  and _45175_ (_27760_, _27585_, _15647_);
  not _45176_ (_27771_, _27760_);
  nor _45177_ (_27782_, _27771_, _16919_);
  not _45178_ (_27793_, _27782_);
  and _45179_ (_27813_, _21023_, _15691_);
  not _45180_ (_27814_, _27813_);
  nor _45181_ (_27825_, _27814_, _17758_);
  and _45182_ (_27836_, _27062_, _21023_);
  not _45183_ (_27847_, _27836_);
  nor _45184_ (_27858_, _27847_, _19360_);
  nor _45185_ (_27869_, _27858_, _27825_);
  and _45186_ (_27880_, _27869_, _27793_);
  not _45187_ (_27891_, _27880_);
  nor _45188_ (_27902_, _27891_, _27749_);
  and _45189_ (_27913_, _27902_, _27716_);
  not _45190_ (_27923_, _27913_);
  nor _45191_ (_27934_, _27923_, _27563_);
  and _45192_ (_27945_, _27934_, _27389_);
  not _45193_ (_27956_, _27945_);
  nor _45194_ (_27967_, _27956_, _27051_);
  and _45195_ (_27978_, _27967_, _26626_);
  not _45196_ (_27989_, _27978_);
  nor _45197_ (_28000_, _27989_, _25320_);
  and _45198_ (_28011_, _28000_, _25309_);
  not _45199_ (_28022_, _28011_);
  or _45200_ (_28033_, _28022_, _25287_);
  not _45201_ (_28044_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _45202_ (_28054_, \oc8051_top_1.oc8051_decoder1.wr , _15636_);
  not _45203_ (_28065_, _28054_);
  nor _45204_ (_28076_, _28065_, _23932_);
  and _45205_ (_28087_, _28076_, _28044_);
  not _45206_ (_28098_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _45207_ (_28109_, _25287_, _28098_);
  and _45208_ (_28120_, _28109_, _28087_);
  and _45209_ (_28131_, _28120_, _28033_);
  nor _45210_ (_28142_, _28076_, _28098_);
  not _45211_ (_28153_, _26659_);
  nor _45212_ (_28164_, _27007_, _25386_);
  nor _45213_ (_28175_, _28164_, _25375_);
  nor _45214_ (_28185_, _28175_, _28153_);
  not _45215_ (_28196_, _28185_);
  and _45216_ (_28207_, _17758_, _27302_);
  nor _45217_ (_28218_, _28207_, _26583_);
  nor _45218_ (_28229_, _28218_, _25374_);
  and _45219_ (_28250_, _26419_, _16919_);
  and _45220_ (_28251_, _28250_, _27466_);
  nor _45221_ (_28262_, _28251_, _27335_);
  nor _45222_ (_28273_, _26419_, _17758_);
  not _45223_ (_28284_, _28273_);
  nor _45224_ (_28295_, _28284_, _27476_);
  nor _45225_ (_28306_, _28295_, _27411_);
  and _45226_ (_28317_, _28306_, _28262_);
  or _45227_ (_28327_, _28317_, _27444_);
  nor _45228_ (_28338_, _27814_, _26419_);
  not _45229_ (_28349_, _28338_);
  and _45230_ (_28360_, _26376_, _26354_);
  and _45231_ (_28371_, _27585_, _25342_);
  and _45232_ (_28382_, _27618_, _26354_);
  nor _45233_ (_28393_, _28382_, _28371_);
  nor _45234_ (_28404_, _28393_, _28360_);
  nor _45235_ (_28415_, _27738_, _19360_);
  and _45236_ (_28435_, _27585_, _15658_);
  not _45237_ (_28436_, _28435_);
  nor _45238_ (_28447_, _28436_, _17758_);
  nor _45239_ (_28458_, _28447_, _28415_);
  not _45240_ (_28469_, _28458_);
  nor _45241_ (_28480_, _28469_, _28404_);
  and _45242_ (_28491_, _28480_, _28349_);
  nor _45243_ (_28502_, _26408_, _26354_);
  not _45244_ (_28513_, _27596_);
  nor _45245_ (_28524_, _28513_, _26398_);
  nor _45246_ (_28535_, _28524_, _27640_);
  nor _45247_ (_28545_, _28535_, _28502_);
  nor _45248_ (_28556_, _27672_, _27160_);
  and _45249_ (_28567_, _27847_, _26408_);
  nor _45250_ (_28578_, _28567_, _26398_);
  not _45251_ (_28589_, _28578_);
  nor _45252_ (_28600_, _28589_, _28556_);
  nor _45253_ (_28611_, _28600_, _28545_);
  and _45254_ (_28622_, _28611_, _28491_);
  not _45255_ (_28633_, _28622_);
  nor _45256_ (_28644_, _28633_, _28327_);
  not _45257_ (_28654_, _28644_);
  nor _45258_ (_28665_, _28654_, _28229_);
  and _45259_ (_28676_, _28665_, _28196_);
  not _45260_ (_28687_, _24197_);
  nor _45261_ (_28698_, _24434_, _24313_);
  and _45262_ (_28709_, _28698_, _28687_);
  and _45263_ (_28720_, _28709_, _25277_);
  nand _45264_ (_28731_, _28720_, _28676_);
  and _45265_ (_28742_, _28076_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or _45266_ (_28753_, _28720_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _45267_ (_28764_, _28753_, _28742_);
  and _45268_ (_28774_, _28764_, _28731_);
  or _45269_ (_28785_, _28774_, _28142_);
  or _45270_ (_28796_, _28785_, _28131_);
  and _45271_ (_06695_, _28796_, _41806_);
  and _45272_ (_28817_, _23499_, _21055_);
  not _45273_ (_28828_, _28817_);
  and _45274_ (_28839_, _20779_, _15702_);
  and _45275_ (_28850_, _26419_, _26800_);
  nor _45276_ (_28861_, _28850_, _26811_);
  not _45277_ (_28872_, _28861_);
  nor _45278_ (_28883_, _26659_, _25353_);
  nor _45279_ (_28893_, _28883_, _28872_);
  not _45280_ (_28904_, _28893_);
  and _45281_ (_28915_, _27596_, _26028_);
  not _45282_ (_28926_, _28915_);
  and _45283_ (_28937_, _27618_, _26006_);
  not _45284_ (_28948_, _28937_);
  nor _45285_ (_28969_, _27651_, _26017_);
  and _45286_ (_28970_, _27672_, _19360_);
  nor _45287_ (_28981_, _28970_, _28969_);
  and _45288_ (_28992_, _28981_, _28948_);
  and _45289_ (_29002_, _28992_, _28926_);
  nor _45290_ (_29013_, _28436_, _26419_);
  not _45291_ (_29024_, _29013_);
  nor _45292_ (_29035_, _27356_, _16425_);
  and _45293_ (_29046_, _27073_, _19360_);
  nor _45294_ (_29057_, _29046_, _29035_);
  and _45295_ (_29068_, _27062_, _26647_);
  not _45296_ (_29079_, _29068_);
  nor _45297_ (_29090_, _29079_, _18815_);
  not _45298_ (_29101_, _29090_);
  and _45299_ (_29112_, _28371_, _18215_);
  nor _45300_ (_29122_, _27813_, _27400_);
  nor _45301_ (_29133_, _29122_, _19360_);
  nor _45302_ (_29144_, _29133_, _29112_);
  and _45303_ (_29155_, _29144_, _29101_);
  and _45304_ (_29166_, _29155_, _29057_);
  and _45305_ (_29177_, _29166_, _29024_);
  and _45306_ (_29188_, _29177_, _29002_);
  and _45307_ (_29198_, _29188_, _28904_);
  not _45308_ (_29209_, _29198_);
  nor _45309_ (_29220_, _29209_, _28839_);
  and _45310_ (_29231_, _29220_, _28828_);
  not _45311_ (_29242_, _29231_);
  or _45312_ (_29253_, _29242_, _25287_);
  not _45313_ (_29264_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _45314_ (_29275_, _25287_, _29264_);
  and _45315_ (_29285_, _29275_, _28087_);
  and _45316_ (_29296_, _29285_, _29253_);
  nor _45317_ (_29307_, _28076_, _29264_);
  not _45318_ (_29318_, _28676_);
  or _45319_ (_29329_, _29318_, _25287_);
  and _45320_ (_29340_, _29275_, _28742_);
  and _45321_ (_29351_, _29340_, _29329_);
  or _45322_ (_29362_, _29351_, _29307_);
  or _45323_ (_29372_, _29362_, _29296_);
  and _45324_ (_08932_, _29372_, _41806_);
  and _45325_ (_29393_, _20811_, _15702_);
  not _45326_ (_29404_, _29393_);
  and _45327_ (_29415_, _23564_, _21055_);
  nor _45328_ (_29426_, _26006_, _25778_);
  or _45329_ (_29437_, _29426_, _26724_);
  and _45330_ (_29448_, _29437_, _26811_);
  nor _45331_ (_29458_, _29437_, _26811_);
  or _45332_ (_29469_, _29458_, _29448_);
  and _45333_ (_29480_, _29469_, _26659_);
  nor _45334_ (_29491_, _26430_, _25995_);
  nor _45335_ (_29512_, _29491_, _26441_);
  nor _45336_ (_29513_, _29512_, _25374_);
  not _45337_ (_29524_, _29513_);
  nor _45338_ (_29535_, _27433_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _45339_ (_29546_, _29535_, _27400_);
  and _45340_ (_29556_, _29546_, _27814_);
  or _45341_ (_29567_, _29556_, _18815_);
  and _45342_ (_29578_, _27596_, _25778_);
  nor _45343_ (_29589_, _27651_, _25767_);
  or _45344_ (_29600_, _29589_, _29578_);
  not _45345_ (_29611_, _29600_);
  and _45346_ (_29622_, _27618_, _25756_);
  and _45347_ (_29633_, _27672_, _18815_);
  nor _45348_ (_29643_, _29633_, _29622_);
  and _45349_ (_29654_, _29643_, _29611_);
  nor _45350_ (_29665_, _29535_, _19022_);
  nand _45351_ (_29676_, _29665_, _27400_);
  nor _45352_ (_29687_, _29079_, _18978_);
  nor _45353_ (_29698_, _27771_, _19360_);
  nor _45354_ (_29709_, _29698_, _29687_);
  and _45355_ (_29720_, _29709_, _29676_);
  and _45356_ (_29730_, _29720_, _29654_);
  and _45357_ (_29741_, _29730_, _29567_);
  and _45358_ (_29752_, _29741_, _29524_);
  nor _45359_ (_29773_, _27356_, _17410_);
  nor _45360_ (_29774_, _27182_, _27084_);
  not _45361_ (_29785_, _29774_);
  nor _45362_ (_29796_, _29785_, _26419_);
  and _45363_ (_29806_, _29785_, _26419_);
  nor _45364_ (_29817_, _29806_, _29796_);
  and _45365_ (_29828_, _29817_, _27073_);
  nor _45366_ (_29839_, _29828_, _29773_);
  nand _45367_ (_29850_, _29839_, _29752_);
  nor _45368_ (_29861_, _29850_, _29480_);
  not _45369_ (_29872_, _29861_);
  nor _45370_ (_29883_, _29872_, _29415_);
  and _45371_ (_29893_, _29883_, _29404_);
  not _45372_ (_29904_, _29893_);
  or _45373_ (_29915_, _29904_, _25287_);
  not _45374_ (_29926_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _45375_ (_29937_, _25287_, _29926_);
  and _45376_ (_29948_, _29937_, _28087_);
  and _45377_ (_29959_, _29948_, _29915_);
  nor _45378_ (_29970_, _28076_, _29926_);
  not _45379_ (_29980_, _24434_);
  and _45380_ (_29991_, _29980_, _24313_);
  and _45381_ (_30002_, _29991_, _24197_);
  and _45382_ (_30013_, _30002_, _25277_);
  or _45383_ (_30024_, _30013_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _45384_ (_30035_, _30024_, _28742_);
  nand _45385_ (_30046_, _30013_, _28676_);
  and _45386_ (_30057_, _30046_, _30035_);
  or _45387_ (_30077_, _30057_, _29970_);
  or _45388_ (_30078_, _30077_, _29959_);
  and _45389_ (_08943_, _30078_, _41806_);
  and _45390_ (_30099_, _20842_, _15702_);
  not _45391_ (_30110_, _30099_);
  and _45392_ (_30121_, _23629_, _21055_);
  nor _45393_ (_30132_, _27356_, _16096_);
  and _45394_ (_30143_, _27084_, _26419_);
  and _45395_ (_30153_, _27182_, _27160_);
  nor _45396_ (_30164_, _30153_, _30143_);
  and _45397_ (_30175_, _30164_, _18978_);
  nor _45398_ (_30186_, _30164_, _18978_);
  nor _45399_ (_30197_, _30186_, _30175_);
  and _45400_ (_30208_, _30197_, _27073_);
  nor _45401_ (_30219_, _30208_, _30132_);
  nor _45402_ (_30230_, _26441_, _25963_);
  nor _45403_ (_30240_, _30230_, _26452_);
  nor _45404_ (_30251_, _30240_, _25374_);
  not _45405_ (_30262_, _30251_);
  nor _45406_ (_30273_, _29079_, _18477_);
  and _45407_ (_30284_, _27618_, _25723_);
  and _45408_ (_30295_, _27672_, _18978_);
  nor _45409_ (_30306_, _30295_, _30284_);
  nor _45410_ (_30317_, _27651_, _25744_);
  and _45411_ (_30327_, _27596_, _25745_);
  nor _45412_ (_30338_, _30327_, _30317_);
  nor _45413_ (_30349_, _27771_, _18815_);
  nor _45414_ (_30360_, _27814_, _18978_);
  nor _45415_ (_30371_, _30360_, _30349_);
  and _45416_ (_30382_, _30371_, _30338_);
  nand _45417_ (_30402_, _30382_, _30306_);
  nor _45418_ (_30403_, _30402_, _30273_);
  and _45419_ (_30414_, _30403_, _30262_);
  nor _45420_ (_30425_, _26844_, _26822_);
  nor _45421_ (_30436_, _30425_, _28153_);
  and _45422_ (_30447_, _30436_, _26866_);
  and _45423_ (_30458_, _27422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45424_ (_30470_, _29665_, _18978_);
  nor _45425_ (_30491_, _30470_, _30458_);
  nor _45426_ (_30501_, _30491_, _27411_);
  nor _45427_ (_30512_, _30501_, _30447_);
  and _45428_ (_30523_, _30512_, _30414_);
  and _45429_ (_30534_, _30523_, _30219_);
  not _45430_ (_30545_, _30534_);
  nor _45431_ (_30556_, _30545_, _30121_);
  and _45432_ (_30567_, _30556_, _30110_);
  not _45433_ (_30578_, _30567_);
  or _45434_ (_30589_, _30578_, _25287_);
  not _45435_ (_30599_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _45436_ (_30610_, _25287_, _30599_);
  and _45437_ (_30621_, _30610_, _28087_);
  and _45438_ (_30632_, _30621_, _30589_);
  nor _45439_ (_30643_, _28076_, _30599_);
  nand _45440_ (_30654_, _25277_, _24197_);
  or _45441_ (_30665_, _28698_, _30654_);
  and _45442_ (_30676_, _30665_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _45443_ (_30686_, _24313_);
  and _45444_ (_30697_, _24197_, _24434_);
  and _45445_ (_30708_, _30697_, _30686_);
  and _45446_ (_30719_, _30708_, _29318_);
  and _45447_ (_30730_, _24197_, _24313_);
  and _45448_ (_30741_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _45449_ (_30752_, _30741_, _30719_);
  and _45450_ (_30763_, _30752_, _25277_);
  or _45451_ (_30773_, _30763_, _30676_);
  and _45452_ (_30784_, _30773_, _28742_);
  or _45453_ (_30795_, _30784_, _30643_);
  or _45454_ (_30806_, _30795_, _30632_);
  and _45455_ (_08954_, _30806_, _41806_);
  and _45456_ (_30827_, _20885_, _15702_);
  not _45457_ (_30838_, _30827_);
  and _45458_ (_30849_, _23694_, _21055_);
  and _45459_ (_30859_, _26866_, _26789_);
  or _45460_ (_30870_, _30859_, _28153_);
  nor _45461_ (_30891_, _30870_, _26877_);
  not _45462_ (_30892_, _30891_);
  nor _45463_ (_30903_, _26452_, _25930_);
  nor _45464_ (_30914_, _30903_, _26463_);
  nor _45465_ (_30925_, _30914_, _25374_);
  not _45466_ (_30936_, _30925_);
  nor _45467_ (_30946_, _27356_, _17094_);
  nor _45468_ (_30957_, _27193_, _26419_);
  nor _45469_ (_30968_, _27095_, _27160_);
  nor _45470_ (_30979_, _30968_, _30957_);
  and _45471_ (_30990_, _30979_, _18488_);
  not _45472_ (_31001_, _30990_);
  not _45473_ (_31012_, _27073_);
  nor _45474_ (_31022_, _30979_, _18488_);
  nor _45475_ (_31033_, _31022_, _31012_);
  and _45476_ (_31044_, _31033_, _31001_);
  nor _45477_ (_31055_, _31044_, _30946_);
  not _45478_ (_31066_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45479_ (_31077_, _27422_, _31066_);
  nor _45480_ (_31088_, _31077_, _18488_);
  nor _45481_ (_31099_, _27814_, _18477_);
  nor _45482_ (_31119_, _27433_, _27411_);
  nor _45483_ (_31120_, _31119_, _31099_);
  nor _45484_ (_31131_, _31120_, _31088_);
  not _45485_ (_31142_, _31131_);
  nor _45486_ (_31153_, _27651_, _25691_);
  and _45487_ (_31164_, _27596_, _25713_);
  nor _45488_ (_31175_, _31164_, _31153_);
  and _45489_ (_31186_, _27618_, _25702_);
  and _45490_ (_31197_, _27672_, _18477_);
  nor _45491_ (_31207_, _31197_, _31186_);
  nor _45492_ (_31218_, _29079_, _18107_);
  nor _45493_ (_31229_, _27771_, _18978_);
  nor _45494_ (_31240_, _31229_, _31218_);
  and _45495_ (_31251_, _31240_, _31207_);
  and _45496_ (_31262_, _31251_, _31175_);
  and _45497_ (_31273_, _31262_, _31142_);
  and _45498_ (_31284_, _31273_, _31055_);
  and _45499_ (_31294_, _31284_, _30936_);
  and _45500_ (_31305_, _31294_, _30892_);
  not _45501_ (_31316_, _31305_);
  nor _45502_ (_31327_, _31316_, _30849_);
  and _45503_ (_31338_, _31327_, _30838_);
  not _45504_ (_31349_, _31338_);
  or _45505_ (_31360_, _31349_, _25287_);
  not _45506_ (_31371_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _45507_ (_31381_, _25287_, _31371_);
  and _45508_ (_31392_, _31381_, _28087_);
  and _45509_ (_31403_, _31392_, _31360_);
  nor _45510_ (_31414_, _28076_, _31371_);
  and _45511_ (_31425_, _30654_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _45512_ (_31436_, _28698_, _24197_);
  not _45513_ (_31447_, _31436_);
  nor _45514_ (_31458_, _31447_, _28676_);
  nor _45515_ (_31468_, _30730_, _30697_);
  nor _45516_ (_31479_, _31468_, _31371_);
  or _45517_ (_31490_, _31479_, _31458_);
  and _45518_ (_31501_, _31490_, _25277_);
  or _45519_ (_31512_, _31501_, _31425_);
  and _45520_ (_31523_, _31512_, _28742_);
  or _45521_ (_31534_, _31523_, _31414_);
  or _45522_ (_31545_, _31534_, _31403_);
  and _45523_ (_08965_, _31545_, _41806_);
  and _45524_ (_31565_, _23759_, _21055_);
  not _45525_ (_31576_, _31565_);
  and _45526_ (_31587_, _20917_, _15702_);
  or _45527_ (_31598_, _26909_, _25669_);
  nor _45528_ (_31609_, _28153_, _26920_);
  and _45529_ (_31620_, _31609_, _31598_);
  nor _45530_ (_31630_, _26528_, _25669_);
  and _45531_ (_31641_, _26528_, _25669_);
  nor _45532_ (_31652_, _31641_, _31630_);
  and _45533_ (_31663_, _31652_, _25353_);
  and _45534_ (_31674_, _26419_, _18117_);
  nor _45535_ (_31695_, _26419_, _16260_);
  or _45536_ (_31696_, _31695_, _31674_);
  and _45537_ (_31707_, _31696_, _27346_);
  and _45538_ (_31717_, _27106_, _26419_);
  and _45539_ (_31728_, _27204_, _27160_);
  nor _45540_ (_31739_, _31728_, _31717_);
  nor _45541_ (_31750_, _31739_, _18107_);
  and _45542_ (_31761_, _31739_, _18107_);
  or _45543_ (_31772_, _31761_, _31012_);
  nor _45544_ (_31783_, _31772_, _31750_);
  nor _45545_ (_31794_, _31783_, _31707_);
  or _45546_ (_31804_, _27444_, _18117_);
  nor _45547_ (_31815_, _27455_, _27411_);
  and _45548_ (_31826_, _31815_, _31804_);
  and _45549_ (_31837_, _27596_, _25669_);
  nor _45550_ (_31848_, _27651_, _25658_);
  not _45551_ (_31859_, _31848_);
  and _45552_ (_31870_, _27618_, _25647_);
  and _45553_ (_31881_, _27672_, _18107_);
  nor _45554_ (_31891_, _31881_, _31870_);
  nand _45555_ (_31902_, _31891_, _31859_);
  nor _45556_ (_31913_, _31902_, _31837_);
  nor _45557_ (_31924_, _29079_, _17943_);
  nor _45558_ (_31935_, _27814_, _18107_);
  nor _45559_ (_31946_, _27771_, _18477_);
  or _45560_ (_31957_, _31946_, _31935_);
  nor _45561_ (_31968_, _31957_, _31924_);
  nand _45562_ (_31979_, _31968_, _31913_);
  nor _45563_ (_31989_, _31979_, _31826_);
  nand _45564_ (_32000_, _31989_, _31794_);
  or _45565_ (_32011_, _32000_, _31663_);
  or _45566_ (_32022_, _32011_, _31620_);
  nor _45567_ (_32033_, _32022_, _31587_);
  and _45568_ (_32044_, _32033_, _31576_);
  not _45569_ (_32055_, _32044_);
  or _45570_ (_32065_, _32055_, _25287_);
  not _45571_ (_32076_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _45572_ (_32087_, _25287_, _32076_);
  and _45573_ (_32098_, _32087_, _28087_);
  and _45574_ (_32109_, _32098_, _32065_);
  nor _45575_ (_32120_, _28076_, _32076_);
  and _45576_ (_32131_, _24445_, _28687_);
  nor _45577_ (_32142_, _24445_, _28687_);
  nor _45578_ (_32152_, _32142_, _32131_);
  not _45579_ (_32163_, _32152_);
  nand _45580_ (_32174_, _32163_, _25277_);
  and _45581_ (_32185_, _32174_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _45582_ (_32196_, _32131_, _29318_);
  and _45583_ (_32207_, _32142_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _45584_ (_32218_, _32207_, _32196_);
  and _45585_ (_32229_, _32218_, _25277_);
  or _45586_ (_32240_, _32229_, _32185_);
  and _45587_ (_32251_, _32240_, _28742_);
  or _45588_ (_32262_, _32251_, _32120_);
  or _45589_ (_32273_, _32262_, _32109_);
  and _45590_ (_08976_, _32273_, _41806_);
  and _45591_ (_32294_, _23824_, _21055_);
  not _45592_ (_32305_, _32294_);
  and _45593_ (_32326_, _20959_, _15702_);
  nor _45594_ (_32327_, _26942_, _26920_);
  not _45595_ (_32338_, _32327_);
  nor _45596_ (_32349_, _28153_, _26953_);
  and _45597_ (_32360_, _32349_, _32338_);
  not _45598_ (_32371_, _32360_);
  nor _45599_ (_32382_, _26539_, _25636_);
  nor _45600_ (_32393_, _32382_, _26550_);
  nor _45601_ (_32404_, _32393_, _25374_);
  nor _45602_ (_32415_, _26419_, _17247_);
  and _45603_ (_32425_, _26419_, _18520_);
  nor _45604_ (_32436_, _32425_, _32415_);
  nor _45605_ (_32447_, _32436_, _27356_);
  nor _45606_ (_32458_, _27117_, _27160_);
  nor _45607_ (_32469_, _27215_, _26419_);
  nor _45608_ (_32480_, _32469_, _32458_);
  and _45609_ (_32491_, _32480_, _18520_);
  nor _45610_ (_32502_, _32480_, _18520_);
  or _45611_ (_32513_, _32502_, _31012_);
  nor _45612_ (_32524_, _32513_, _32491_);
  nor _45613_ (_32535_, _32524_, _32447_);
  not _45614_ (_32546_, _27509_);
  and _45615_ (_32557_, _32546_, _27466_);
  nor _45616_ (_32568_, _27509_, _27455_);
  nor _45617_ (_32579_, _32568_, _17943_);
  nor _45618_ (_32590_, _32579_, _32557_);
  nor _45619_ (_32601_, _32590_, _27411_);
  nor _45620_ (_32612_, _27651_, _25495_);
  and _45621_ (_32633_, _27596_, _25506_);
  nor _45622_ (_32634_, _32633_, _32612_);
  and _45623_ (_32645_, _27618_, _25484_);
  and _45624_ (_32656_, _27672_, _17943_);
  nor _45625_ (_32667_, _32656_, _32645_);
  nor _45626_ (_32678_, _29079_, _16919_);
  not _45627_ (_32689_, _32678_);
  nor _45628_ (_32700_, _27814_, _17943_);
  nor _45629_ (_32711_, _27771_, _18107_);
  nor _45630_ (_32722_, _32711_, _32700_);
  and _45631_ (_32733_, _32722_, _32689_);
  and _45632_ (_32744_, _32733_, _32667_);
  and _45633_ (_32755_, _32744_, _32634_);
  not _45634_ (_32766_, _32755_);
  nor _45635_ (_32777_, _32766_, _32601_);
  and _45636_ (_32788_, _32777_, _32535_);
  not _45637_ (_32798_, _32788_);
  nor _45638_ (_32809_, _32798_, _32404_);
  and _45639_ (_32820_, _32809_, _32371_);
  not _45640_ (_32831_, _32820_);
  nor _45641_ (_32842_, _32831_, _32326_);
  and _45642_ (_32853_, _32842_, _32305_);
  not _45643_ (_32864_, _32853_);
  or _45644_ (_32875_, _32864_, _25287_);
  not _45645_ (_32886_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _45646_ (_32897_, _25287_, _32886_);
  and _45647_ (_32908_, _32897_, _28087_);
  and _45648_ (_32919_, _32908_, _32875_);
  nor _45649_ (_32930_, _28076_, _32886_);
  and _45650_ (_32941_, _29991_, _28687_);
  and _45651_ (_32952_, _32941_, _25277_);
  nand _45652_ (_32963_, _32952_, _28676_);
  or _45653_ (_32984_, _32952_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _45654_ (_32985_, _32984_, _28742_);
  and _45655_ (_32996_, _32985_, _32963_);
  or _45656_ (_33007_, _32996_, _32930_);
  or _45657_ (_33018_, _33007_, _32919_);
  and _45658_ (_08987_, _33018_, _41806_);
  and _45659_ (_33039_, _23889_, _21055_);
  not _45660_ (_33050_, _33039_);
  and _45661_ (_33061_, _20991_, _15702_);
  nor _45662_ (_33072_, _26975_, _26953_);
  not _45663_ (_33083_, _33072_);
  nor _45664_ (_33094_, _28153_, _26986_);
  and _45665_ (_33105_, _33094_, _33083_);
  not _45666_ (_33116_, _33105_);
  nor _45667_ (_33127_, _26550_, _25604_);
  nor _45668_ (_33138_, _33127_, _26561_);
  nor _45669_ (_33148_, _33138_, _25374_);
  nor _45670_ (_33159_, _26419_, _25408_);
  or _45671_ (_33170_, _33159_, _27356_);
  nor _45672_ (_33181_, _33170_, _28250_);
  nor _45673_ (_33192_, _26419_, _18520_);
  nand _45674_ (_33203_, _33192_, _27215_);
  nand _45675_ (_33214_, _27127_, _26419_);
  and _45676_ (_33225_, _33214_, _33203_);
  nor _45677_ (_33236_, _33225_, _16919_);
  not _45678_ (_33247_, _33236_);
  and _45679_ (_33258_, _33225_, _16919_);
  nor _45680_ (_33269_, _33258_, _31012_);
  and _45681_ (_33280_, _33269_, _33247_);
  nor _45682_ (_33291_, _33280_, _33181_);
  nor _45683_ (_33302_, _32557_, _16919_);
  and _45684_ (_33313_, _32557_, _16919_);
  nor _45685_ (_33324_, _33313_, _33302_);
  nor _45686_ (_33335_, _33324_, _27411_);
  and _45687_ (_33356_, _27596_, _25452_);
  nor _45688_ (_33357_, _27651_, _25441_);
  not _45689_ (_33368_, _33357_);
  and _45690_ (_33379_, _27618_, _25430_);
  and _45691_ (_33390_, _27672_, _16919_);
  nor _45692_ (_33401_, _33390_, _33379_);
  nand _45693_ (_33412_, _33401_, _33368_);
  nor _45694_ (_33423_, _33412_, _33356_);
  nor _45695_ (_33434_, _29079_, _17758_);
  not _45696_ (_33445_, _33434_);
  nor _45697_ (_33456_, _27814_, _16919_);
  nor _45698_ (_33467_, _27771_, _17943_);
  nor _45699_ (_33478_, _33467_, _33456_);
  and _45700_ (_33489_, _33478_, _33445_);
  and _45701_ (_33499_, _33489_, _33423_);
  not _45702_ (_33510_, _33499_);
  nor _45703_ (_33521_, _33510_, _33335_);
  and _45704_ (_33532_, _33521_, _33291_);
  not _45705_ (_33543_, _33532_);
  nor _45706_ (_33554_, _33543_, _33148_);
  and _45707_ (_33565_, _33554_, _33116_);
  not _45708_ (_33576_, _33565_);
  nor _45709_ (_33587_, _33576_, _33061_);
  and _45710_ (_33598_, _33587_, _33050_);
  not _45711_ (_33609_, _33598_);
  or _45712_ (_33620_, _33609_, _25287_);
  not _45713_ (_33631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _45714_ (_33642_, _25287_, _33631_);
  and _45715_ (_33653_, _33642_, _28087_);
  and _45716_ (_33664_, _33653_, _33620_);
  nor _45717_ (_33675_, _28076_, _33631_);
  nor _45718_ (_33686_, _24197_, _24313_);
  and _45719_ (_33697_, _33686_, _24434_);
  and _45720_ (_33708_, _33697_, _25277_);
  nand _45721_ (_33719_, _33708_, _28676_);
  or _45722_ (_33730_, _33708_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _45723_ (_33741_, _33730_, _28742_);
  and _45724_ (_33752_, _33741_, _33719_);
  or _45725_ (_33763_, _33752_, _33675_);
  or _45726_ (_33774_, _33763_, _33664_);
  and _45727_ (_08998_, _33774_, _41806_);
  and _45728_ (_33795_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45729_ (_33806_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor _45730_ (_33817_, _33806_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _45731_ (_33828_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _45732_ (_33839_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _45733_ (_33849_, _33839_, _33828_);
  and _45734_ (_33860_, _33806_, _15636_);
  and _45735_ (_33881_, _33860_, _33849_);
  not _45736_ (_33882_, _33881_);
  and _45737_ (_33893_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and _45738_ (_33904_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _45739_ (_33915_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _45740_ (_33926_, _33915_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _45741_ (_33937_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _45742_ (_33948_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _45743_ (_33959_, _33948_, _33937_);
  and _45744_ (_33970_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not _45745_ (_33981_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _45746_ (_33992_, _33981_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45747_ (_34003_, _33992_, _33937_);
  and _45748_ (_34014_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _45749_ (_34025_, _34014_, _33970_);
  and _45750_ (_34036_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45751_ (_34047_, _34036_, _33937_);
  and _45752_ (_34058_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not _45753_ (_34069_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45754_ (_34080_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _34069_);
  and _45755_ (_34091_, _34080_, _33937_);
  and _45756_ (_34102_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _45757_ (_34113_, _34102_, _34058_);
  and _45758_ (_34124_, _33948_, _33937_);
  and _45759_ (_34135_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and _45760_ (_34156_, _33948_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45761_ (_34157_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _45762_ (_34168_, _34157_, _34135_);
  and _45763_ (_34179_, _34168_, _34113_);
  and _45764_ (_34190_, _34179_, _34025_);
  nor _45765_ (_34200_, _34190_, _33926_);
  nor _45766_ (_34211_, _34200_, _33904_);
  nor _45767_ (_34222_, _34211_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45768_ (_34233_, _34222_, _33893_);
  nor _45769_ (_34244_, _34233_, _33882_);
  and _45770_ (_34255_, _33849_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _45771_ (_34266_, _34255_, _33882_);
  nor _45772_ (_34277_, _34266_, _34244_);
  and _45773_ (_34288_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45774_ (_34299_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _45775_ (_34310_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45776_ (_34321_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _45777_ (_34332_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _45778_ (_34343_, _34332_, _34321_);
  and _45779_ (_34354_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _45780_ (_34365_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _45781_ (_34376_, _34365_, _34354_);
  and _45782_ (_34387_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and _45783_ (_34398_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _45784_ (_34409_, _34398_, _34387_);
  and _45785_ (_34420_, _34409_, _34376_);
  and _45786_ (_34431_, _34420_, _34343_);
  nor _45787_ (_34442_, _34431_, _33915_);
  and _45788_ (_34453_, _34442_, _34310_);
  nor _45789_ (_34464_, _34453_, _34299_);
  nor _45790_ (_34475_, _34464_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45791_ (_34486_, _34475_, _34288_);
  nor _45792_ (_34497_, _34486_, _33882_);
  and _45793_ (_34508_, _33849_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _45794_ (_34519_, _34508_, _33882_);
  nor _45795_ (_34530_, _34519_, _34497_);
  not _45796_ (_34540_, _34530_);
  and _45797_ (_34551_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45798_ (_34562_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45799_ (_34573_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _45800_ (_34584_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _45801_ (_34595_, _34584_, _34573_);
  and _45802_ (_34606_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _45803_ (_34617_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _45804_ (_34628_, _34617_, _34606_);
  and _45805_ (_34639_, _34628_, _34595_);
  and _45806_ (_34650_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _45807_ (_34661_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _45808_ (_34672_, _34661_, _34650_);
  and _45809_ (_34683_, _34672_, _34639_);
  nor _45810_ (_34694_, _34683_, _33926_);
  nor _45811_ (_34705_, _34694_, _34562_);
  nor _45812_ (_34716_, _34705_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45813_ (_34727_, _34716_, _34551_);
  nor _45814_ (_34738_, _34727_, _33882_);
  and _45815_ (_34749_, _33849_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _45816_ (_34760_, _34749_, _33882_);
  nor _45817_ (_34781_, _34760_, _34738_);
  nor _45818_ (_34782_, _34781_, _34540_);
  and _45819_ (_34793_, _34782_, _34277_);
  and _45820_ (_34804_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not _45821_ (_34815_, _34804_);
  and _45822_ (_34826_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _45823_ (_34837_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _45824_ (_34848_, _34837_, _34826_);
  and _45825_ (_34859_, _34848_, _34815_);
  and _45826_ (_34870_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _45827_ (_34881_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _45828_ (_34891_, _34881_, _34870_);
  and _45829_ (_34902_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _45830_ (_34913_, _33915_, _34902_);
  and _45831_ (_34924_, _34913_, _34891_);
  and _45832_ (_34935_, _34924_, _34859_);
  and _45833_ (_34946_, _34935_, _34310_);
  nor _45834_ (_34957_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _34310_);
  nor _45835_ (_34968_, _34957_, _34946_);
  nor _45836_ (_34979_, _34968_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _45837_ (_34990_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45838_ (_35001_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _34990_);
  nor _45839_ (_35012_, _35001_, _34979_);
  and _45840_ (_35023_, _35012_, _33881_);
  and _45841_ (_35034_, _33849_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _45842_ (_35045_, _35034_, _33882_);
  nor _45843_ (_35056_, _35045_, _35023_);
  and _45844_ (_35067_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45845_ (_35078_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45846_ (_35089_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _45847_ (_35100_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _45848_ (_35111_, _35100_, _35089_);
  and _45849_ (_35122_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _45850_ (_35133_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _45851_ (_35144_, _35133_, _35122_);
  and _45852_ (_35155_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _45853_ (_35166_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _45854_ (_35177_, _35166_, _35155_);
  and _45855_ (_35188_, _35177_, _35144_);
  and _45856_ (_35199_, _35188_, _35111_);
  nor _45857_ (_35209_, _35199_, _33926_);
  nor _45858_ (_35220_, _35209_, _35078_);
  nor _45859_ (_35231_, _35220_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45860_ (_35242_, _35231_, _35067_);
  nor _45861_ (_35253_, _35242_, _33882_);
  and _45862_ (_35264_, _33849_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _45863_ (_35275_, _35264_, _33882_);
  nor _45864_ (_35286_, _35275_, _35253_);
  nor _45865_ (_35297_, _35286_, _35056_);
  and _45866_ (_35308_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45867_ (_35319_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45868_ (_35330_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and _45869_ (_35341_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _45870_ (_35352_, _35341_, _35330_);
  and _45871_ (_35363_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _45872_ (_35374_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _45873_ (_35385_, _35374_, _35363_);
  and _45874_ (_35396_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _45875_ (_35407_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _45876_ (_35418_, _35407_, _35396_);
  and _45877_ (_35429_, _35418_, _35385_);
  and _45878_ (_35440_, _35429_, _35352_);
  nor _45879_ (_35451_, _35440_, _33915_);
  and _45880_ (_35462_, _35451_, _34310_);
  or _45881_ (_35473_, _35462_, _35319_);
  and _45882_ (_35495_, _35473_, _34990_);
  nor _45883_ (_35496_, _35495_, _35308_);
  nor _45884_ (_35518_, _35496_, _33882_);
  and _45885_ (_35519_, _33849_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _45886_ (_35541_, _35519_, _33882_);
  nor _45887_ (_35542_, _35541_, _35518_);
  and _45888_ (_35563_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and _45889_ (_35564_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _45890_ (_35575_, _35564_, _35563_);
  and _45891_ (_35586_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _45892_ (_35597_, _35586_, _33915_);
  and _45893_ (_35608_, _35597_, _35575_);
  and _45894_ (_35619_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not _45895_ (_35630_, _35619_);
  and _45896_ (_35641_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _45897_ (_35652_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _45898_ (_35663_, _35652_, _35641_);
  and _45899_ (_35674_, _35663_, _35630_);
  and _45900_ (_35685_, _35674_, _35608_);
  and _45901_ (_35696_, _35685_, _34310_);
  nor _45902_ (_35707_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _34310_);
  or _45903_ (_35718_, _35707_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45904_ (_35729_, _35718_, _35696_);
  and _45905_ (_35740_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _45906_ (_35751_, _35740_, _35729_);
  and _45907_ (_35762_, _35751_, _33881_);
  and _45908_ (_35773_, _33849_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _45909_ (_35784_, _35773_, _33882_);
  nor _45910_ (_35795_, _35784_, _35762_);
  not _45911_ (_35806_, _35795_);
  and _45912_ (_35817_, _35806_, _35542_);
  and _45913_ (_35828_, _35817_, _35297_);
  and _45914_ (_35839_, _35828_, _34793_);
  and _45915_ (_35850_, _35297_, _35542_);
  and _45916_ (_35860_, _34781_, _34277_);
  and _45917_ (_35871_, _35860_, _34540_);
  and _45918_ (_35882_, _35871_, _35850_);
  or _45919_ (_35893_, _35882_, _35839_);
  not _45920_ (_35904_, _35893_);
  and _45921_ (_35915_, _35860_, _34530_);
  and _45922_ (_35926_, _35915_, _35850_);
  not _45923_ (_35937_, _34277_);
  and _45924_ (_35948_, _34781_, _35937_);
  and _45925_ (_35959_, _35948_, _34540_);
  and _45926_ (_35970_, _35959_, _35828_);
  nor _45927_ (_35981_, _35970_, _35926_);
  and _45928_ (_35992_, _35948_, _34530_);
  and _45929_ (_36003_, _35992_, _35806_);
  and _45930_ (_36014_, _36003_, _35850_);
  and _45931_ (_36025_, _34782_, _35937_);
  and _45932_ (_36036_, _36025_, _35850_);
  nor _45933_ (_36047_, _36036_, _36014_);
  and _45934_ (_36058_, _36047_, _35981_);
  and _45935_ (_36069_, _35795_, _35850_);
  nor _45936_ (_36080_, _34781_, _34530_);
  and _45937_ (_36091_, _36080_, _35937_);
  or _45938_ (_36102_, _36091_, _34793_);
  and _45939_ (_36113_, _36102_, _36069_);
  and _45940_ (_36124_, _35992_, _35795_);
  and _45941_ (_36135_, _36124_, _35850_);
  nor _45942_ (_36146_, _36135_, _36113_);
  and _45943_ (_36157_, _36146_, _36058_);
  and _45944_ (_36167_, _36157_, _35904_);
  and _45945_ (_36178_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45946_ (_36189_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45947_ (_36200_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _45948_ (_36211_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _45949_ (_36222_, _36211_, _36200_);
  and _45950_ (_36233_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _45951_ (_36244_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _45952_ (_36255_, _36244_, _36233_);
  and _45953_ (_36266_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _45954_ (_36277_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _45955_ (_36288_, _36277_, _36266_);
  and _45956_ (_36299_, _36288_, _36255_);
  and _45957_ (_36310_, _36299_, _36222_);
  nor _45958_ (_36321_, _36310_, _33915_);
  and _45959_ (_36332_, _36321_, _34310_);
  nor _45960_ (_36343_, _36332_, _36189_);
  nor _45961_ (_36354_, _36343_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45962_ (_36365_, _36354_, _36178_);
  nor _45963_ (_36376_, _36365_, _33882_);
  and _45964_ (_36387_, _33849_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _45965_ (_36398_, _36387_, _33882_);
  nor _45966_ (_36409_, _36398_, _36376_);
  not _45967_ (_36420_, _36409_);
  not _45968_ (_36431_, _35056_);
  and _45969_ (_36442_, _35542_, _35286_);
  and _45970_ (_36453_, _36442_, _36431_);
  and _45971_ (_36464_, _36453_, _36420_);
  and _45972_ (_36474_, _35959_, _35795_);
  and _45973_ (_36485_, _36474_, _36464_);
  and _45974_ (_36496_, _36464_, _36003_);
  and _45975_ (_36507_, _36080_, _34277_);
  and _45976_ (_36518_, _36507_, _35806_);
  and _45977_ (_36529_, _36518_, _36464_);
  nor _45978_ (_36540_, _36529_, _36496_);
  not _45979_ (_36551_, _36540_);
  nor _45980_ (_36562_, _36551_, _36485_);
  and _45981_ (_36573_, _36409_, _35056_);
  and _45982_ (_36584_, _36573_, _36442_);
  and _45983_ (_36595_, _36025_, _35806_);
  and _45984_ (_36606_, _36595_, _36584_);
  not _45985_ (_36617_, _36606_);
  and _45986_ (_36628_, _36453_, _36409_);
  and _45987_ (_36639_, _36628_, _35871_);
  and _45988_ (_36650_, _36507_, _35795_);
  and _45989_ (_36661_, _36650_, _35850_);
  nor _45990_ (_36672_, _36661_, _36639_);
  and _45991_ (_36683_, _36672_, _36617_);
  and _45992_ (_36694_, _36683_, _36562_);
  and _45993_ (_36705_, _36694_, _36167_);
  nor _45994_ (_36716_, _36705_, _33817_);
  not _45995_ (_36727_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _45996_ (_36738_, _15636_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _45997_ (_36749_, _36738_, _36727_);
  and _45998_ (_36760_, _36749_, _36507_);
  and _45999_ (_36771_, _36760_, _36584_);
  and _46000_ (_36781_, _36639_, _36738_);
  and _46001_ (_36792_, _36781_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or _46002_ (_36803_, _36792_, _36771_);
  nor _46003_ (_36814_, _36803_, _36716_);
  nor _46004_ (_36825_, _36814_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46005_ (_36836_, _36825_, _33795_);
  and _46006_ (_36847_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _46007_ (_36858_, _33817_);
  not _46008_ (_36869_, _35286_);
  and _46009_ (_36880_, _35542_, _36869_);
  nor _46010_ (_36891_, _36409_, _36431_);
  and _46011_ (_36902_, _36891_, _36880_);
  and _46012_ (_36913_, _35948_, _35806_);
  and _46013_ (_36924_, _36913_, _36902_);
  and _46014_ (_36935_, _36091_, _35795_);
  and _46015_ (_36946_, _36935_, _36902_);
  and _46016_ (_36957_, _35959_, _36069_);
  or _46017_ (_36968_, _36957_, _36946_);
  or _46018_ (_36979_, _36968_, _36924_);
  and _46019_ (_36990_, _34793_, _35806_);
  or _46020_ (_37001_, _36990_, _35871_);
  and _46021_ (_37012_, _36902_, _37001_);
  nor _46022_ (_37023_, _35806_, _35542_);
  and _46023_ (_37034_, _37023_, _35959_);
  and _46024_ (_37045_, _35915_, _35795_);
  and _46025_ (_37056_, _37045_, _36902_);
  or _46026_ (_37067_, _37056_, _37034_);
  or _46027_ (_37078_, _37067_, _36639_);
  or _46028_ (_37087_, _37078_, _37012_);
  and _46029_ (_37095_, _36902_, _36650_);
  and _46030_ (_37102_, _36025_, _35795_);
  and _46031_ (_37110_, _37102_, _36902_);
  or _46032_ (_37118_, _37110_, _37095_);
  and _46033_ (_37125_, _36628_, _36474_);
  and _46034_ (_37133_, _36628_, _36595_);
  nor _46035_ (_37141_, _37133_, _37125_);
  not _46036_ (_37148_, _37141_);
  or _46037_ (_37149_, _37148_, _37118_);
  or _46038_ (_37150_, _37149_, _37087_);
  or _46039_ (_37153_, _37150_, _36979_);
  and _46040_ (_37164_, _34793_, _35795_);
  and _46041_ (_37175_, _37164_, _36453_);
  and _46042_ (_37186_, _35915_, _35806_);
  and _46043_ (_37197_, _37186_, _36902_);
  and _46044_ (_37208_, _35959_, _35806_);
  and _46045_ (_37219_, _36584_, _37208_);
  or _46046_ (_37230_, _37219_, _37197_);
  nor _46047_ (_37241_, _37230_, _37175_);
  and _46048_ (_37252_, _36628_, _36518_);
  and _46049_ (_37263_, _36902_, _36595_);
  nor _46050_ (_37274_, _37263_, _37252_);
  and _46051_ (_37285_, _37274_, _37241_);
  and _46052_ (_37296_, _36584_, _36474_);
  and _46053_ (_37307_, _37164_, _36902_);
  nor _46054_ (_37318_, _37307_, _37296_);
  and _46055_ (_37329_, _36628_, _37208_);
  and _46056_ (_37340_, _37102_, _36628_);
  nor _46057_ (_37351_, _37340_, _37329_);
  and _46058_ (_37362_, _37351_, _37318_);
  and _46059_ (_37373_, _37362_, _37285_);
  and _46060_ (_37384_, _36628_, _36003_);
  and _46061_ (_37394_, _36902_, _36124_);
  or _46062_ (_37405_, _37394_, _37384_);
  and _46063_ (_37416_, _36584_, _36025_);
  and _46064_ (_37421_, _36650_, _36453_);
  or _46065_ (_37432_, _37421_, _37416_);
  or _46066_ (_37443_, _37432_, _37405_);
  and _46067_ (_37454_, _36628_, _36124_);
  and _46068_ (_37464_, _36453_, _36990_);
  or _46069_ (_37475_, _37464_, _37454_);
  and _46070_ (_37485_, _36584_, _35871_);
  and _46071_ (_37496_, _37485_, _35795_);
  and _46072_ (_37507_, _35806_, _35871_);
  or _46073_ (_37518_, _37186_, _37507_);
  and _46074_ (_37528_, _37518_, _36584_);
  nor _46075_ (_37539_, _37528_, _37496_);
  not _46076_ (_37550_, _37539_);
  or _46077_ (_37560_, _37550_, _37475_);
  nor _46078_ (_37571_, _37560_, _37443_);
  nand _46079_ (_37582_, _37571_, _37373_);
  or _46080_ (_37592_, _37582_, _37153_);
  and _46081_ (_37603_, _37592_, _36858_);
  and _46082_ (_37614_, _36738_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _46083_ (_37624_, _37614_, _36639_);
  not _46084_ (_37635_, _37624_);
  nor _46085_ (_37646_, _34781_, _35937_);
  and _46086_ (_37657_, _36584_, _37646_);
  and _46087_ (_37668_, _37657_, _36749_);
  not _46088_ (_37679_, _36749_);
  and _46089_ (_37690_, _35795_, _35871_);
  and _46090_ (_37701_, _37690_, _36584_);
  and _46091_ (_37712_, _37186_, _36584_);
  nor _46092_ (_37723_, _37712_, _37701_);
  nor _46093_ (_37734_, _37723_, _37679_);
  nor _46094_ (_37745_, _37734_, _37668_);
  and _46095_ (_37756_, _37745_, _37635_);
  not _46096_ (_37767_, _37756_);
  nor _46097_ (_37778_, _37767_, _37603_);
  nor _46098_ (_37789_, _37778_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46099_ (_37800_, _37789_, _36847_);
  nor _46100_ (_37811_, _37800_, _36836_);
  and _46101_ (_37822_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _46102_ (_37833_, _36573_, _36880_);
  and _46103_ (_37844_, _37833_, _36124_);
  and _46104_ (_37855_, _37833_, _36474_);
  nor _46105_ (_37866_, _37855_, _37844_);
  and _46106_ (_37877_, _37866_, _36562_);
  nor _46107_ (_37888_, _37877_, _33817_);
  nor _46108_ (_37899_, _37888_, _37668_);
  nor _46109_ (_37910_, _37866_, _36858_);
  not _46110_ (_37921_, _37910_);
  and _46111_ (_37932_, _37921_, _37899_);
  nor _46112_ (_37943_, _37932_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46113_ (_37954_, _37943_, _37822_);
  and _46114_ (_37965_, _37954_, _41806_);
  and _46115_ (_09544_, _37965_, _37811_);
  and _46116_ (_37986_, _24796_, _24665_);
  and _46117_ (_37997_, _37986_, _25244_);
  and _46118_ (_38008_, _37997_, _24960_);
  and _46119_ (_38019_, _38008_, _25112_);
  and _46120_ (_38030_, _38019_, _30002_);
  and _46121_ (_38041_, _38030_, _28076_);
  and _46122_ (_38052_, _38041_, _28044_);
  nor _46123_ (_38063_, _21055_, _15702_);
  and _46124_ (_38074_, _26648_, _21034_);
  nor _46125_ (_38085_, _27813_, _38074_);
  and _46126_ (_38096_, _38085_, _27771_);
  and _46127_ (_38107_, _38096_, _38063_);
  and _46128_ (_38118_, _38107_, _29079_);
  nor _46129_ (_38129_, _38118_, _17758_);
  not _46130_ (_38140_, _38129_);
  and _46131_ (_38151_, _38140_, _27716_);
  and _46132_ (_38162_, _38151_, _27389_);
  not _46133_ (_38173_, _38162_);
  and _46134_ (_38183_, _38173_, _38052_);
  and _46135_ (_38194_, _38019_, _24197_);
  and _46136_ (_38205_, _38194_, _29991_);
  and _46137_ (_38216_, _38205_, _28087_);
  not _46138_ (_38226_, _38216_);
  and _46139_ (_38237_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _46140_ (_38248_, _38118_, _16919_);
  not _46141_ (_38258_, _38248_);
  and _46142_ (_38269_, _38258_, _33423_);
  and _46143_ (_38280_, _38269_, _33291_);
  nor _46144_ (_38290_, _38280_, _38226_);
  nor _46145_ (_38301_, _38290_, _38237_);
  and _46146_ (_38312_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _46147_ (_38322_, _38118_, _17943_);
  not _46148_ (_38333_, _38322_);
  and _46149_ (_38344_, _38333_, _32667_);
  and _46150_ (_38355_, _38344_, _32634_);
  and _46151_ (_38366_, _38355_, _32535_);
  nor _46152_ (_38377_, _38366_, _38226_);
  nor _46153_ (_38388_, _38377_, _38312_);
  and _46154_ (_38390_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _46155_ (_38391_, _38118_, _18107_);
  not _46156_ (_38392_, _38391_);
  and _46157_ (_38393_, _38392_, _31913_);
  and _46158_ (_38394_, _38393_, _31794_);
  nor _46159_ (_38395_, _38394_, _38226_);
  nor _46160_ (_38396_, _38395_, _38390_);
  and _46161_ (_38397_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _46162_ (_38398_, _38118_, _18477_);
  not _46163_ (_38399_, _38398_);
  and _46164_ (_38400_, _38399_, _31207_);
  and _46165_ (_38401_, _38400_, _31175_);
  and _46166_ (_38402_, _38401_, _31055_);
  nor _46167_ (_38403_, _38402_, _38226_);
  nor _46168_ (_38404_, _38403_, _38397_);
  and _46169_ (_38405_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _46170_ (_38406_, _38118_, _18978_);
  not _46171_ (_38407_, _38406_);
  and _46172_ (_38408_, _38407_, _30306_);
  and _46173_ (_38409_, _38408_, _30338_);
  and _46174_ (_38410_, _38409_, _30219_);
  nor _46175_ (_38411_, _38410_, _38226_);
  nor _46176_ (_38412_, _38411_, _38405_);
  and _46177_ (_38413_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _46178_ (_38414_, _38118_, _18815_);
  not _46179_ (_38415_, _38414_);
  and _46180_ (_38416_, _38415_, _29654_);
  and _46181_ (_38417_, _38416_, _29839_);
  not _46182_ (_38418_, _38417_);
  and _46183_ (_38419_, _38418_, _38216_);
  nor _46184_ (_38420_, _38419_, _38413_);
  nor _46185_ (_38421_, _38216_, _24379_);
  nor _46186_ (_38422_, _38118_, _19360_);
  not _46187_ (_38423_, _38422_);
  and _46188_ (_38424_, _38423_, _29057_);
  and _46189_ (_38425_, _38424_, _29002_);
  not _46190_ (_38426_, _38425_);
  and _46191_ (_38427_, _38426_, _38216_);
  nor _46192_ (_38428_, _38427_, _38421_);
  and _46193_ (_38429_, _38428_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46194_ (_38430_, _38429_, _38420_);
  and _46195_ (_38431_, _38430_, _38412_);
  and _46196_ (_38432_, _38431_, _38404_);
  and _46197_ (_38433_, _38432_, _38396_);
  and _46198_ (_38434_, _38433_, _38388_);
  and _46199_ (_38435_, _38434_, _38301_);
  nor _46200_ (_38436_, _38216_, _24818_);
  and _46201_ (_38437_, _38436_, _38435_);
  nor _46202_ (_38438_, _38436_, _38435_);
  nor _46203_ (_38439_, _38438_, _38437_);
  and _46204_ (_38440_, _38439_, _24522_);
  nor _46205_ (_38441_, _38440_, _24862_);
  nor _46206_ (_38442_, _38441_, _38216_);
  nor _46207_ (_38443_, _38442_, _38183_);
  nor _46208_ (_09564_, _38443_, rst);
  not _46209_ (_38444_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46210_ (_38445_, _38428_, _38444_);
  nor _46211_ (_38446_, _38428_, _38444_);
  nor _46212_ (_38447_, _38446_, _38445_);
  and _46213_ (_38448_, _38447_, _24522_);
  nor _46214_ (_38449_, _38448_, _24390_);
  nor _46215_ (_38450_, _38449_, _38216_);
  nor _46216_ (_38451_, _38450_, _38427_);
  nand _46217_ (_10690_, _38451_, _41806_);
  nor _46218_ (_38452_, _38429_, _38420_);
  nor _46219_ (_38453_, _38452_, _38430_);
  nor _46220_ (_38454_, _38453_, _23943_);
  nor _46221_ (_38455_, _38454_, _24245_);
  nor _46222_ (_38456_, _38455_, _38216_);
  nor _46223_ (_38457_, _38456_, _38419_);
  nand _46224_ (_10701_, _38457_, _41806_);
  nor _46225_ (_38458_, _38430_, _38412_);
  nor _46226_ (_38459_, _38458_, _38431_);
  nor _46227_ (_38460_, _38459_, _23943_);
  nor _46228_ (_38461_, _38460_, _23998_);
  nor _46229_ (_38462_, _38461_, _38216_);
  nor _46230_ (_38463_, _38462_, _38411_);
  nand _46231_ (_10712_, _38463_, _41806_);
  nor _46232_ (_38464_, _38431_, _38404_);
  nor _46233_ (_38465_, _38464_, _38432_);
  nor _46234_ (_38466_, _38465_, _23943_);
  nor _46235_ (_38467_, _38466_, _25004_);
  nor _46236_ (_38468_, _38467_, _38216_);
  nor _46237_ (_38469_, _38468_, _38403_);
  nor _46238_ (_10723_, _38469_, rst);
  nor _46239_ (_38470_, _38432_, _38396_);
  nor _46240_ (_38471_, _38470_, _38433_);
  nor _46241_ (_38472_, _38471_, _23943_);
  nor _46242_ (_38473_, _38472_, _25156_);
  nor _46243_ (_38474_, _38473_, _38216_);
  nor _46244_ (_38475_, _38474_, _38395_);
  nor _46245_ (_10734_, _38475_, rst);
  nor _46246_ (_38476_, _38433_, _38388_);
  nor _46247_ (_38477_, _38476_, _38434_);
  nor _46248_ (_38478_, _38477_, _23943_);
  nor _46249_ (_38479_, _38478_, _24708_);
  nor _46250_ (_38480_, _38479_, _38216_);
  nor _46251_ (_38481_, _38480_, _38377_);
  nor _46252_ (_10745_, _38481_, rst);
  nor _46253_ (_38482_, _38434_, _38301_);
  nor _46254_ (_38483_, _38482_, _38435_);
  nor _46255_ (_38484_, _38483_, _23943_);
  nor _46256_ (_38485_, _38484_, _24555_);
  nor _46257_ (_38486_, _38485_, _38216_);
  nor _46258_ (_38487_, _38486_, _38290_);
  nor _46259_ (_10756_, _38487_, rst);
  and _46260_ (_38488_, _28087_, _25112_);
  and _46261_ (_38489_, _38488_, _31436_);
  nand _46262_ (_38490_, _38489_, _38008_);
  nor _46263_ (_38491_, _38490_, _28011_);
  and _46264_ (_38492_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15636_);
  and _46265_ (_38493_, _38492_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46266_ (_38494_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _46267_ (_38495_, _38494_, _38493_);
  or _46268_ (_38496_, _38495_, _38491_);
  nor _46269_ (_38497_, _27814_, _17584_);
  nor _46270_ (_38498_, _28436_, _18477_);
  and _46271_ (_38499_, _26419_, _17247_);
  not _46272_ (_38500_, _38499_);
  nor _46273_ (_38501_, _17758_, _16425_);
  and _46274_ (_38502_, _38501_, _27138_);
  and _46275_ (_38503_, _38502_, _25821_);
  and _46276_ (_38504_, _38503_, _25865_);
  and _46277_ (_38505_, _38504_, _26474_);
  nor _46278_ (_38506_, _38505_, _27160_);
  and _46279_ (_38507_, _26419_, _16260_);
  nor _46280_ (_38508_, _38507_, _38506_);
  and _46281_ (_38509_, _38508_, _38500_);
  and _46282_ (_38510_, _27226_, _17758_);
  and _46283_ (_38511_, _17094_, _16096_);
  and _46284_ (_38512_, _17410_, _16425_);
  and _46285_ (_38513_, _38512_, _38511_);
  and _46286_ (_38514_, _38513_, _38510_);
  and _46287_ (_38515_, _17247_, _16260_);
  and _46288_ (_38516_, _38515_, _38514_);
  nor _46289_ (_38517_, _38516_, _26419_);
  not _46290_ (_38518_, _38517_);
  and _46291_ (_38519_, _38518_, _38509_);
  nor _46292_ (_38520_, _26419_, _16601_);
  and _46293_ (_38521_, _26419_, _16601_);
  nor _46294_ (_38522_, _38521_, _38520_);
  and _46295_ (_38523_, _38522_, _38519_);
  nor _46296_ (_38524_, _38523_, _27302_);
  and _46297_ (_38525_, _38523_, _27302_);
  nor _46298_ (_38526_, _38525_, _38524_);
  and _46299_ (_38527_, _38526_, _27073_);
  and _46300_ (_38528_, _26419_, _27302_);
  nor _46301_ (_38529_, _38528_, _28273_);
  nor _46302_ (_38530_, _38529_, _27356_);
  or _46303_ (_38531_, _38530_, _38527_);
  or _46304_ (_38532_, _38531_, _38498_);
  and _46305_ (_38533_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor _46306_ (_38534_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _46307_ (_38535_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _46308_ (_38536_, _38535_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46309_ (_38537_, _38536_, _38534_);
  nor _46310_ (_38538_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _46311_ (_38539_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _46312_ (_38540_, _38539_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46313_ (_38541_, _38540_, _38538_);
  nor _46314_ (_38542_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _46315_ (_38543_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _46316_ (_38544_, _38543_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46317_ (_38545_, _38544_, _38542_);
  not _46318_ (_38546_, _38545_);
  nor _46319_ (_38547_, _38546_, _28175_);
  nor _46320_ (_38548_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _46321_ (_38549_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _46322_ (_38550_, _38549_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46323_ (_38551_, _38550_, _38548_);
  and _46324_ (_38552_, _38551_, _38547_);
  nor _46325_ (_38553_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _46326_ (_38554_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _46327_ (_38555_, _38554_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46328_ (_38556_, _38555_, _38553_);
  and _46329_ (_38557_, _38556_, _38552_);
  and _46330_ (_38558_, _38557_, _38541_);
  nor _46331_ (_38559_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _46332_ (_38560_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _46333_ (_38561_, _38560_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46334_ (_38562_, _38561_, _38559_);
  and _46335_ (_38563_, _38562_, _38558_);
  and _46336_ (_38564_, _38563_, _38537_);
  nor _46337_ (_38565_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _46338_ (_38566_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _46339_ (_38567_, _38566_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46340_ (_38568_, _38567_, _38565_);
  and _46341_ (_38569_, _38568_, _38564_);
  nor _46342_ (_38570_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _46343_ (_38571_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _46344_ (_38572_, _38571_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46345_ (_38573_, _38572_, _38570_);
  nor _46346_ (_38574_, _38573_, _38569_);
  and _46347_ (_38575_, _38573_, _38569_);
  or _46348_ (_38576_, _38575_, _38574_);
  nor _46349_ (_38577_, _38576_, _28153_);
  and _46350_ (_38578_, _20747_, _15702_);
  or _46351_ (_38579_, _38578_, _38577_);
  or _46352_ (_38580_, _38579_, _38533_);
  or _46353_ (_38581_, _38580_, _38532_);
  nor _46354_ (_38582_, _38581_, _38497_);
  nand _46355_ (_38583_, _38582_, _38493_);
  and _46356_ (_38584_, _38583_, _41806_);
  and _46357_ (_12702_, _38584_, _38496_);
  and _46358_ (_38585_, _38488_, _30708_);
  and _46359_ (_38586_, _38585_, _38008_);
  nor _46360_ (_38587_, _38586_, _38493_);
  not _46361_ (_38588_, _38587_);
  nand _46362_ (_38589_, _38588_, _28011_);
  not _46363_ (_38590_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand _46364_ (_38591_, _38587_, _38590_);
  and _46365_ (_38592_, _38591_, _41806_);
  and _46366_ (_12723_, _38592_, _38589_);
  nor _46367_ (_38593_, _38490_, _29231_);
  and _46368_ (_38594_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _46369_ (_38595_, _38594_, _38493_);
  or _46370_ (_38596_, _38595_, _38593_);
  nor _46371_ (_38597_, _27814_, _16425_);
  nor _46372_ (_38598_, _28436_, _18107_);
  nor _46373_ (_38599_, _27356_, _19360_);
  nor _46374_ (_38600_, _28273_, _27335_);
  not _46375_ (_38601_, _38600_);
  nor _46376_ (_38602_, _38601_, _27247_);
  nor _46377_ (_38603_, _38602_, _25789_);
  and _46378_ (_38604_, _38602_, _25789_);
  nor _46379_ (_38605_, _38604_, _38603_);
  and _46380_ (_38606_, _38605_, _27073_);
  or _46381_ (_38607_, _38606_, _38599_);
  or _46382_ (_38608_, _38607_, _38598_);
  and _46383_ (_38609_, _23373_, _21055_);
  and _46384_ (_38610_, _38546_, _28175_);
  nor _46385_ (_38611_, _38610_, _38547_);
  and _46386_ (_38612_, _38611_, _26659_);
  and _46387_ (_38613_, _20525_, _15702_);
  or _46388_ (_38614_, _38613_, _38612_);
  or _46389_ (_38615_, _38614_, _38609_);
  or _46390_ (_38616_, _38615_, _38608_);
  nor _46391_ (_38617_, _38616_, _38597_);
  nand _46392_ (_38618_, _38617_, _38493_);
  and _46393_ (_38619_, _38618_, _41806_);
  and _46394_ (_13612_, _38619_, _38596_);
  nor _46395_ (_38620_, _38490_, _29893_);
  and _46396_ (_38621_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _46397_ (_38622_, _38621_, _38493_);
  or _46398_ (_38623_, _38622_, _38620_);
  nor _46399_ (_38624_, _27814_, _17410_);
  nor _46400_ (_38625_, _28436_, _17943_);
  and _46401_ (_38626_, _38502_, _26419_);
  and _46402_ (_38627_, _38510_, _16425_);
  and _46403_ (_38628_, _38627_, _27160_);
  nor _46404_ (_38629_, _38628_, _38626_);
  and _46405_ (_38630_, _38629_, _17410_);
  nor _46406_ (_38631_, _38629_, _17410_);
  or _46407_ (_38632_, _38631_, _31012_);
  nor _46408_ (_38633_, _38632_, _38630_);
  nor _46409_ (_38634_, _27356_, _18815_);
  or _46410_ (_38635_, _38634_, _38633_);
  or _46411_ (_38636_, _38635_, _38625_);
  and _46412_ (_38637_, _22369_, _21055_);
  nor _46413_ (_38638_, _38551_, _38547_);
  nor _46414_ (_38639_, _38638_, _38552_);
  and _46415_ (_38640_, _38639_, _26659_);
  and _46416_ (_38641_, _20557_, _15702_);
  or _46417_ (_38642_, _38641_, _38640_);
  or _46418_ (_38643_, _38642_, _38637_);
  or _46419_ (_38644_, _38643_, _38636_);
  nor _46420_ (_38645_, _38644_, _38624_);
  nand _46421_ (_38646_, _38645_, _38493_);
  and _46422_ (_38647_, _38646_, _41806_);
  and _46423_ (_13621_, _38647_, _38623_);
  nor _46424_ (_38648_, _38490_, _30567_);
  and _46425_ (_38649_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _46426_ (_38650_, _38649_, _38493_);
  or _46427_ (_38651_, _38650_, _38648_);
  nor _46428_ (_38652_, _27814_, _16096_);
  nor _46429_ (_38653_, _28436_, _16919_);
  and _46430_ (_38654_, _38627_, _17410_);
  and _46431_ (_38655_, _38654_, _27160_);
  and _46432_ (_38656_, _38503_, _26419_);
  nor _46433_ (_38657_, _38656_, _38655_);
  and _46434_ (_38658_, _38657_, _16096_);
  nor _46435_ (_38659_, _38657_, _16096_);
  nor _46436_ (_38660_, _38659_, _38658_);
  and _46437_ (_38661_, _38660_, _27073_);
  nor _46438_ (_38662_, _27356_, _18978_);
  or _46439_ (_38663_, _38662_, _38661_);
  or _46440_ (_38664_, _38663_, _38653_);
  and _46441_ (_38665_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _46442_ (_38666_, _38556_, _38552_);
  nor _46443_ (_38667_, _38666_, _38557_);
  and _46444_ (_38668_, _38667_, _26659_);
  and _46445_ (_38669_, _20589_, _15702_);
  or _46446_ (_38670_, _38669_, _38668_);
  or _46447_ (_38671_, _38670_, _38665_);
  or _46448_ (_38672_, _38671_, _38664_);
  nor _46449_ (_38673_, _38672_, _38652_);
  nand _46450_ (_38674_, _38673_, _38493_);
  and _46451_ (_38675_, _38674_, _41806_);
  and _46452_ (_13631_, _38675_, _38651_);
  nor _46453_ (_38676_, _38490_, _31338_);
  and _46454_ (_38677_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _46455_ (_38678_, _38677_, _38493_);
  or _46456_ (_38679_, _38678_, _38676_);
  nor _46457_ (_38680_, _27814_, _17094_);
  nor _46458_ (_38681_, _38504_, _26474_);
  not _46459_ (_38682_, _38681_);
  and _46460_ (_38683_, _38682_, _38506_);
  and _46461_ (_38684_, _38654_, _16096_);
  nor _46462_ (_38685_, _38684_, _17094_);
  nor _46463_ (_38686_, _38685_, _38514_);
  nor _46464_ (_38687_, _38686_, _26419_);
  nor _46465_ (_38688_, _38687_, _38683_);
  nor _46466_ (_38689_, _38688_, _31012_);
  nor _46467_ (_38690_, _27356_, _18477_);
  or _46468_ (_38691_, _38690_, _38689_);
  or _46469_ (_38692_, _38691_, _28447_);
  and _46470_ (_38693_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _46471_ (_38694_, _38557_, _38541_);
  not _46472_ (_38695_, _38694_);
  nor _46473_ (_38696_, _38558_, _28153_);
  and _46474_ (_38697_, _38696_, _38695_);
  and _46475_ (_38698_, _20620_, _15702_);
  or _46476_ (_38699_, _38698_, _38697_);
  or _46477_ (_38700_, _38699_, _38693_);
  or _46478_ (_38701_, _38700_, _38692_);
  nor _46479_ (_38702_, _38701_, _38680_);
  nand _46480_ (_38703_, _38702_, _38493_);
  and _46481_ (_38704_, _38703_, _41806_);
  and _46482_ (_13640_, _38704_, _38679_);
  nor _46483_ (_38705_, _38490_, _32044_);
  and _46484_ (_38706_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _46485_ (_38707_, _38706_, _38493_);
  or _46486_ (_38708_, _38707_, _38705_);
  nor _46487_ (_38709_, _27814_, _16260_);
  nor _46488_ (_38710_, _28436_, _19360_);
  nor _46489_ (_38711_, _38514_, _26419_);
  nor _46490_ (_38712_, _38711_, _38506_);
  nor _46491_ (_38713_, _38712_, _25517_);
  and _46492_ (_38714_, _38712_, _25517_);
  nor _46493_ (_38715_, _38714_, _38713_);
  and _46494_ (_38716_, _38715_, _27073_);
  nor _46495_ (_38717_, _26419_, _18117_);
  or _46496_ (_38718_, _38717_, _27356_);
  nor _46497_ (_38719_, _38718_, _38507_);
  or _46498_ (_38720_, _38719_, _38716_);
  or _46499_ (_38721_, _38720_, _38710_);
  and _46500_ (_38722_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _46501_ (_38723_, _38562_, _38558_);
  not _46502_ (_38724_, _38723_);
  nor _46503_ (_38725_, _38563_, _28153_);
  and _46504_ (_38726_, _38725_, _38724_);
  and _46505_ (_38727_, _20652_, _15702_);
  or _46506_ (_38728_, _38727_, _38726_);
  or _46507_ (_38729_, _38728_, _38722_);
  or _46508_ (_38730_, _38729_, _38721_);
  nor _46509_ (_38731_, _38730_, _38709_);
  nand _46510_ (_38732_, _38731_, _38493_);
  and _46511_ (_38733_, _38732_, _41806_);
  and _46512_ (_13650_, _38733_, _38708_);
  nor _46513_ (_38734_, _38490_, _32853_);
  and _46514_ (_38735_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _46515_ (_38736_, _38735_, _38493_);
  or _46516_ (_38737_, _38736_, _38734_);
  nor _46517_ (_38738_, _27814_, _17247_);
  nor _46518_ (_38739_, _28436_, _18815_);
  and _46519_ (_38740_, _38514_, _16260_);
  nor _46520_ (_38741_, _38740_, _26419_);
  not _46521_ (_38742_, _38741_);
  and _46522_ (_38743_, _38742_, _38508_);
  and _46523_ (_38744_, _38743_, _17247_);
  nor _46524_ (_38745_, _38743_, _17247_);
  or _46525_ (_38746_, _38745_, _38744_);
  and _46526_ (_38747_, _38746_, _27073_);
  nor _46527_ (_38748_, _33192_, _27356_);
  and _46528_ (_38749_, _38748_, _38500_);
  or _46529_ (_38750_, _38749_, _38747_);
  or _46530_ (_38751_, _38750_, _38739_);
  and _46531_ (_38752_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _46532_ (_38753_, _38563_, _38537_);
  nor _46533_ (_38754_, _38753_, _38564_);
  and _46534_ (_38755_, _38754_, _26659_);
  and _46535_ (_38756_, _20684_, _15702_);
  or _46536_ (_38757_, _38756_, _38755_);
  or _46537_ (_38758_, _38757_, _38752_);
  or _46538_ (_38759_, _38758_, _38751_);
  nor _46539_ (_38760_, _38759_, _38738_);
  nand _46540_ (_38761_, _38760_, _38493_);
  and _46541_ (_38762_, _38761_, _41806_);
  and _46542_ (_13660_, _38762_, _38737_);
  nor _46543_ (_38763_, _38490_, _33598_);
  and _46544_ (_38764_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _46545_ (_38765_, _38764_, _38493_);
  or _46546_ (_38766_, _38765_, _38763_);
  nor _46547_ (_38767_, _27814_, _16601_);
  nor _46548_ (_38768_, _28436_, _18978_);
  and _46549_ (_38769_, _38519_, _16601_);
  nor _46550_ (_38770_, _38519_, _16601_);
  nor _46551_ (_38771_, _38770_, _38769_);
  nor _46552_ (_38772_, _38771_, _31012_);
  nor _46553_ (_38773_, _26419_, _16930_);
  or _46554_ (_38774_, _38773_, _27356_);
  nor _46555_ (_38775_, _38774_, _38521_);
  or _46556_ (_38776_, _38775_, _38772_);
  or _46557_ (_38777_, _38776_, _38768_);
  and _46558_ (_38778_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _46559_ (_38779_, _38568_, _38564_);
  not _46560_ (_38780_, _38779_);
  nor _46561_ (_38781_, _38569_, _28153_);
  and _46562_ (_38782_, _38781_, _38780_);
  and _46563_ (_38783_, _20715_, _15702_);
  or _46564_ (_38784_, _38783_, _38782_);
  or _46565_ (_38785_, _38784_, _38778_);
  or _46566_ (_38786_, _38785_, _38777_);
  nor _46567_ (_38787_, _38786_, _38767_);
  nand _46568_ (_38788_, _38787_, _38493_);
  and _46569_ (_38789_, _38788_, _41806_);
  and _46570_ (_13670_, _38789_, _38766_);
  nand _46571_ (_38790_, _38588_, _29231_);
  not _46572_ (_38791_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _46573_ (_38792_, _38587_, _38791_);
  and _46574_ (_38793_, _38792_, _41806_);
  and _46575_ (_13679_, _38793_, _38790_);
  nand _46576_ (_38794_, _38588_, _29893_);
  not _46577_ (_38795_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand _46578_ (_38796_, _38587_, _38795_);
  and _46579_ (_38797_, _38796_, _41806_);
  and _46580_ (_13688_, _38797_, _38794_);
  nand _46581_ (_38798_, _38588_, _30567_);
  not _46582_ (_38799_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand _46583_ (_38800_, _38587_, _38799_);
  and _46584_ (_38801_, _38800_, _41806_);
  and _46585_ (_13698_, _38801_, _38798_);
  nand _46586_ (_38802_, _38588_, _31338_);
  or _46587_ (_38803_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _46588_ (_38804_, _38803_, _41806_);
  and _46589_ (_13708_, _38804_, _38802_);
  nand _46590_ (_38805_, _38588_, _32044_);
  or _46591_ (_38806_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _46592_ (_38807_, _38806_, _41806_);
  and _46593_ (_13718_, _38807_, _38805_);
  nand _46594_ (_38808_, _38588_, _32853_);
  or _46595_ (_38809_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _46596_ (_38810_, _38809_, _41806_);
  and _46597_ (_13727_, _38810_, _38808_);
  nand _46598_ (_38812_, _38588_, _33598_);
  or _46599_ (_38815_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _46600_ (_38816_, _38815_, _41806_);
  and _46601_ (_13736_, _38816_, _38812_);
  and _46602_ (_38817_, _28087_, _24456_);
  nor _46603_ (_38818_, _24665_, _24949_);
  and _46604_ (_38819_, _25255_, _24796_);
  and _46605_ (_38820_, _38819_, _38818_);
  and _46606_ (_38821_, _38820_, _38817_);
  nor _46607_ (_38822_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _46608_ (_38823_, _38822_);
  and _46609_ (_38824_, _38823_, _28676_);
  and _46610_ (_38833_, _38820_, _28742_);
  not _46611_ (_38839_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _46612_ (_38845_, _38822_, _38839_);
  nor _46613_ (_38849_, _38845_, _38833_);
  not _46614_ (_38850_, _38849_);
  nor _46615_ (_38851_, _38850_, _38824_);
  not _46616_ (_38852_, _38833_);
  not _46617_ (_38853_, _28709_);
  nor _46618_ (_38854_, _38853_, _28676_);
  nor _46619_ (_38855_, _28709_, _38839_);
  nor _46620_ (_38856_, _38855_, _38854_);
  nor _46621_ (_38857_, _38856_, _38852_);
  nor _46622_ (_38858_, _38857_, _38851_);
  or _46623_ (_38859_, _38858_, _38821_);
  not _46624_ (_38860_, _38821_);
  or _46625_ (_38861_, _38860_, _38162_);
  and _46626_ (_38862_, _38861_, _38859_);
  nor _46627_ (_16545_, _38862_, rst);
  nor _46628_ (_38863_, _38860_, _38417_);
  not _46629_ (_38864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand _46630_ (_38865_, _38833_, _30002_);
  nand _46631_ (_38866_, _38865_, _38864_);
  and _46632_ (_38867_, _38866_, _38860_);
  or _46633_ (_38868_, _38865_, _29318_);
  and _46634_ (_38869_, _38868_, _38867_);
  or _46635_ (_38870_, _38869_, _38863_);
  and _46636_ (_21479_, _38870_, _41806_);
  nand _46637_ (_38871_, _38821_, _38410_);
  or _46638_ (_38873_, _20811_, _20779_);
  or _46639_ (_38875_, _38873_, _20842_);
  or _46640_ (_38876_, _38875_, _20885_);
  or _46641_ (_38877_, _38876_, _20959_);
  or _46642_ (_38878_, _38877_, _20991_);
  or _46643_ (_38879_, _38878_, _20451_);
  and _46644_ (_38880_, _38879_, _15702_);
  or _46645_ (_38881_, _28218_, _26572_);
  not _46646_ (_38882_, _28207_);
  nand _46647_ (_38883_, _38882_, _26572_);
  and _46648_ (_38884_, _38883_, _25353_);
  and _46649_ (_38885_, _38884_, _38881_);
  not _46650_ (_38886_, _25375_);
  nand _46651_ (_38887_, _27007_, _38886_);
  nor _46652_ (_38888_, _28153_, _28164_);
  and _46653_ (_38889_, _38888_, _38887_);
  and _46654_ (_38890_, _38515_, _22269_);
  and _46655_ (_38891_, _38513_, _21055_);
  nand _46656_ (_38892_, _38891_, _38890_);
  nand _46657_ (_38893_, _38892_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _46658_ (_38894_, _38893_, _38889_);
  or _46659_ (_38895_, _38894_, _38885_);
  or _46660_ (_38896_, _38895_, _31587_);
  or _46661_ (_38897_, _38896_, _38880_);
  nor _46662_ (_38898_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _46663_ (_38899_, _38898_, _38833_);
  and _46664_ (_38900_, _38899_, _38897_);
  not _46665_ (_38901_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _46666_ (_38902_, _30708_, _38901_);
  or _46667_ (_38903_, _38902_, _30719_);
  and _46668_ (_38904_, _38903_, _38833_);
  or _46669_ (_38905_, _38904_, _38821_);
  or _46670_ (_38906_, _38905_, _38900_);
  and _46671_ (_38907_, _38906_, _38871_);
  and _46672_ (_21490_, _38907_, _41806_);
  nor _46673_ (_38908_, _38860_, _38402_);
  and _46674_ (_38909_, _38833_, _31436_);
  and _46675_ (_38910_, _38909_, _28676_);
  nor _46676_ (_38912_, _38909_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _46677_ (_38915_, _38912_, _38821_);
  not _46678_ (_38921_, _38915_);
  nor _46679_ (_38926_, _38921_, _38910_);
  nor _46680_ (_38933_, _38926_, _38908_);
  nor _46681_ (_21502_, _38933_, rst);
  not _46682_ (_38949_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  not _46683_ (_38950_, _24665_);
  nand _46684_ (_38951_, _38819_, _38950_);
  not _46685_ (_38952_, _28742_);
  nor _46686_ (_38953_, _38952_, _24949_);
  not _46687_ (_38954_, _38953_);
  nor _46688_ (_38955_, _38954_, _38951_);
  and _46689_ (_38956_, _38955_, _32163_);
  nor _46690_ (_38957_, _38956_, _38949_);
  and _46691_ (_38958_, _32142_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _46692_ (_38959_, _38958_, _32196_);
  nor _46693_ (_38960_, _38959_, _38852_);
  nor _46694_ (_38961_, _38960_, _38957_);
  nor _46695_ (_38962_, _38961_, _38821_);
  nor _46696_ (_38963_, _38860_, _38394_);
  nor _46697_ (_38964_, _38963_, _38962_);
  nor _46698_ (_21514_, _38964_, rst);
  nand _46699_ (_38965_, _38833_, _32941_);
  nor _46700_ (_38966_, _38965_, _28676_);
  and _46701_ (_38967_, _38965_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _46702_ (_38968_, _38967_, _38821_);
  or _46703_ (_38969_, _38968_, _38966_);
  nand _46704_ (_38970_, _38821_, _38366_);
  and _46705_ (_38971_, _38970_, _38969_);
  and _46706_ (_21526_, _38971_, _41806_);
  and _46707_ (_38972_, _33697_, _29318_);
  nor _46708_ (_38973_, _33697_, _31066_);
  nor _46709_ (_38974_, _38973_, _38972_);
  nor _46710_ (_38975_, _38974_, _38852_);
  and _46711_ (_38976_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _46712_ (_38977_, _38976_);
  nor _46713_ (_38978_, _38977_, _27813_);
  nor _46714_ (_38979_, _38978_, _31066_);
  and _46715_ (_38980_, _26659_, _26909_);
  and _46716_ (_38981_, _26528_, _25353_);
  nor _46717_ (_38982_, _38981_, _38980_);
  nor _46718_ (_38983_, _38982_, _38977_);
  nor _46719_ (_38984_, _38983_, _38979_);
  nor _46720_ (_38988_, _38984_, _38833_);
  nor _46721_ (_38999_, _38988_, _38975_);
  nor _46722_ (_39002_, _38999_, _38821_);
  nor _46723_ (_39003_, _38860_, _38280_);
  nor _46724_ (_39004_, _39003_, _39002_);
  nor _46725_ (_21538_, _39004_, rst);
  not _46726_ (_39020_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46727_ (_39021_, _38492_, _39020_);
  not _46728_ (_39022_, _39021_);
  or _46729_ (_39023_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _46730_ (_39024_, _39023_, _39020_);
  and _46731_ (_39025_, _24197_, _25112_);
  and _46732_ (_39026_, _39025_, _24445_);
  not _46733_ (_39027_, _24796_);
  and _46734_ (_39028_, _25244_, _39027_);
  and _46735_ (_39029_, _39028_, _28087_);
  and _46736_ (_39030_, _39029_, _39026_);
  nand _46737_ (_39031_, _39030_, _38818_);
  and _46738_ (_39032_, _39031_, _39024_);
  nor _46739_ (_39033_, _39032_, _28011_);
  and _46740_ (_39034_, _25244_, _25112_);
  and _46741_ (_39035_, _39034_, _24807_);
  and _46742_ (_39036_, _39035_, _38953_);
  and _46743_ (_39037_, _39036_, _28709_);
  and _46744_ (_39038_, _39037_, _28676_);
  nor _46745_ (_39039_, _39037_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _46746_ (_39040_, _39039_);
  and _46747_ (_39041_, _39032_, _39022_);
  and _46748_ (_39042_, _39041_, _39040_);
  not _46749_ (_39043_, _39042_);
  nor _46750_ (_39044_, _39043_, _39038_);
  or _46751_ (_39045_, _39044_, _39033_);
  and _46752_ (_39046_, _39045_, _39022_);
  nor _46753_ (_39047_, _39022_, _38582_);
  or _46754_ (_39048_, _39047_, _39046_);
  and _46755_ (_22313_, _39048_, _41806_);
  nor _46756_ (_39049_, _39032_, _29231_);
  and _46757_ (_39050_, _39036_, _24456_);
  and _46758_ (_39051_, _39050_, _28676_);
  nor _46759_ (_39052_, _39050_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not _46760_ (_39053_, _39052_);
  and _46761_ (_39054_, _39053_, _39041_);
  not _46762_ (_39055_, _39054_);
  nor _46763_ (_39056_, _39055_, _39051_);
  or _46764_ (_39057_, _39056_, _39049_);
  and _46765_ (_39058_, _39057_, _39022_);
  nor _46766_ (_39059_, _39022_, _38617_);
  or _46767_ (_39060_, _39059_, _39058_);
  and _46768_ (_24174_, _39060_, _41806_);
  and _46769_ (_39061_, _39021_, _38645_);
  nor _46770_ (_39062_, _39032_, _29893_);
  and _46771_ (_39063_, _39036_, _30002_);
  and _46772_ (_39064_, _39063_, _28676_);
  nor _46773_ (_39065_, _39063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not _46774_ (_39066_, _39065_);
  and _46775_ (_39067_, _39066_, _39041_);
  not _46776_ (_39068_, _39067_);
  nor _46777_ (_39069_, _39068_, _39064_);
  nor _46778_ (_39070_, _39069_, _39021_);
  not _46779_ (_39071_, _39070_);
  nor _46780_ (_39072_, _39071_, _39062_);
  nor _46781_ (_39073_, _39072_, _39061_);
  and _46782_ (_24186_, _39073_, _41806_);
  nor _46783_ (_39074_, _39032_, _30567_);
  nor _46784_ (_39075_, _25113_, _24949_);
  and _46785_ (_39076_, _39075_, _25244_);
  and _46786_ (_39077_, _28742_, _24807_);
  and _46787_ (_39078_, _39077_, _39076_);
  not _46788_ (_39079_, _39078_);
  and _46789_ (_39080_, _39041_, _39079_);
  and _46790_ (_39081_, _39080_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _46791_ (_39082_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _46792_ (_39083_, _30708_, _39082_);
  nor _46793_ (_39084_, _39083_, _30719_);
  and _46794_ (_39085_, _39041_, _39078_);
  not _46795_ (_39086_, _39085_);
  nor _46796_ (_39087_, _39086_, _39084_);
  nor _46797_ (_39088_, _39087_, _39081_);
  and _46798_ (_39089_, _39088_, _39022_);
  not _46799_ (_39090_, _39089_);
  nor _46800_ (_39091_, _39090_, _39074_);
  and _46801_ (_39092_, _39021_, _38673_);
  or _46802_ (_39093_, _39092_, _39091_);
  nor _46803_ (_24198_, _39093_, rst);
  nor _46804_ (_39094_, _39032_, _31338_);
  and _46805_ (_39095_, _39080_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _46806_ (_39096_, _31447_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _46807_ (_39097_, _39096_, _31458_);
  nor _46808_ (_39098_, _39097_, _39086_);
  nor _46809_ (_39099_, _39098_, _39095_);
  not _46810_ (_39100_, _39099_);
  nor _46811_ (_39101_, _39100_, _39094_);
  nor _46812_ (_39102_, _39101_, _39021_);
  nor _46813_ (_39103_, _39022_, _38702_);
  nor _46814_ (_39104_, _39103_, _39102_);
  nor _46815_ (_24210_, _39104_, rst);
  nor _46816_ (_39105_, _39032_, _32044_);
  and _46817_ (_39106_, _39036_, _32131_);
  and _46818_ (_39107_, _39106_, _28676_);
  nor _46819_ (_39108_, _39106_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not _46820_ (_39109_, _39108_);
  and _46821_ (_39110_, _39109_, _39041_);
  not _46822_ (_39111_, _39110_);
  nor _46823_ (_39112_, _39111_, _39107_);
  or _46824_ (_39113_, _39112_, _39105_);
  and _46825_ (_39114_, _39113_, _39022_);
  nor _46826_ (_39115_, _39022_, _38731_);
  or _46827_ (_39116_, _39115_, _39114_);
  and _46828_ (_24222_, _39116_, _41806_);
  nor _46829_ (_39117_, _39032_, _32853_);
  and _46830_ (_39118_, _39036_, _32941_);
  and _46831_ (_39119_, _39118_, _28676_);
  nor _46832_ (_39120_, _39118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not _46833_ (_39121_, _39120_);
  and _46834_ (_39122_, _39121_, _39041_);
  not _46835_ (_39123_, _39122_);
  nor _46836_ (_39124_, _39123_, _39119_);
  or _46837_ (_39125_, _39124_, _39117_);
  and _46838_ (_39126_, _39125_, _39022_);
  nor _46839_ (_39127_, _39022_, _38760_);
  or _46840_ (_39128_, _39127_, _39126_);
  and _46841_ (_24234_, _39128_, _41806_);
  nor _46842_ (_39129_, _39032_, _33598_);
  and _46843_ (_39130_, _39036_, _33697_);
  and _46844_ (_39131_, _39130_, _28676_);
  nor _46845_ (_39132_, _39130_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not _46846_ (_39133_, _39132_);
  and _46847_ (_39134_, _39133_, _39041_);
  not _46848_ (_39135_, _39134_);
  nor _46849_ (_39136_, _39135_, _39131_);
  or _46850_ (_39137_, _39136_, _39129_);
  and _46851_ (_39138_, _39137_, _39022_);
  nor _46852_ (_39139_, _39022_, _38787_);
  or _46853_ (_39140_, _39139_, _39138_);
  and _46854_ (_24246_, _39140_, _41806_);
  and _46855_ (_39141_, _38019_, _28709_);
  nand _46856_ (_39142_, _39141_, _28676_);
  or _46857_ (_39143_, _39141_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46858_ (_39144_, _39143_, _28742_);
  and _46859_ (_39145_, _39144_, _39142_);
  and _46860_ (_39146_, _38008_, _39026_);
  nand _46861_ (_39147_, _39146_, _38162_);
  or _46862_ (_39148_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46863_ (_39149_, _39148_, _28087_);
  and _46864_ (_39150_, _39149_, _39147_);
  not _46865_ (_39151_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor _46866_ (_39152_, _28076_, _39151_);
  or _46867_ (_39153_, _39152_, rst);
  or _46868_ (_39154_, _39153_, _39150_);
  or _46869_ (_35484_, _39154_, _39145_);
  nor _46870_ (_39155_, _38950_, _24949_);
  and _46871_ (_39156_, _38819_, _39155_);
  and _46872_ (_39157_, _39156_, _28709_);
  nand _46873_ (_39158_, _39157_, _28676_);
  or _46874_ (_39159_, _39157_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46875_ (_39160_, _39159_, _28742_);
  and _46876_ (_39161_, _39160_, _39158_);
  and _46877_ (_39162_, _39156_, _24456_);
  not _46878_ (_39163_, _39162_);
  nor _46879_ (_39164_, _39163_, _38162_);
  not _46880_ (_39165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor _46881_ (_39166_, _39162_, _39165_);
  or _46882_ (_39167_, _39166_, _39164_);
  and _46883_ (_39168_, _39167_, _28087_);
  nor _46884_ (_39169_, _28076_, _39165_);
  or _46885_ (_39170_, _39169_, rst);
  or _46886_ (_39171_, _39170_, _39168_);
  or _46887_ (_35507_, _39171_, _39161_);
  and _46888_ (_39172_, _39027_, _24665_);
  and _46889_ (_39173_, _39172_, _39076_);
  and _46890_ (_39174_, _39173_, _28709_);
  nand _46891_ (_39175_, _39174_, _28676_);
  or _46892_ (_39176_, _39174_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _46893_ (_39177_, _39176_, _28742_);
  and _46894_ (_39178_, _39177_, _39175_);
  and _46895_ (_39179_, _39028_, _39155_);
  and _46896_ (_39180_, _39179_, _39026_);
  not _46897_ (_39181_, _39180_);
  nor _46898_ (_39182_, _39181_, _38162_);
  not _46899_ (_39183_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor _46900_ (_39184_, _39180_, _39183_);
  or _46901_ (_39185_, _39184_, _39182_);
  and _46902_ (_39186_, _39185_, _28087_);
  nor _46903_ (_39187_, _28076_, _39183_);
  or _46904_ (_39188_, _39187_, rst);
  or _46905_ (_39189_, _39188_, _39186_);
  or _46906_ (_35530_, _39189_, _39178_);
  and _46907_ (_39190_, _39172_, _25266_);
  and _46908_ (_39191_, _39190_, _28709_);
  nand _46909_ (_39192_, _39191_, _28676_);
  or _46910_ (_39193_, _39191_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _46911_ (_39194_, _39193_, _28742_);
  and _46912_ (_39195_, _39194_, _39192_);
  nor _46913_ (_39196_, _25244_, _24796_);
  and _46914_ (_39203_, _39155_, _39196_);
  and _46915_ (_39214_, _39203_, _39026_);
  not _46916_ (_39225_, _39214_);
  nor _46917_ (_39235_, _39225_, _38162_);
  not _46918_ (_39241_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor _46919_ (_39251_, _39214_, _39241_);
  or _46920_ (_39262_, _39251_, _39235_);
  and _46921_ (_39273_, _39262_, _28087_);
  nor _46922_ (_39284_, _28076_, _39241_);
  or _46923_ (_39295_, _39284_, rst);
  or _46924_ (_39306_, _39295_, _39273_);
  or _46925_ (_35552_, _39306_, _39195_);
  not _46926_ (_39327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _46927_ (_39338_, _39146_, _39327_);
  nand _46928_ (_39349_, _38019_, _24456_);
  nor _46929_ (_39360_, _39349_, _28676_);
  or _46930_ (_39371_, _39360_, _39338_);
  and _46931_ (_39382_, _39371_, _28742_);
  and _46932_ (_39393_, _39146_, _38426_);
  or _46933_ (_39404_, _39393_, _39338_);
  and _46934_ (_39410_, _39404_, _28087_);
  nor _46935_ (_39411_, _28076_, _39327_);
  or _46936_ (_39412_, _39411_, rst);
  or _46937_ (_39413_, _39412_, _39410_);
  or _46938_ (_41207_, _39413_, _39382_);
  or _46939_ (_39414_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46940_ (_39415_, _39414_, _28742_);
  nand _46941_ (_39416_, _38205_, _28676_);
  and _46942_ (_39417_, _39416_, _39415_);
  nand _46943_ (_39418_, _39146_, _38417_);
  or _46944_ (_39419_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46945_ (_39420_, _39419_, _28087_);
  and _46946_ (_39421_, _39420_, _39418_);
  not _46947_ (_39422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor _46948_ (_39423_, _28076_, _39422_);
  or _46949_ (_39424_, _39423_, rst);
  or _46950_ (_39425_, _39424_, _39421_);
  or _46951_ (_41209_, _39425_, _39417_);
  not _46952_ (_39426_, _31468_);
  nand _46953_ (_39427_, _38019_, _39426_);
  and _46954_ (_39428_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46955_ (_39429_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _46956_ (_39430_, _39429_, _30719_);
  and _46957_ (_39431_, _39430_, _38019_);
  or _46958_ (_39432_, _39431_, _39428_);
  and _46959_ (_39433_, _39432_, _28742_);
  nand _46960_ (_39434_, _39146_, _38410_);
  or _46961_ (_39435_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46962_ (_39436_, _39435_, _28087_);
  and _46963_ (_39437_, _39436_, _39434_);
  not _46964_ (_39438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor _46965_ (_39439_, _28076_, _39438_);
  or _46966_ (_39440_, _39439_, rst);
  or _46967_ (_39441_, _39440_, _39437_);
  or _46968_ (_41211_, _39441_, _39433_);
  not _46969_ (_39442_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor _46970_ (_39443_, _38194_, _39442_);
  nor _46971_ (_39444_, _31468_, _39442_);
  or _46972_ (_39445_, _39444_, _31458_);
  and _46973_ (_39446_, _39445_, _38019_);
  or _46974_ (_39447_, _39446_, _39443_);
  and _46975_ (_39448_, _39447_, _28742_);
  nand _46976_ (_39449_, _39146_, _38402_);
  or _46977_ (_39450_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46978_ (_39451_, _39450_, _28087_);
  and _46979_ (_39452_, _39451_, _39449_);
  nor _46980_ (_39453_, _28076_, _39442_);
  or _46981_ (_39454_, _39453_, rst);
  or _46982_ (_39455_, _39454_, _39452_);
  or _46983_ (_41213_, _39455_, _39448_);
  nand _46984_ (_39456_, _38019_, _32163_);
  and _46985_ (_39457_, _39456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46986_ (_39458_, _32142_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46987_ (_39459_, _39458_, _32196_);
  and _46988_ (_39460_, _39459_, _38019_);
  or _46989_ (_39461_, _39460_, _39457_);
  and _46990_ (_39462_, _39461_, _28742_);
  nand _46991_ (_39463_, _39146_, _38394_);
  or _46992_ (_39464_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46993_ (_39465_, _39464_, _28087_);
  and _46994_ (_39466_, _39465_, _39463_);
  not _46995_ (_39467_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor _46996_ (_39468_, _28076_, _39467_);
  or _46997_ (_39469_, _39468_, rst);
  or _46998_ (_39470_, _39469_, _39466_);
  or _46999_ (_41214_, _39470_, _39462_);
  and _47000_ (_39471_, _38019_, _32941_);
  nand _47001_ (_39472_, _39471_, _28676_);
  or _47002_ (_39473_, _39471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _47003_ (_39474_, _39473_, _28742_);
  and _47004_ (_39475_, _39474_, _39472_);
  nand _47005_ (_39476_, _39146_, _38366_);
  or _47006_ (_39477_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _47007_ (_39478_, _39477_, _28087_);
  and _47008_ (_39479_, _39478_, _39476_);
  not _47009_ (_39480_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor _47010_ (_39481_, _28076_, _39480_);
  or _47011_ (_39482_, _39481_, rst);
  or _47012_ (_39483_, _39482_, _39479_);
  or _47013_ (_41216_, _39483_, _39475_);
  and _47014_ (_39484_, _38019_, _33697_);
  nand _47015_ (_39485_, _39484_, _28676_);
  or _47016_ (_39486_, _39484_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _47017_ (_39487_, _39486_, _28742_);
  and _47018_ (_39488_, _39487_, _39485_);
  nand _47019_ (_39489_, _39146_, _38280_);
  or _47020_ (_39490_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _47021_ (_39491_, _39490_, _28087_);
  and _47022_ (_39492_, _39491_, _39489_);
  not _47023_ (_39493_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _47024_ (_39494_, _28076_, _39493_);
  or _47025_ (_39495_, _39494_, rst);
  or _47026_ (_39496_, _39495_, _39492_);
  or _47027_ (_41218_, _39496_, _39488_);
  nand _47028_ (_39497_, _39162_, _28676_);
  or _47029_ (_39498_, _39162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _47030_ (_39499_, _39498_, _28742_);
  and _47031_ (_39500_, _39499_, _39497_);
  nor _47032_ (_39501_, _39163_, _38425_);
  not _47033_ (_39502_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _47034_ (_39503_, _39162_, _39502_);
  or _47035_ (_39504_, _39503_, _39501_);
  and _47036_ (_39505_, _39504_, _28087_);
  nor _47037_ (_39506_, _28076_, _39502_);
  or _47038_ (_39507_, _39506_, rst);
  or _47039_ (_39508_, _39507_, _39505_);
  or _47040_ (_41220_, _39508_, _39500_);
  and _47041_ (_39509_, _39156_, _30002_);
  nand _47042_ (_39510_, _39509_, _28676_);
  or _47043_ (_39511_, _39509_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _47044_ (_39512_, _39511_, _28742_);
  and _47045_ (_39513_, _39512_, _39510_);
  nor _47046_ (_39514_, _39163_, _38417_);
  not _47047_ (_39515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor _47048_ (_39516_, _39162_, _39515_);
  or _47049_ (_39517_, _39516_, _39514_);
  and _47050_ (_39518_, _39517_, _28087_);
  nor _47051_ (_39519_, _28076_, _39515_);
  or _47052_ (_39520_, _39519_, rst);
  or _47053_ (_39521_, _39520_, _39518_);
  or _47054_ (_41221_, _39521_, _39513_);
  and _47055_ (_39522_, _39156_, _30708_);
  nand _47056_ (_39523_, _39522_, _28676_);
  or _47057_ (_39524_, _39522_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _47058_ (_39525_, _39524_, _28742_);
  and _47059_ (_39526_, _39525_, _39523_);
  nor _47060_ (_39527_, _39163_, _38410_);
  not _47061_ (_39528_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor _47062_ (_39529_, _39162_, _39528_);
  or _47063_ (_39530_, _39529_, _39527_);
  and _47064_ (_39531_, _39530_, _28087_);
  nor _47065_ (_39532_, _28076_, _39528_);
  or _47066_ (_39533_, _39532_, rst);
  or _47067_ (_39534_, _39533_, _39531_);
  or _47068_ (_41223_, _39534_, _39526_);
  and _47069_ (_39535_, _39156_, _31436_);
  nand _47070_ (_39536_, _39535_, _28676_);
  or _47071_ (_39537_, _39535_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _47072_ (_39538_, _39537_, _28742_);
  and _47073_ (_39539_, _39538_, _39536_);
  nor _47074_ (_39540_, _39163_, _38402_);
  not _47075_ (_39541_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor _47076_ (_39542_, _39162_, _39541_);
  or _47077_ (_39543_, _39542_, _39540_);
  and _47078_ (_39544_, _39543_, _28087_);
  nor _47079_ (_39545_, _28076_, _39541_);
  or _47080_ (_39546_, _39545_, rst);
  or _47081_ (_39547_, _39546_, _39544_);
  or _47082_ (_41225_, _39547_, _39539_);
  and _47083_ (_39548_, _39156_, _32131_);
  nand _47084_ (_39549_, _39548_, _28676_);
  or _47085_ (_39550_, _39548_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47086_ (_39551_, _39550_, _28742_);
  and _47087_ (_39552_, _39551_, _39549_);
  nor _47088_ (_39553_, _39163_, _38394_);
  not _47089_ (_39554_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor _47090_ (_39555_, _39162_, _39554_);
  or _47091_ (_39556_, _39555_, _39553_);
  and _47092_ (_39557_, _39556_, _28087_);
  nor _47093_ (_39558_, _28076_, _39554_);
  or _47094_ (_39559_, _39558_, rst);
  or _47095_ (_39560_, _39559_, _39557_);
  or _47096_ (_41227_, _39560_, _39552_);
  and _47097_ (_39561_, _39156_, _32941_);
  nand _47098_ (_39562_, _39561_, _28676_);
  or _47099_ (_39563_, _39561_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _47100_ (_39564_, _39563_, _28742_);
  and _47101_ (_39565_, _39564_, _39562_);
  nor _47102_ (_39566_, _39163_, _38366_);
  not _47103_ (_39567_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor _47104_ (_39568_, _39162_, _39567_);
  or _47105_ (_39569_, _39568_, _39566_);
  and _47106_ (_39570_, _39569_, _28087_);
  nor _47107_ (_39571_, _28076_, _39567_);
  or _47108_ (_39572_, _39571_, rst);
  or _47109_ (_39573_, _39572_, _39570_);
  or _47110_ (_41228_, _39573_, _39565_);
  and _47111_ (_39574_, _39156_, _33697_);
  nand _47112_ (_39575_, _39574_, _28676_);
  or _47113_ (_39576_, _39574_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _47114_ (_39577_, _39576_, _28742_);
  and _47115_ (_39578_, _39577_, _39575_);
  nor _47116_ (_39579_, _39163_, _38280_);
  not _47117_ (_39580_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _47118_ (_39581_, _39162_, _39580_);
  or _47119_ (_39582_, _39581_, _39579_);
  and _47120_ (_39583_, _39582_, _28087_);
  nor _47121_ (_39584_, _28076_, _39580_);
  or _47122_ (_39585_, _39584_, rst);
  or _47123_ (_39586_, _39585_, _39583_);
  or _47124_ (_41230_, _39586_, _39578_);
  nand _47125_ (_39587_, _39180_, _28676_);
  or _47126_ (_39588_, _39180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _47127_ (_39589_, _39588_, _28742_);
  and _47128_ (_39590_, _39589_, _39587_);
  nor _47129_ (_39591_, _39181_, _38425_);
  not _47130_ (_39592_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _47131_ (_39593_, _39180_, _39592_);
  or _47132_ (_39594_, _39593_, _39591_);
  and _47133_ (_39595_, _39594_, _28087_);
  nor _47134_ (_39596_, _28076_, _39592_);
  or _47135_ (_39597_, _39596_, rst);
  or _47136_ (_39598_, _39597_, _39595_);
  or _47137_ (_41232_, _39598_, _39590_);
  and _47138_ (_39599_, _39173_, _30002_);
  nand _47139_ (_39600_, _39599_, _28676_);
  or _47140_ (_39601_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _47141_ (_39602_, _39601_, _28742_);
  and _47142_ (_39603_, _39602_, _39600_);
  nor _47143_ (_39604_, _39181_, _38417_);
  not _47144_ (_39605_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor _47145_ (_39606_, _39180_, _39605_);
  or _47146_ (_39607_, _39606_, _39604_);
  and _47147_ (_39608_, _39607_, _28087_);
  nor _47148_ (_39609_, _28076_, _39605_);
  or _47149_ (_39610_, _39609_, rst);
  or _47150_ (_39611_, _39610_, _39608_);
  or _47151_ (_41234_, _39611_, _39603_);
  and _47152_ (_39612_, _39173_, _30708_);
  nand _47153_ (_39613_, _39612_, _28676_);
  or _47154_ (_39614_, _39612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _47155_ (_39615_, _39614_, _28742_);
  and _47156_ (_39616_, _39615_, _39613_);
  nor _47157_ (_39618_, _39181_, _38410_);
  not _47158_ (_39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor _47159_ (_39620_, _39180_, _39619_);
  or _47160_ (_39621_, _39620_, _39618_);
  and _47161_ (_39622_, _39621_, _28087_);
  nor _47162_ (_39623_, _28076_, _39619_);
  or _47163_ (_39624_, _39623_, rst);
  or _47164_ (_39625_, _39624_, _39622_);
  or _47165_ (_41235_, _39625_, _39616_);
  and _47166_ (_39626_, _39173_, _31436_);
  nand _47167_ (_39627_, _39626_, _28676_);
  or _47168_ (_39628_, _39626_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _47169_ (_39629_, _39628_, _28742_);
  and _47170_ (_39630_, _39629_, _39627_);
  nor _47171_ (_39631_, _39181_, _38402_);
  not _47172_ (_39632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor _47173_ (_39633_, _39180_, _39632_);
  or _47174_ (_39634_, _39633_, _39631_);
  and _47175_ (_39635_, _39634_, _28087_);
  nor _47176_ (_39636_, _28076_, _39632_);
  or _47177_ (_39637_, _39636_, rst);
  or _47178_ (_39638_, _39637_, _39635_);
  or _47179_ (_41237_, _39638_, _39630_);
  and _47180_ (_39639_, _39173_, _32131_);
  nand _47181_ (_39640_, _39639_, _28676_);
  or _47182_ (_39641_, _39639_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _47183_ (_39642_, _39641_, _28742_);
  and _47184_ (_39643_, _39642_, _39640_);
  nor _47185_ (_39644_, _39181_, _38394_);
  not _47186_ (_39645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _47187_ (_39646_, _39180_, _39645_);
  or _47188_ (_39647_, _39646_, _39644_);
  and _47189_ (_39652_, _39647_, _28087_);
  nor _47190_ (_39653_, _28076_, _39645_);
  or _47191_ (_39654_, _39653_, rst);
  or _47192_ (_39655_, _39654_, _39652_);
  or _47193_ (_41239_, _39655_, _39643_);
  and _47194_ (_39656_, _39173_, _32941_);
  nand _47195_ (_39657_, _39656_, _28676_);
  or _47196_ (_39658_, _39656_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _47197_ (_39659_, _39658_, _28742_);
  and _47198_ (_39660_, _39659_, _39657_);
  nor _47199_ (_39661_, _39181_, _38366_);
  not _47200_ (_39662_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor _47201_ (_39663_, _39180_, _39662_);
  or _47202_ (_39664_, _39663_, _39661_);
  and _47203_ (_39665_, _39664_, _28087_);
  nor _47204_ (_39666_, _28076_, _39662_);
  or _47205_ (_39667_, _39666_, rst);
  or _47206_ (_39668_, _39667_, _39665_);
  or _47207_ (_41240_, _39668_, _39660_);
  and _47208_ (_39669_, _39173_, _33697_);
  nand _47209_ (_39670_, _39669_, _28676_);
  or _47210_ (_39671_, _39669_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47211_ (_39672_, _39671_, _28742_);
  and _47212_ (_39673_, _39672_, _39670_);
  nor _47213_ (_39674_, _39181_, _38280_);
  not _47214_ (_39675_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor _47215_ (_39676_, _39180_, _39675_);
  or _47216_ (_39677_, _39676_, _39674_);
  and _47217_ (_39678_, _39677_, _28087_);
  nor _47218_ (_39679_, _28076_, _39675_);
  or _47219_ (_39680_, _39679_, rst);
  or _47220_ (_39681_, _39680_, _39678_);
  or _47221_ (_41242_, _39681_, _39673_);
  and _47222_ (_39682_, _39190_, _24456_);
  nand _47223_ (_39683_, _39682_, _28676_);
  or _47224_ (_39684_, _39682_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _47225_ (_39685_, _39684_, _28742_);
  and _47226_ (_39686_, _39685_, _39683_);
  nor _47227_ (_39687_, _39225_, _38425_);
  not _47228_ (_39688_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _47229_ (_39689_, _39214_, _39688_);
  or _47230_ (_39690_, _39689_, _39687_);
  and _47231_ (_39691_, _39690_, _28087_);
  nor _47232_ (_39692_, _28076_, _39688_);
  or _47233_ (_39693_, _39692_, rst);
  or _47234_ (_39694_, _39693_, _39691_);
  or _47235_ (_41244_, _39694_, _39686_);
  and _47236_ (_39695_, _39190_, _30002_);
  nand _47237_ (_39696_, _39695_, _28676_);
  or _47238_ (_39697_, _39695_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _47239_ (_39698_, _39697_, _28742_);
  and _47240_ (_39699_, _39698_, _39696_);
  nor _47241_ (_39700_, _39225_, _38417_);
  not _47242_ (_39701_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor _47243_ (_39702_, _39214_, _39701_);
  or _47244_ (_39703_, _39702_, _39700_);
  and _47245_ (_39704_, _39703_, _28087_);
  nor _47246_ (_39705_, _28076_, _39701_);
  or _47247_ (_39706_, _39705_, rst);
  or _47248_ (_39707_, _39706_, _39704_);
  or _47249_ (_41245_, _39707_, _39699_);
  and _47250_ (_39708_, _39190_, _30708_);
  nand _47251_ (_39709_, _39708_, _28676_);
  or _47252_ (_39710_, _39708_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _47253_ (_39711_, _39710_, _28742_);
  and _47254_ (_39712_, _39711_, _39709_);
  nor _47255_ (_39720_, _39225_, _38410_);
  not _47256_ (_39721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor _47257_ (_39722_, _39214_, _39721_);
  or _47258_ (_39723_, _39722_, _39720_);
  and _47259_ (_39724_, _39723_, _28087_);
  nor _47260_ (_39725_, _28076_, _39721_);
  or _47261_ (_39726_, _39725_, rst);
  or _47262_ (_39727_, _39726_, _39724_);
  or _47263_ (_41247_, _39727_, _39712_);
  and _47264_ (_39728_, _39190_, _31436_);
  nand _47265_ (_39729_, _39728_, _28676_);
  or _47266_ (_39730_, _39728_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _47267_ (_39731_, _39730_, _28742_);
  and _47268_ (_39732_, _39731_, _39729_);
  nor _47269_ (_39733_, _39225_, _38402_);
  not _47270_ (_39734_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor _47271_ (_39735_, _39214_, _39734_);
  or _47272_ (_39736_, _39735_, _39733_);
  and _47273_ (_39737_, _39736_, _28087_);
  nor _47274_ (_39738_, _28076_, _39734_);
  or _47275_ (_39739_, _39738_, rst);
  or _47276_ (_39740_, _39739_, _39737_);
  or _47277_ (_41249_, _39740_, _39732_);
  and _47278_ (_39741_, _39190_, _32131_);
  nand _47279_ (_39742_, _39741_, _28676_);
  or _47280_ (_39743_, _39741_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47281_ (_39744_, _39743_, _28742_);
  and _47282_ (_39745_, _39744_, _39742_);
  nor _47283_ (_39746_, _39225_, _38394_);
  not _47284_ (_39747_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor _47285_ (_39748_, _39214_, _39747_);
  or _47286_ (_39749_, _39748_, _39746_);
  and _47287_ (_39750_, _39749_, _28087_);
  nor _47288_ (_39751_, _28076_, _39747_);
  or _47289_ (_39752_, _39751_, rst);
  or _47290_ (_39753_, _39752_, _39750_);
  or _47291_ (_41251_, _39753_, _39745_);
  and _47292_ (_39754_, _39190_, _32941_);
  nand _47293_ (_39755_, _39754_, _28676_);
  or _47294_ (_39756_, _39754_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _47295_ (_39757_, _39756_, _28742_);
  and _47296_ (_39758_, _39757_, _39755_);
  nor _47297_ (_39759_, _39225_, _38366_);
  not _47298_ (_39760_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor _47299_ (_39761_, _39214_, _39760_);
  or _47300_ (_39762_, _39761_, _39759_);
  and _47301_ (_39763_, _39762_, _28087_);
  nor _47302_ (_39768_, _28076_, _39760_);
  or _47303_ (_39769_, _39768_, rst);
  or _47304_ (_39770_, _39769_, _39763_);
  or _47305_ (_41252_, _39770_, _39758_);
  and _47306_ (_39771_, _39190_, _33697_);
  nand _47307_ (_39772_, _39771_, _28676_);
  or _47308_ (_39773_, _39771_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _47309_ (_39774_, _39773_, _28742_);
  and _47310_ (_39775_, _39774_, _39772_);
  nor _47311_ (_39776_, _39225_, _38280_);
  not _47312_ (_39777_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _47313_ (_39778_, _39214_, _39777_);
  or _47314_ (_39779_, _39778_, _39776_);
  and _47315_ (_39780_, _39779_, _28087_);
  nor _47316_ (_39781_, _28076_, _39777_);
  or _47317_ (_39782_, _39781_, rst);
  or _47318_ (_39792_, _39782_, _39780_);
  or _47319_ (_41254_, _39792_, _39775_);
  and _47320_ (_39793_, _38817_, _25113_);
  and _47321_ (_39794_, _39793_, _39203_);
  nor _47322_ (_39795_, _25244_, _25112_);
  and _47323_ (_39796_, _39795_, _39172_);
  and _47324_ (_39797_, _39796_, _38953_);
  and _47325_ (_39798_, _39797_, _28709_);
  nand _47326_ (_39799_, _39798_, _28676_);
  or _47327_ (_39800_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _47328_ (_39801_, _39800_, _39799_);
  or _47329_ (_39802_, _39801_, _39794_);
  nand _47330_ (_39803_, _39794_, _38162_);
  and _47331_ (_39804_, _39803_, _41806_);
  and _47332_ (_41748_, _39804_, _39802_);
  and _47333_ (_39805_, _39793_, _39179_);
  and _47334_ (_39806_, _25244_, _25113_);
  and _47335_ (_39807_, _39806_, _38953_);
  and _47336_ (_39808_, _39807_, _39172_);
  and _47337_ (_39809_, _39808_, _28709_);
  nand _47338_ (_39810_, _39809_, _28676_);
  or _47339_ (_39811_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47340_ (_39812_, _39811_, _39810_);
  or _47341_ (_39813_, _39812_, _39805_);
  nand _47342_ (_39814_, _39805_, _38162_);
  and _47343_ (_39815_, _39814_, _41806_);
  and _47344_ (_41751_, _39815_, _39813_);
  or _47345_ (_39816_, _24445_, _30697_);
  and _47346_ (_39817_, _39816_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47347_ (_39818_, _39817_, _38972_);
  and _47348_ (_39819_, _39807_, _37986_);
  and _47349_ (_39820_, _39819_, _39818_);
  and _47350_ (_39821_, _39793_, _38008_);
  nand _47351_ (_39822_, _39819_, _24434_);
  and _47352_ (_39823_, _39822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47353_ (_39824_, _39823_, _39821_);
  or _47354_ (_39825_, _39824_, _39820_);
  nand _47355_ (_39826_, _39821_, _38280_);
  and _47356_ (_39827_, _39826_, _41806_);
  and _47357_ (_41753_, _39827_, _39825_);
  not _47358_ (_39828_, _39821_);
  not _47359_ (_39829_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _47360_ (_39830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _47361_ (_39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47362_ (_39832_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39831_);
  and _47363_ (_39833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47364_ (_39834_, _39833_, _39832_);
  nor _47365_ (_39835_, _39834_, _39830_);
  or _47366_ (_39836_, _39835_, _39829_);
  and _47367_ (_39837_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _47368_ (_39838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _47369_ (_39839_, _39838_, _39837_);
  nor _47370_ (_39840_, _39839_, _39830_);
  and _47371_ (_39841_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39831_);
  and _47372_ (_39842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47373_ (_39843_, _39842_, _39841_);
  nand _47374_ (_39844_, _39843_, _39840_);
  or _47375_ (_39845_, _39844_, _39836_);
  and _47376_ (_39846_, _39845_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor _47377_ (_39847_, _24197_, _25112_);
  and _47378_ (_39848_, _28742_, _28698_);
  and _47379_ (_39849_, _39848_, _38008_);
  and _47380_ (_39850_, _39849_, _39847_);
  or _47381_ (_39851_, _39850_, _39846_);
  and _47382_ (_39852_, _39851_, _39828_);
  nand _47383_ (_39853_, _39850_, _28676_);
  and _47384_ (_39854_, _39853_, _39852_);
  nor _47385_ (_39855_, _39828_, _38162_);
  or _47386_ (_39856_, _39855_, _39854_);
  and _47387_ (_41755_, _39856_, _41806_);
  nor _47388_ (_39857_, _39843_, _39830_);
  nand _47389_ (_39858_, _39857_, _39839_);
  or _47390_ (_39859_, _39858_, _39836_);
  and _47391_ (_39860_, _39859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _47392_ (_39861_, _28742_, _29991_);
  and _47393_ (_39862_, _39861_, _38008_);
  and _47394_ (_39863_, _39862_, _39847_);
  or _47395_ (_39864_, _39863_, _39860_);
  and _47396_ (_39865_, _39864_, _39828_);
  nand _47397_ (_39866_, _39863_, _28676_);
  and _47398_ (_39867_, _39866_, _39865_);
  nor _47399_ (_39868_, _39828_, _38366_);
  or _47400_ (_39869_, _39868_, _39867_);
  and _47401_ (_41757_, _39869_, _41806_);
  not _47402_ (_39870_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _47403_ (_39871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _39870_);
  nand _47404_ (_39872_, _39835_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _47405_ (_39873_, _39857_, _39840_);
  or _47406_ (_39874_, _39873_, _39872_);
  and _47407_ (_39875_, _39874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _47408_ (_39876_, _39875_, _39871_);
  nor _47409_ (_39877_, _28687_, _25112_);
  and _47410_ (_39878_, _39862_, _39877_);
  or _47411_ (_39879_, _39878_, _39876_);
  and _47412_ (_39880_, _39879_, _39828_);
  nand _47413_ (_39881_, _39878_, _28676_);
  and _47414_ (_39882_, _39881_, _39880_);
  nor _47415_ (_39883_, _39828_, _38417_);
  or _47416_ (_39884_, _39883_, _39882_);
  and _47417_ (_41759_, _39884_, _41806_);
  and _47418_ (_39885_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _47419_ (_39886_, _39872_, _39858_);
  and _47420_ (_39887_, _39886_, _39885_);
  and _47421_ (_39888_, _39849_, _39877_);
  or _47422_ (_39889_, _39888_, _39887_);
  and _47423_ (_39890_, _39889_, _39828_);
  nand _47424_ (_39891_, _39888_, _28676_);
  and _47425_ (_39892_, _39891_, _39890_);
  nor _47426_ (_39893_, _39828_, _38402_);
  or _47427_ (_39894_, _39893_, _39892_);
  and _47428_ (_41761_, _39894_, _41806_);
  and _47429_ (_39895_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _47430_ (_39896_, _39895_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _47431_ (_39897_, _39896_);
  and _47432_ (_39898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47433_ (_39899_, _39898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47434_ (_39900_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _47435_ (_39901_, _39900_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _47436_ (_39902_, _39901_, _39899_);
  and _47437_ (_39903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _47438_ (_39904_, _39903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not _47439_ (_39905_, _39904_);
  and _47440_ (_39906_, _39905_, _39902_);
  and _47441_ (_39907_, _39906_, _39897_);
  not _47442_ (_39908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47443_ (_39909_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47444_ (_39910_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39831_);
  or _47445_ (_39911_, _39910_, _39909_);
  nor _47446_ (_39912_, _39911_, _39908_);
  nor _47447_ (_39913_, _39912_, _39830_);
  nor _47448_ (_39914_, _39913_, _39907_);
  and _47449_ (_39915_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _47450_ (_39916_, _39915_, _39831_);
  and _47451_ (_39917_, _39916_, _39914_);
  and _47452_ (_39918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39830_);
  not _47453_ (_39919_, _39918_);
  not _47454_ (_39920_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47455_ (_39921_, _39898_, _39920_);
  not _47456_ (_39922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47457_ (_39923_, _39900_, _39922_);
  nor _47458_ (_39924_, _39923_, _39921_);
  not _47459_ (_39925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _47460_ (_39926_, _39903_, _39925_);
  not _47461_ (_39927_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _47462_ (_39928_, _39895_, _39927_);
  nor _47463_ (_39929_, _39928_, _39926_);
  and _47464_ (_39930_, _39929_, _39924_);
  nor _47465_ (_39931_, _39930_, _39919_);
  nand _47466_ (_39932_, _39931_, _39916_);
  and _47467_ (_39933_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41806_);
  nand _47468_ (_39934_, _39933_, _39932_);
  nor _47469_ (_41793_, _39934_, _39917_);
  nor _47470_ (_39935_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _47471_ (_39936_, _39935_);
  nor _47472_ (_39937_, _39931_, _39914_);
  nor _47473_ (_39938_, _39937_, _39936_);
  nand _47474_ (_39939_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41806_);
  nor _47475_ (_41795_, _39939_, _39938_);
  and _47476_ (_39940_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _47477_ (_39941_, _39902_);
  or _47478_ (_39942_, _39941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _47479_ (_39943_, _39942_, _39940_);
  or _47480_ (_39944_, _39906_, _39837_);
  and _47481_ (_39945_, _39944_, _39943_);
  and _47482_ (_39946_, _39945_, _39914_);
  or _47483_ (_39947_, _39946_, _39915_);
  and _47484_ (_39948_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _47485_ (_39949_, _39914_);
  and _47486_ (_39950_, _39931_, _39949_);
  and _47487_ (_39951_, _39928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47488_ (_39952_, _39951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _47489_ (_39953_, _39924_);
  and _47490_ (_39954_, _39926_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47491_ (_39955_, _39954_, _39953_);
  and _47492_ (_39956_, _39955_, _39952_);
  and _47493_ (_39957_, _39953_, _39837_);
  or _47494_ (_39958_, _39957_, _39956_);
  and _47495_ (_39959_, _39958_, _39950_);
  or _47496_ (_39960_, _39959_, _39948_);
  or _47497_ (_39961_, _39960_, _39947_);
  not _47498_ (_39962_, _39915_);
  or _47499_ (_39963_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _47500_ (_39964_, _39963_, _41806_);
  and _47501_ (_41796_, _39964_, _39961_);
  and _47502_ (_39965_, _39896_, _39831_);
  or _47503_ (_39966_, _39941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _47504_ (_39967_, _39966_, _39965_);
  or _47505_ (_39968_, _39906_, _39838_);
  and _47506_ (_39969_, _39968_, _39967_);
  and _47507_ (_39970_, _39969_, _39914_);
  or _47508_ (_39971_, _39970_, _39915_);
  and _47509_ (_39972_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47510_ (_39973_, _39928_, _39831_);
  or _47511_ (_39974_, _39973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47512_ (_39975_, _39926_, _39831_);
  nor _47513_ (_39976_, _39975_, _39953_);
  and _47514_ (_39977_, _39976_, _39974_);
  and _47515_ (_39978_, _39953_, _39838_);
  or _47516_ (_39979_, _39978_, _39977_);
  and _47517_ (_39980_, _39979_, _39950_);
  or _47518_ (_39981_, _39980_, _39972_);
  or _47519_ (_39982_, _39981_, _39971_);
  or _47520_ (_39983_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47521_ (_39984_, _39983_, _41806_);
  and _47522_ (_41798_, _39984_, _39982_);
  nand _47523_ (_39985_, _39937_, _39830_);
  nor _47524_ (_39986_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _47525_ (_39987_, _39986_, _39915_);
  and _47526_ (_39988_, _39987_, _41806_);
  and _47527_ (_41800_, _39988_, _39985_);
  and _47528_ (_39989_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _47529_ (_39990_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _47530_ (_39991_, _39990_, _39986_);
  nor _47531_ (_39992_, _39991_, _39949_);
  or _47532_ (_39993_, _39992_, _39915_);
  or _47533_ (_39994_, _39993_, _39989_);
  or _47534_ (_39995_, _39991_, _39962_);
  and _47535_ (_39996_, _39995_, _41806_);
  and _47536_ (_41802_, _39996_, _39994_);
  and _47537_ (_39997_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41806_);
  and _47538_ (_41804_, _39997_, _39915_);
  nor _47539_ (_39998_, _39937_, _39915_);
  and _47540_ (_39999_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _47541_ (_40000_, _39999_, _39998_);
  and _47542_ (_42729_, _40000_, _41806_);
  and _47543_ (_40001_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _47544_ (_40002_, _40001_, _39998_);
  and _47545_ (_42731_, _40002_, _41806_);
  and _47546_ (_40003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _41806_);
  and _47547_ (_42733_, _40003_, _39915_);
  not _47548_ (_40004_, _39921_);
  nor _47549_ (_40005_, _39928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _47550_ (_40006_, _40005_, _39926_);
  or _47551_ (_40007_, _40006_, _39923_);
  and _47552_ (_40008_, _40007_, _40004_);
  and _47553_ (_40009_, _40008_, _39950_);
  not _47554_ (_40010_, _39899_);
  or _47555_ (_40011_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _47556_ (_40012_, _40011_, _39905_);
  or _47557_ (_40013_, _40012_, _39901_);
  and _47558_ (_40014_, _40013_, _40010_);
  and _47559_ (_40015_, _40014_, _39914_);
  or _47560_ (_40016_, _40015_, _39915_);
  or _47561_ (_40017_, _40016_, _40009_);
  or _47562_ (_40018_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _47563_ (_40019_, _40018_, _41806_);
  and _47564_ (_42734_, _40019_, _40017_);
  nand _47565_ (_40020_, _39924_, _39918_);
  nor _47566_ (_40021_, _40020_, _39929_);
  or _47567_ (_40022_, _40021_, _39914_);
  nand _47568_ (_40023_, _39914_, _39941_);
  and _47569_ (_40024_, _40023_, _40022_);
  or _47570_ (_40025_, _40024_, _39915_);
  or _47571_ (_40026_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _47572_ (_40027_, _40026_, _41806_);
  and _47573_ (_42736_, _40027_, _40025_);
  and _47574_ (_40028_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _41806_);
  and _47575_ (_42738_, _40028_, _39915_);
  and _47576_ (_40029_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _41806_);
  and _47577_ (_42740_, _40029_, _39915_);
  nand _47578_ (_40030_, _39937_, _39935_);
  nor _47579_ (_40031_, _39915_, _39914_);
  or _47580_ (_40032_, _40031_, _39831_);
  and _47581_ (_40033_, _40032_, _41806_);
  and _47582_ (_42742_, _40033_, _40030_);
  not _47583_ (_40034_, _39998_);
  and _47584_ (_40035_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _47585_ (_40036_, _39965_);
  and _47586_ (_40037_, _40036_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _47587_ (_40038_, _39904_, _39831_);
  or _47588_ (_40039_, _40038_, _39901_);
  or _47589_ (_40040_, _40039_, _40037_);
  not _47590_ (_40041_, _39901_);
  or _47591_ (_40042_, _40041_, _39833_);
  and _47592_ (_40043_, _40042_, _40040_);
  or _47593_ (_40044_, _40043_, _39899_);
  or _47594_ (_40045_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39831_);
  or _47595_ (_40046_, _40045_, _40010_);
  and _47596_ (_40047_, _40046_, _39914_);
  and _47597_ (_40048_, _40047_, _40044_);
  not _47598_ (_40049_, _39973_);
  and _47599_ (_40050_, _40049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _47600_ (_40051_, _39975_, _39923_);
  or _47601_ (_40052_, _40051_, _40050_);
  not _47602_ (_40053_, _39923_);
  or _47603_ (_40054_, _40053_, _39833_);
  and _47604_ (_40055_, _40054_, _40004_);
  and _47605_ (_40056_, _40055_, _40052_);
  and _47606_ (_40057_, _40045_, _39921_);
  or _47607_ (_40058_, _40057_, _40056_);
  and _47608_ (_40059_, _40058_, _39950_);
  or _47609_ (_40060_, _40059_, _40048_);
  and _47610_ (_40061_, _40060_, _39962_);
  or _47611_ (_40062_, _40061_, _40035_);
  and _47612_ (_42744_, _40062_, _41806_);
  and _47613_ (_40063_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _47614_ (_40064_, _40036_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _47615_ (_40065_, _40064_, _40039_);
  or _47616_ (_40066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39831_);
  or _47617_ (_40067_, _40066_, _40041_);
  and _47618_ (_40068_, _40067_, _40010_);
  and _47619_ (_40069_, _40068_, _40065_);
  and _47620_ (_40070_, _39899_, _39842_);
  or _47621_ (_40071_, _40070_, _40069_);
  and _47622_ (_40072_, _40071_, _39914_);
  and _47623_ (_40073_, _40049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _47624_ (_40074_, _40073_, _40051_);
  or _47625_ (_40075_, _40066_, _40053_);
  and _47626_ (_40076_, _40075_, _40004_);
  and _47627_ (_40077_, _40076_, _40074_);
  and _47628_ (_40078_, _39921_, _39842_);
  or _47629_ (_40079_, _40078_, _40077_);
  and _47630_ (_40080_, _40079_, _39950_);
  or _47631_ (_40081_, _40080_, _40072_);
  and _47632_ (_40082_, _40081_, _39962_);
  or _47633_ (_40083_, _40082_, _40063_);
  and _47634_ (_42746_, _40083_, _41806_);
  and _47635_ (_40084_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not _47636_ (_40085_, _39940_);
  and _47637_ (_40086_, _40085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _47638_ (_40087_, _39904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47639_ (_40088_, _40087_, _39901_);
  or _47640_ (_40089_, _40088_, _40086_);
  or _47641_ (_40090_, _40041_, _39832_);
  and _47642_ (_40091_, _40090_, _40089_);
  or _47643_ (_40092_, _40091_, _39899_);
  or _47644_ (_40093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47645_ (_40094_, _40093_, _40010_);
  and _47646_ (_40095_, _40094_, _39914_);
  and _47647_ (_40096_, _40095_, _40092_);
  not _47648_ (_40097_, _39951_);
  and _47649_ (_40098_, _40097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _47650_ (_40099_, _39954_, _39923_);
  or _47651_ (_40100_, _40099_, _40098_);
  or _47652_ (_40101_, _40053_, _39832_);
  and _47653_ (_40102_, _40101_, _40004_);
  and _47654_ (_40103_, _40102_, _40100_);
  and _47655_ (_40104_, _40093_, _39921_);
  or _47656_ (_40105_, _40104_, _40103_);
  and _47657_ (_40106_, _40105_, _39950_);
  or _47658_ (_40107_, _40106_, _40096_);
  and _47659_ (_40108_, _40107_, _39962_);
  or _47660_ (_40109_, _40108_, _40084_);
  and _47661_ (_42748_, _40109_, _41806_);
  and _47662_ (_40110_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _47663_ (_40111_, _40085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _47664_ (_40112_, _40111_, _40088_);
  or _47665_ (_40113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47666_ (_40114_, _40113_, _40041_);
  and _47667_ (_40115_, _40114_, _40010_);
  and _47668_ (_40116_, _40115_, _40112_);
  and _47669_ (_40117_, _39899_, _39841_);
  or _47670_ (_40118_, _40117_, _40116_);
  and _47671_ (_40119_, _40118_, _39914_);
  and _47672_ (_40120_, _40097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _47673_ (_40121_, _40120_, _40099_);
  or _47674_ (_40122_, _40113_, _40053_);
  and _47675_ (_40123_, _40122_, _40004_);
  and _47676_ (_40124_, _40123_, _40121_);
  and _47677_ (_40125_, _39921_, _39841_);
  or _47678_ (_40126_, _40125_, _40124_);
  and _47679_ (_40127_, _40126_, _39950_);
  or _47680_ (_40128_, _40127_, _40119_);
  and _47681_ (_40129_, _40128_, _39962_);
  or _47682_ (_40130_, _40129_, _40110_);
  and _47683_ (_42750_, _40130_, _41806_);
  and _47684_ (_40131_, _39935_, _39914_);
  nand _47685_ (_40132_, _39935_, _39931_);
  and _47686_ (_40133_, _40132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _47687_ (_40134_, _40133_, _40131_);
  and _47688_ (_42752_, _40134_, _41806_);
  and _47689_ (_40135_, _39932_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _47690_ (_40136_, _40135_, _39917_);
  and _47691_ (_42754_, _40136_, _41806_);
  and _47692_ (_40137_, _39819_, _24456_);
  or _47693_ (_40138_, _40137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _47694_ (_40139_, _40138_, _39828_);
  nand _47695_ (_40140_, _40137_, _28676_);
  and _47696_ (_40141_, _40140_, _40139_);
  nor _47697_ (_40142_, _39828_, _38425_);
  or _47698_ (_40143_, _40142_, _40141_);
  and _47699_ (_42756_, _40143_, _41806_);
  and _47700_ (_40144_, _39819_, _30708_);
  nand _47701_ (_40145_, _40144_, _28676_);
  or _47702_ (_40146_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _47703_ (_40147_, _40146_, _39828_);
  and _47704_ (_40148_, _40147_, _40145_);
  nor _47705_ (_40149_, _39828_, _38410_);
  or _47706_ (_40150_, _40149_, _40148_);
  and _47707_ (_42758_, _40150_, _41806_);
  and _47708_ (_40151_, _39819_, _32131_);
  nand _47709_ (_40152_, _40151_, _28676_);
  or _47710_ (_40153_, _40151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _47711_ (_40154_, _40153_, _39828_);
  and _47712_ (_40155_, _40154_, _40152_);
  nor _47713_ (_40156_, _39828_, _38394_);
  or _47714_ (_40157_, _40156_, _40155_);
  and _47715_ (_42760_, _40157_, _41806_);
  and _47716_ (_40158_, _39808_, _24456_);
  nand _47717_ (_40159_, _40158_, _28676_);
  not _47718_ (_40160_, _39805_);
  or _47719_ (_40161_, _40158_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47720_ (_40162_, _40161_, _40160_);
  and _47721_ (_40163_, _40162_, _40159_);
  nor _47722_ (_40164_, _40160_, _38425_);
  or _47723_ (_40165_, _40164_, _40163_);
  and _47724_ (_42762_, _40165_, _41806_);
  and _47725_ (_40166_, _39808_, _30002_);
  nand _47726_ (_40167_, _40166_, _28676_);
  or _47727_ (_40168_, _40166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _47728_ (_40169_, _40168_, _40160_);
  and _47729_ (_40170_, _40169_, _40167_);
  nor _47730_ (_40171_, _40160_, _38417_);
  or _47731_ (_40172_, _40171_, _40170_);
  and _47732_ (_42764_, _40172_, _41806_);
  and _47733_ (_40173_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _47734_ (_40174_, _40173_, _30719_);
  and _47735_ (_40175_, _40174_, _39808_);
  nand _47736_ (_40176_, _39808_, _39426_);
  and _47737_ (_40177_, _40176_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _47738_ (_40178_, _40177_, _39805_);
  or _47739_ (_40179_, _40178_, _40175_);
  nand _47740_ (_40180_, _39805_, _38410_);
  and _47741_ (_40181_, _40180_, _41806_);
  and _47742_ (_42766_, _40181_, _40179_);
  and _47743_ (_40182_, _39808_, _31436_);
  nand _47744_ (_40183_, _40182_, _28676_);
  or _47745_ (_40184_, _40182_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _47746_ (_40185_, _40184_, _40183_);
  or _47747_ (_40186_, _40185_, _39805_);
  nand _47748_ (_40187_, _39805_, _38402_);
  and _47749_ (_40188_, _40187_, _41806_);
  and _47750_ (_42768_, _40188_, _40186_);
  and _47751_ (_40189_, _39808_, _32131_);
  nand _47752_ (_40190_, _40189_, _28676_);
  or _47753_ (_40191_, _40189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _47754_ (_40192_, _40191_, _40160_);
  and _47755_ (_40193_, _40192_, _40190_);
  nor _47756_ (_40194_, _40160_, _38394_);
  or _47757_ (_40195_, _40194_, _40193_);
  and _47758_ (_42770_, _40195_, _41806_);
  and _47759_ (_40196_, _39808_, _32941_);
  nand _47760_ (_40197_, _40196_, _28676_);
  or _47761_ (_40198_, _40196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _47762_ (_40199_, _40198_, _40160_);
  and _47763_ (_40200_, _40199_, _40197_);
  nor _47764_ (_40201_, _40160_, _38366_);
  or _47765_ (_40202_, _40201_, _40200_);
  and _47766_ (_42772_, _40202_, _41806_);
  and _47767_ (_40203_, _39808_, _33697_);
  nand _47768_ (_40204_, _40203_, _28676_);
  or _47769_ (_40205_, _40203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _47770_ (_40206_, _40205_, _40160_);
  and _47771_ (_40207_, _40206_, _40204_);
  nor _47772_ (_40208_, _40160_, _38280_);
  or _47773_ (_40209_, _40208_, _40207_);
  and _47774_ (_42774_, _40209_, _41806_);
  and _47775_ (_40210_, _39797_, _24456_);
  nand _47776_ (_40211_, _40210_, _28676_);
  or _47777_ (_40212_, _40210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47778_ (_40213_, _40212_, _40211_);
  or _47779_ (_40214_, _40213_, _39794_);
  nand _47780_ (_40215_, _39794_, _38425_);
  and _47781_ (_40216_, _40215_, _41806_);
  and _47782_ (_42776_, _40216_, _40214_);
  and _47783_ (_40217_, _39797_, _30002_);
  nand _47784_ (_40218_, _40217_, _28676_);
  not _47785_ (_40219_, _39794_);
  or _47786_ (_40220_, _40217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47787_ (_40221_, _40220_, _40219_);
  and _47788_ (_40222_, _40221_, _40218_);
  nor _47789_ (_40223_, _40219_, _38417_);
  or _47790_ (_40224_, _40223_, _40222_);
  and _47791_ (_42778_, _40224_, _41806_);
  and _47792_ (_40225_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _47793_ (_40226_, _40225_, _30719_);
  and _47794_ (_40227_, _40226_, _39797_);
  nand _47795_ (_40228_, _39797_, _39426_);
  and _47796_ (_40229_, _40228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _47797_ (_40230_, _40229_, _39794_);
  or _47798_ (_40231_, _40230_, _40227_);
  nand _47799_ (_40232_, _39794_, _38410_);
  and _47800_ (_40233_, _40232_, _41806_);
  and _47801_ (_42780_, _40233_, _40231_);
  and _47802_ (_40234_, _39797_, _31436_);
  nand _47803_ (_40235_, _40234_, _28676_);
  or _47804_ (_40236_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _47805_ (_40237_, _40236_, _40219_);
  and _47806_ (_40238_, _40237_, _40235_);
  nor _47807_ (_40239_, _40219_, _38402_);
  or _47808_ (_40240_, _40239_, _40238_);
  and _47809_ (_42782_, _40240_, _41806_);
  and _47810_ (_40241_, _39797_, _32131_);
  nand _47811_ (_40242_, _40241_, _28676_);
  or _47812_ (_40243_, _40241_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _47813_ (_40244_, _40243_, _40219_);
  and _47814_ (_40245_, _40244_, _40242_);
  nor _47815_ (_40246_, _40219_, _38394_);
  or _47816_ (_40247_, _40246_, _40245_);
  and _47817_ (_42784_, _40247_, _41806_);
  and _47818_ (_40248_, _39797_, _32941_);
  nand _47819_ (_40249_, _40248_, _28676_);
  or _47820_ (_40250_, _40248_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _47821_ (_40251_, _40250_, _40219_);
  and _47822_ (_40252_, _40251_, _40249_);
  nor _47823_ (_40253_, _40219_, _38366_);
  or _47824_ (_40254_, _40253_, _40252_);
  and _47825_ (_42786_, _40254_, _41806_);
  and _47826_ (_40255_, _39797_, _33697_);
  nand _47827_ (_40256_, _40255_, _28676_);
  or _47828_ (_40257_, _40255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _47829_ (_40258_, _40257_, _40219_);
  and _47830_ (_40259_, _40258_, _40256_);
  nor _47831_ (_40260_, _40219_, _38280_);
  or _47832_ (_40261_, _40260_, _40259_);
  and _47833_ (_42788_, _40261_, _41806_);
  nor _47834_ (_40262_, _24949_, _23932_);
  nor _47835_ (_40263_, _40262_, _28065_);
  not _47836_ (_40264_, _40263_);
  and _47837_ (_40265_, _37954_, _37811_);
  not _47838_ (_40266_, _38443_);
  and _47839_ (_40267_, _40266_, _40265_);
  not _47840_ (_40268_, _40267_);
  not _47841_ (_40269_, _36836_);
  and _47842_ (_40270_, _37800_, _40269_);
  and _47843_ (_40271_, _40270_, _37954_);
  not _47844_ (_40272_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _47845_ (_40273_, _36409_, _29980_);
  nor _47846_ (_40274_, _36409_, _29980_);
  nor _47847_ (_40275_, _40274_, _40273_);
  and _47848_ (_40276_, _40275_, _24313_);
  not _47849_ (_40277_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _47850_ (_40278_, _38821_, _40277_);
  nor _47851_ (_40279_, _40278_, _38908_);
  and _47852_ (_40280_, _40279_, _25113_);
  nor _47853_ (_40281_, _40279_, _25113_);
  nor _47854_ (_40282_, _40281_, _40280_);
  and _47855_ (_40283_, _40282_, _24197_);
  and _47856_ (_40284_, _40283_, _40276_);
  and _47857_ (_40285_, _40284_, _40263_);
  and _47858_ (_40286_, _40285_, _40272_);
  and _47859_ (_40287_, _40286_, _38173_);
  and _47860_ (_40288_, _40279_, _36420_);
  and _47861_ (_40289_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _47862_ (_40290_, _40279_, _36420_);
  and _47863_ (_40291_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor _47864_ (_40292_, _40291_, _40289_);
  nor _47865_ (_40293_, _40279_, _36409_);
  and _47866_ (_40294_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _47867_ (_40295_, _40279_, _36409_);
  and _47868_ (_40296_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _47869_ (_40297_, _40296_, _40294_);
  and _47870_ (_40298_, _40297_, _40292_);
  nor _47871_ (_40299_, _40298_, _40286_);
  nor _47872_ (_40300_, _40299_, _40287_);
  not _47873_ (_40301_, _40300_);
  and _47874_ (_40302_, _40301_, _40271_);
  not _47875_ (_40303_, _37954_);
  nor _47876_ (_40304_, _37800_, _40269_);
  not _47877_ (_40305_, _33860_);
  and _47878_ (_40306_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _47879_ (_40307_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _47880_ (_40308_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _47881_ (_40309_, _40308_, _40307_);
  and _47882_ (_40310_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _47883_ (_40311_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _47884_ (_40312_, _40311_, _40310_);
  and _47885_ (_40313_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _47886_ (_40314_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _47887_ (_40315_, _40314_, _40313_);
  and _47888_ (_40316_, _40315_, _40312_);
  and _47889_ (_40317_, _40316_, _40309_);
  nor _47890_ (_40318_, _33915_, _40305_);
  not _47891_ (_40319_, _40318_);
  nor _47892_ (_40320_, _40319_, _40317_);
  nor _47893_ (_40321_, _40320_, _40306_);
  not _47894_ (_40322_, _40321_);
  and _47895_ (_40323_, _40322_, _40304_);
  nor _47896_ (_40324_, _40323_, _40303_);
  not _47897_ (_40325_, _40324_);
  nor _47898_ (_40326_, _40325_, _40302_);
  and _47899_ (_40327_, _40326_, _40268_);
  nor _47900_ (_40328_, _37384_, _37148_);
  nor _47901_ (_40329_, _37296_, _37252_);
  nor _47902_ (_40330_, _37454_, _37219_);
  and _47903_ (_40331_, _40330_, _40329_);
  and _47904_ (_40332_, _37539_, _37351_);
  and _47905_ (_40333_, _40332_, _40331_);
  and _47906_ (_40334_, _40333_, _40328_);
  nor _47907_ (_40335_, _40334_, _33817_);
  and _47908_ (_40336_, _37507_, _36584_);
  nor _47909_ (_40337_, _37712_, _40336_);
  nor _47910_ (_40338_, _40337_, _37679_);
  nor _47911_ (_40339_, _40338_, _40335_);
  not _47912_ (_40340_, _40339_);
  and _47913_ (_40341_, _40340_, _40327_);
  and _47914_ (_40342_, _40304_, _37954_);
  and _47915_ (_40343_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _47916_ (_40344_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _47917_ (_40345_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _47918_ (_40346_, _40345_, _40344_);
  and _47919_ (_40347_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _47920_ (_40348_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _47921_ (_40349_, _40348_, _40347_);
  and _47922_ (_40350_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _47923_ (_40351_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _47924_ (_40352_, _40351_, _40350_);
  and _47925_ (_40353_, _40352_, _40349_);
  and _47926_ (_40354_, _40353_, _40346_);
  nor _47927_ (_40355_, _40354_, _40319_);
  nor _47928_ (_40356_, _40355_, _40343_);
  not _47929_ (_40357_, _40356_);
  and _47930_ (_40358_, _40357_, _40342_);
  not _47931_ (_40359_, _40271_);
  not _47932_ (_40360_, _38402_);
  and _47933_ (_40361_, _40286_, _40360_);
  and _47934_ (_40362_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _47935_ (_40363_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _47936_ (_40364_, _40363_, _40362_);
  and _47937_ (_40365_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _47938_ (_40366_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _47939_ (_40367_, _40366_, _40365_);
  and _47940_ (_40368_, _40367_, _40364_);
  nor _47941_ (_40369_, _40368_, _40286_);
  nor _47942_ (_40370_, _40369_, _40361_);
  nor _47943_ (_40371_, _40370_, _40359_);
  nor _47944_ (_40372_, _40371_, _40358_);
  not _47945_ (_40373_, _38469_);
  and _47946_ (_40374_, _40373_, _40265_);
  not _47947_ (_40375_, _40279_);
  and _47948_ (_40376_, _37800_, _36836_);
  and _47949_ (_40377_, _40376_, _37954_);
  and _47950_ (_40378_, _40377_, _40375_);
  nor _47951_ (_40379_, _40378_, _40374_);
  and _47952_ (_40380_, _40379_, _40372_);
  not _47953_ (_40381_, _40380_);
  and _47954_ (_40382_, _40381_, _40341_);
  and _47955_ (_40383_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _47956_ (_40384_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _47957_ (_40385_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _47958_ (_40386_, _40385_, _40384_);
  and _47959_ (_40387_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _47960_ (_40388_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _47961_ (_40389_, _40388_, _40387_);
  and _47962_ (_40390_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _47963_ (_40391_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _47964_ (_40392_, _40391_, _40390_);
  and _47965_ (_40393_, _40392_, _40389_);
  and _47966_ (_40394_, _40393_, _40386_);
  nor _47967_ (_40395_, _40394_, _40319_);
  nor _47968_ (_40396_, _40395_, _40383_);
  not _47969_ (_40397_, _40396_);
  and _47970_ (_40398_, _40397_, _40342_);
  and _47971_ (_40399_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and _47972_ (_40400_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _47973_ (_40401_, _40400_, _40399_);
  and _47974_ (_40402_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _47975_ (_40403_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _47976_ (_40404_, _40403_, _40402_);
  and _47977_ (_40405_, _40404_, _40401_);
  nor _47978_ (_40406_, _40405_, _40286_);
  and _47979_ (_40407_, _40286_, _38426_);
  nor _47980_ (_40408_, _40407_, _40406_);
  nor _47981_ (_40409_, _40408_, _40359_);
  nor _47982_ (_40410_, _40409_, _40398_);
  not _47983_ (_40411_, _38451_);
  and _47984_ (_40412_, _40411_, _40265_);
  and _47985_ (_40413_, _40377_, _36420_);
  nor _47986_ (_40414_, _40413_, _40412_);
  and _47987_ (_40415_, _40414_, _40410_);
  nor _47988_ (_40416_, _40415_, _40340_);
  nor _47989_ (_40417_, _40416_, _40382_);
  and _47990_ (_40418_, _24949_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _47991_ (_40419_, _40418_, _25113_);
  nor _47992_ (_40420_, _24434_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _47993_ (_40421_, _40420_, _40419_);
  not _47994_ (_40422_, _40421_);
  and _47995_ (_40423_, _40422_, _40417_);
  nor _47996_ (_40424_, _40423_, _40264_);
  and _47997_ (_40425_, _40303_, _36836_);
  and _47998_ (_40426_, _40425_, _37800_);
  not _47999_ (_40427_, _38481_);
  and _48000_ (_40428_, _40427_, _40265_);
  nor _48001_ (_40429_, _40428_, _40426_);
  and _48002_ (_40430_, _40303_, _37811_);
  not _48003_ (_40431_, _40430_);
  not _48004_ (_40432_, _38366_);
  and _48005_ (_40433_, _40286_, _40432_);
  and _48006_ (_40434_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _48007_ (_40435_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _48008_ (_40436_, _40435_, _40434_);
  and _48009_ (_40437_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _48010_ (_40438_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _48011_ (_40439_, _40438_, _40437_);
  and _48012_ (_40440_, _40439_, _40436_);
  nor _48013_ (_40441_, _40440_, _40286_);
  nor _48014_ (_40442_, _40441_, _40433_);
  not _48015_ (_40443_, _40442_);
  and _48016_ (_40444_, _40443_, _40271_);
  and _48017_ (_40445_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _48018_ (_40446_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _48019_ (_40447_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _48020_ (_40448_, _40447_, _40446_);
  and _48021_ (_40449_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _48022_ (_40450_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _48023_ (_40451_, _40450_, _40449_);
  and _48024_ (_40452_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _48025_ (_40453_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _48026_ (_40454_, _40453_, _40452_);
  and _48027_ (_40455_, _40454_, _40451_);
  and _48028_ (_40456_, _40455_, _40448_);
  nor _48029_ (_40457_, _40456_, _40319_);
  nor _48030_ (_40458_, _40457_, _40445_);
  not _48031_ (_40459_, _40458_);
  and _48032_ (_40460_, _40459_, _40342_);
  nor _48033_ (_40461_, _40460_, _40444_);
  and _48034_ (_40462_, _40461_, _40431_);
  and _48035_ (_40463_, _40462_, _40429_);
  not _48036_ (_40464_, _40463_);
  and _48037_ (_40465_, _40464_, _40341_);
  and _48038_ (_40466_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _48039_ (_40467_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _48040_ (_40468_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _48041_ (_40469_, _40468_, _40467_);
  and _48042_ (_40470_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _48043_ (_40471_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _48044_ (_40472_, _40471_, _40470_);
  and _48045_ (_40473_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _48046_ (_40474_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _48047_ (_40475_, _40474_, _40473_);
  and _48048_ (_40476_, _40475_, _40472_);
  and _48049_ (_40477_, _40476_, _40469_);
  nor _48050_ (_40478_, _40477_, _40319_);
  nor _48051_ (_40479_, _40478_, _40466_);
  not _48052_ (_40480_, _40479_);
  and _48053_ (_40481_, _40480_, _40342_);
  not _48054_ (_40482_, _38410_);
  and _48055_ (_40483_, _40286_, _40482_);
  and _48056_ (_40484_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _48057_ (_40485_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _48058_ (_40486_, _40485_, _40484_);
  and _48059_ (_40487_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _48060_ (_40488_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _48061_ (_40489_, _40488_, _40487_);
  and _48062_ (_40490_, _40489_, _40486_);
  nor _48063_ (_40491_, _40490_, _40286_);
  nor _48064_ (_40492_, _40491_, _40483_);
  not _48065_ (_40493_, _40492_);
  and _48066_ (_40494_, _40493_, _40271_);
  nor _48067_ (_40495_, _40494_, _40481_);
  not _48068_ (_40496_, _38463_);
  and _48069_ (_40497_, _40496_, _40265_);
  and _48070_ (_40498_, _40377_, _36869_);
  nor _48071_ (_40499_, _40498_, _40497_);
  and _48072_ (_40500_, _40499_, _40495_);
  nor _48073_ (_40501_, _40500_, _40340_);
  nor _48074_ (_40502_, _40501_, _40465_);
  and _48075_ (_40503_, _40418_, _39027_);
  nor _48076_ (_40504_, _24197_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _48077_ (_40505_, _40504_, _40503_);
  not _48078_ (_40506_, _40505_);
  and _48079_ (_40507_, _40506_, _40502_);
  nor _48080_ (_40508_, _40422_, _40417_);
  nor _48081_ (_40509_, _40508_, _40507_);
  and _48082_ (_40510_, _40509_, _40424_);
  not _48083_ (_40511_, _38475_);
  and _48084_ (_40512_, _40511_, _40265_);
  or _48085_ (_40513_, _40512_, _40425_);
  and _48086_ (_40514_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _48087_ (_40515_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _48088_ (_40516_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _48089_ (_40517_, _40516_, _40515_);
  and _48090_ (_40518_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _48091_ (_40519_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _48092_ (_40520_, _40519_, _40518_);
  and _48093_ (_40521_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _48094_ (_40522_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _48095_ (_40523_, _40522_, _40521_);
  and _48096_ (_40524_, _40523_, _40520_);
  and _48097_ (_40525_, _40524_, _40517_);
  nor _48098_ (_40526_, _40525_, _40319_);
  nor _48099_ (_40527_, _40526_, _40514_);
  not _48100_ (_40528_, _40527_);
  and _48101_ (_40529_, _40528_, _40342_);
  and _48102_ (_40530_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and _48103_ (_40531_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and _48104_ (_40532_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _48105_ (_40533_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _48106_ (_40534_, _40533_, _40532_);
  or _48107_ (_40535_, _40534_, _40531_);
  nor _48108_ (_40536_, _40535_, _40530_);
  nor _48109_ (_40537_, _40536_, _40286_);
  not _48110_ (_40538_, _38394_);
  and _48111_ (_40539_, _40286_, _40538_);
  or _48112_ (_40540_, _40539_, _40537_);
  and _48113_ (_40541_, _40540_, _40271_);
  or _48114_ (_40542_, _40541_, _40529_);
  nor _48115_ (_40543_, _38821_, _38949_);
  or _48116_ (_40544_, _40543_, _38963_);
  and _48117_ (_40545_, _40544_, _40377_);
  or _48118_ (_40546_, _40545_, _40542_);
  or _48119_ (_40547_, _40546_, _40513_);
  and _48120_ (_40548_, _40547_, _40341_);
  and _48121_ (_40549_, _40270_, _40303_);
  not _48122_ (_40550_, _38457_);
  and _48123_ (_40551_, _40550_, _40265_);
  nor _48124_ (_40552_, _40551_, _40549_);
  and _48125_ (_40553_, _40377_, _36431_);
  and _48126_ (_40554_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  not _48127_ (_40555_, _40554_);
  and _48128_ (_40556_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _48129_ (_40557_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _48130_ (_40558_, _40557_, _40556_);
  and _48131_ (_40559_, _40558_, _40555_);
  and _48132_ (_40560_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _48133_ (_40561_, _40560_, _40286_);
  and _48134_ (_40562_, _40561_, _40559_);
  and _48135_ (_40563_, _40286_, _38417_);
  or _48136_ (_40564_, _40563_, _40562_);
  nor _48137_ (_40570_, _40564_, _40359_);
  and _48138_ (_40576_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _48139_ (_40582_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _48140_ (_40588_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _48141_ (_40594_, _40588_, _40582_);
  and _48142_ (_40597_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _48143_ (_40598_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _48144_ (_40599_, _40598_, _40597_);
  and _48145_ (_40600_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _48146_ (_40601_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _48147_ (_40602_, _40601_, _40600_);
  and _48148_ (_40603_, _40602_, _40599_);
  and _48149_ (_40604_, _40603_, _40594_);
  nor _48150_ (_40605_, _40604_, _40319_);
  nor _48151_ (_40606_, _40605_, _40576_);
  not _48152_ (_40607_, _40606_);
  and _48153_ (_40608_, _40607_, _40342_);
  or _48154_ (_40609_, _40608_, _40570_);
  nor _48155_ (_40610_, _40609_, _40553_);
  and _48156_ (_40611_, _40610_, _40552_);
  nor _48157_ (_40612_, _40611_, _40340_);
  nor _48158_ (_40613_, _40612_, _40548_);
  not _48159_ (_40614_, _25244_);
  and _48160_ (_40615_, _40418_, _40614_);
  nor _48161_ (_40616_, _24313_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _48162_ (_40617_, _40616_, _40615_);
  nand _48163_ (_40618_, _40617_, _40613_);
  or _48164_ (_40619_, _40617_, _40613_);
  and _48165_ (_40620_, _40619_, _40618_);
  not _48166_ (_40621_, _40620_);
  nor _48167_ (_40622_, _40506_, _40502_);
  not _48168_ (_40623_, _40622_);
  nor _48169_ (_40624_, _40381_, _40341_);
  and _48170_ (_40625_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _48171_ (_40626_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _48172_ (_40627_, _40626_, _40625_);
  and _48173_ (_40628_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _48174_ (_40629_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _48175_ (_40630_, _40629_, _40628_);
  and _48176_ (_40631_, _40630_, _40627_);
  nor _48177_ (_40632_, _40631_, _40286_);
  not _48178_ (_40633_, _38280_);
  and _48179_ (_40636_, _40286_, _40633_);
  nor _48180_ (_40639_, _40636_, _40632_);
  nor _48181_ (_40643_, _40639_, _40359_);
  and _48182_ (_40645_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _48183_ (_40646_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _48184_ (_40647_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _48185_ (_40652_, _40647_, _40646_);
  and _48186_ (_40657_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _48187_ (_40658_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _48188_ (_40659_, _40658_, _40657_);
  and _48189_ (_40660_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _48190_ (_40666_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _48191_ (_40670_, _40666_, _40660_);
  and _48192_ (_40671_, _40670_, _40659_);
  and _48193_ (_40672_, _40671_, _40652_);
  nor _48194_ (_40677_, _40672_, _40319_);
  nor _48195_ (_40682_, _40677_, _40645_);
  not _48196_ (_40683_, _40682_);
  and _48197_ (_40684_, _40683_, _40304_);
  or _48198_ (_40685_, _40684_, _40425_);
  nor _48199_ (_40691_, _40685_, _40643_);
  not _48200_ (_40695_, _38487_);
  and _48201_ (_40696_, _40695_, _40265_);
  nor _48202_ (_40697_, _40696_, _40430_);
  and _48203_ (_40703_, _40697_, _40691_);
  and _48204_ (_40707_, _40703_, _40341_);
  nor _48205_ (_40708_, _40707_, _40624_);
  nor _48206_ (_40709_, _40418_, _25113_);
  and _48207_ (_40714_, _40418_, _24665_);
  nor _48208_ (_40719_, _40714_, _40709_);
  not _48209_ (_40720_, _40719_);
  and _48210_ (_40721_, _40720_, _40708_);
  nor _48211_ (_40726_, _40720_, _40708_);
  nor _48212_ (_40731_, _40726_, _40721_);
  and _48213_ (_40732_, _40731_, _40623_);
  and _48214_ (_40733_, _40732_, _40621_);
  and _48215_ (_40734_, _40733_, _40510_);
  not _48216_ (_40740_, _40502_);
  and _48217_ (_40744_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not _48218_ (_40745_, _40417_);
  and _48219_ (_40746_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _48220_ (_40752_, _40746_, _40744_);
  and _48221_ (_40756_, _40752_, _40613_);
  not _48222_ (_40757_, _40613_);
  not _48223_ (_40758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _48224_ (_40763_, _40417_, _40758_);
  and _48225_ (_40768_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _48226_ (_40769_, _40768_, _40763_);
  and _48227_ (_40770_, _40769_, _40757_);
  or _48228_ (_40775_, _40770_, _40756_);
  or _48229_ (_40780_, _40775_, _40740_);
  not _48230_ (_40781_, _40708_);
  and _48231_ (_40782_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and _48232_ (_40785_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _48233_ (_40791_, _40785_, _40782_);
  and _48234_ (_40793_, _40791_, _40613_);
  not _48235_ (_40794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _48236_ (_40797_, _40417_, _40794_);
  and _48237_ (_40803_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _48238_ (_40805_, _40803_, _40797_);
  and _48239_ (_40806_, _40805_, _40757_);
  or _48240_ (_40808_, _40806_, _40793_);
  or _48241_ (_40814_, _40808_, _40502_);
  and _48242_ (_40817_, _40814_, _40781_);
  and _48243_ (_40818_, _40817_, _40780_);
  or _48244_ (_40820_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _48245_ (_40826_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _48246_ (_40828_, _40826_, _40820_);
  and _48247_ (_40829_, _40828_, _40613_);
  or _48248_ (_40830_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not _48249_ (_40831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand _48250_ (_40832_, _40417_, _40831_);
  and _48251_ (_40833_, _40832_, _40830_);
  and _48252_ (_40834_, _40833_, _40757_);
  or _48253_ (_40835_, _40834_, _40829_);
  or _48254_ (_40836_, _40835_, _40740_);
  or _48255_ (_40837_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _48256_ (_40838_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _48257_ (_40839_, _40838_, _40837_);
  and _48258_ (_40840_, _40839_, _40613_);
  or _48259_ (_40841_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not _48260_ (_40842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand _48261_ (_40843_, _40417_, _40842_);
  and _48262_ (_40844_, _40843_, _40841_);
  and _48263_ (_40845_, _40844_, _40757_);
  or _48264_ (_40846_, _40845_, _40840_);
  or _48265_ (_40847_, _40846_, _40502_);
  and _48266_ (_40848_, _40847_, _40708_);
  and _48267_ (_40849_, _40848_, _40836_);
  or _48268_ (_40850_, _40849_, _40818_);
  or _48269_ (_40851_, _40850_, _40734_);
  not _48270_ (_40852_, _40734_);
  or _48271_ (_40853_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and _48272_ (_40854_, _40853_, _41806_);
  and _48273_ (_42863_, _40854_, _40851_);
  nor _48274_ (_40855_, _40421_, _40264_);
  nor _48275_ (_40856_, _40617_, _40264_);
  and _48276_ (_40857_, _40856_, _40855_);
  and _48277_ (_40858_, _40719_, _40263_);
  nor _48278_ (_40859_, _40505_, _40264_);
  and _48279_ (_40860_, _40859_, _40858_);
  and _48280_ (_40861_, _40860_, _40857_);
  and _48281_ (_40862_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _48282_ (_40863_, _40862_, _26071_);
  nor _48283_ (_40864_, _40863_, _28676_);
  nand _48284_ (_40865_, _26071_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48285_ (_40866_, _17475_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48286_ (_40867_, _40866_, _40865_);
  nor _48287_ (_40868_, _38162_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _48288_ (_40869_, _40868_, _40867_);
  or _48289_ (_40870_, _40869_, _40864_);
  and _48290_ (_40871_, _40870_, _40263_);
  and _48291_ (_40872_, _40871_, _40861_);
  not _48292_ (_40873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor _48293_ (_40874_, _40861_, _40873_);
  or _48294_ (_42875_, _40874_, _40872_);
  nor _48295_ (_40875_, _40859_, _40858_);
  nor _48296_ (_40876_, _40856_, _40855_);
  and _48297_ (_40877_, _40876_, _40263_);
  and _48298_ (_40878_, _40877_, _40875_);
  and _48299_ (_40879_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _26061_);
  and _48300_ (_40880_, _40879_, _26104_);
  not _48301_ (_40881_, _40880_);
  nor _48302_ (_40882_, _40881_, _28676_);
  not _48303_ (_40883_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48304_ (_40884_, _38425_, _40883_);
  or _48305_ (_40885_, _16315_, _40883_);
  and _48306_ (_40886_, _40885_, _40881_);
  and _48307_ (_40887_, _40886_, _40884_);
  or _48308_ (_40888_, _40887_, _40882_);
  and _48309_ (_40889_, _40888_, _40878_);
  not _48310_ (_40890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _48311_ (_40891_, _40878_, _40890_);
  or _48312_ (_43133_, _40891_, _40889_);
  nand _48313_ (_40892_, _40879_, _26180_);
  nor _48314_ (_40893_, _40892_, _28676_);
  nor _48315_ (_40894_, _38417_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48316_ (_40895_, _40879_, _26137_);
  and _48317_ (_40896_, _40879_, _26071_);
  or _48318_ (_40897_, _40896_, _40862_);
  or _48319_ (_40898_, _40897_, _40895_);
  and _48320_ (_40899_, _40898_, _17301_);
  or _48321_ (_40900_, _40899_, _40894_);
  or _48322_ (_40901_, _40900_, _40893_);
  and _48323_ (_40902_, _40901_, _40878_);
  not _48324_ (_40903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _48325_ (_40904_, _40878_, _40903_);
  or _48326_ (_43139_, _40904_, _40902_);
  not _48327_ (_40905_, _40878_);
  and _48328_ (_40906_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand _48329_ (_40907_, _40879_, _26147_);
  nor _48330_ (_40908_, _40907_, _28676_);
  nor _48331_ (_40909_, _38410_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48332_ (_40910_, _40879_, _26169_);
  or _48333_ (_40911_, _40910_, _40897_);
  and _48334_ (_40912_, _40911_, _15953_);
  or _48335_ (_40913_, _40912_, _40909_);
  or _48336_ (_40914_, _40913_, _40908_);
  and _48337_ (_40915_, _40914_, _40878_);
  or _48338_ (_43145_, _40915_, _40906_);
  and _48339_ (_40916_, _40896_, _29318_);
  nor _48340_ (_40917_, _38402_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _48341_ (_40918_, _40895_, _40862_);
  or _48342_ (_40919_, _40918_, _40910_);
  and _48343_ (_40920_, _40919_, _16985_);
  or _48344_ (_40921_, _40920_, _40917_);
  or _48345_ (_40922_, _40921_, _40916_);
  and _48346_ (_40923_, _40922_, _40878_);
  and _48347_ (_40924_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _48348_ (_43151_, _40924_, _40923_);
  nand _48349_ (_40925_, _40862_, _26104_);
  nor _48350_ (_40926_, _40925_, _28676_);
  nor _48351_ (_40927_, _38394_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48352_ (_40928_, _26104_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48353_ (_40929_, _16150_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48354_ (_40930_, _40929_, _40928_);
  or _48355_ (_40931_, _40930_, _40927_);
  or _48356_ (_40932_, _40931_, _40926_);
  and _48357_ (_40933_, _40932_, _40878_);
  and _48358_ (_40934_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _48359_ (_43157_, _40934_, _40933_);
  nand _48360_ (_40935_, _40862_, _26180_);
  nor _48361_ (_40936_, _40935_, _28676_);
  nor _48362_ (_40937_, _38366_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48363_ (_40938_, _26180_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48364_ (_40939_, _17138_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48365_ (_40940_, _40939_, _40938_);
  or _48366_ (_40941_, _40940_, _40937_);
  or _48367_ (_40942_, _40941_, _40936_);
  and _48368_ (_40943_, _40942_, _40878_);
  and _48369_ (_40944_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _48370_ (_43163_, _40944_, _40943_);
  nand _48371_ (_40945_, _40862_, _26147_);
  nor _48372_ (_40946_, _40945_, _28676_);
  nor _48373_ (_40947_, _38280_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48374_ (_40948_, _26147_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48375_ (_40949_, _16490_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48376_ (_40950_, _40949_, _40948_);
  or _48377_ (_40951_, _40950_, _40947_);
  or _48378_ (_40952_, _40951_, _40946_);
  and _48379_ (_40953_, _40952_, _40878_);
  and _48380_ (_40954_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _48381_ (_43169_, _40954_, _40953_);
  and _48382_ (_40955_, _40878_, _40870_);
  and _48383_ (_40956_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _48384_ (_43172_, _40956_, _40955_);
  and _48385_ (_40957_, _40888_, _40263_);
  and _48386_ (_40958_, _40855_, _40617_);
  and _48387_ (_40959_, _40958_, _40875_);
  and _48388_ (_40960_, _40959_, _40957_);
  not _48389_ (_40961_, _40959_);
  and _48390_ (_40962_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _48391_ (_43180_, _40962_, _40960_);
  and _48392_ (_40963_, _40901_, _40263_);
  and _48393_ (_40964_, _40959_, _40963_);
  and _48394_ (_40965_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _48395_ (_43184_, _40965_, _40964_);
  and _48396_ (_40966_, _40914_, _40263_);
  and _48397_ (_40967_, _40959_, _40966_);
  and _48398_ (_40968_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _48399_ (_43188_, _40968_, _40967_);
  and _48400_ (_40969_, _40922_, _40263_);
  and _48401_ (_40970_, _40959_, _40969_);
  and _48402_ (_40971_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _48403_ (_43192_, _40971_, _40970_);
  and _48404_ (_40972_, _40932_, _40263_);
  and _48405_ (_40973_, _40959_, _40972_);
  not _48406_ (_40974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _48407_ (_40975_, _40959_, _40974_);
  or _48408_ (_43196_, _40975_, _40973_);
  and _48409_ (_40976_, _40942_, _40263_);
  and _48410_ (_40977_, _40959_, _40976_);
  not _48411_ (_40978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _48412_ (_40979_, _40959_, _40978_);
  or _48413_ (_43200_, _40979_, _40977_);
  and _48414_ (_40980_, _40952_, _40263_);
  and _48415_ (_40981_, _40959_, _40980_);
  and _48416_ (_40982_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _48417_ (_43204_, _40982_, _40981_);
  and _48418_ (_40983_, _40959_, _40871_);
  and _48419_ (_40984_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _48420_ (_43207_, _40984_, _40983_);
  and _48421_ (_40985_, _40856_, _40421_);
  and _48422_ (_40986_, _40985_, _40875_);
  and _48423_ (_40987_, _40986_, _40957_);
  not _48424_ (_40988_, _40986_);
  and _48425_ (_40989_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _48426_ (_43215_, _40989_, _40987_);
  and _48427_ (_40990_, _40986_, _40963_);
  and _48428_ (_40991_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _48429_ (_43219_, _40991_, _40990_);
  and _48430_ (_40992_, _40986_, _40966_);
  not _48431_ (_40993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _48432_ (_40994_, _40986_, _40993_);
  or _48433_ (_43223_, _40994_, _40992_);
  and _48434_ (_40995_, _40986_, _40969_);
  and _48435_ (_40996_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _48436_ (_43227_, _40996_, _40995_);
  and _48437_ (_40997_, _40986_, _40972_);
  not _48438_ (_40998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _48439_ (_40999_, _40986_, _40998_);
  or _48440_ (_43231_, _40999_, _40997_);
  and _48441_ (_41000_, _40986_, _40976_);
  not _48442_ (_41001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _48443_ (_41002_, _40986_, _41001_);
  or _48444_ (_43235_, _41002_, _41000_);
  and _48445_ (_41003_, _40986_, _40980_);
  and _48446_ (_41004_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _48447_ (_43239_, _41004_, _41003_);
  and _48448_ (_41005_, _40986_, _40871_);
  not _48449_ (_41006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _48450_ (_41007_, _40986_, _41006_);
  or _48451_ (_43242_, _41007_, _41005_);
  and _48452_ (_41008_, _40875_, _40857_);
  and _48453_ (_41009_, _41008_, _40957_);
  not _48454_ (_41010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _48455_ (_41011_, _41008_, _41010_);
  or _48456_ (_43248_, _41011_, _41009_);
  and _48457_ (_41012_, _41008_, _40963_);
  not _48458_ (_41013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _48459_ (_41014_, _41008_, _41013_);
  or _48460_ (_43252_, _41014_, _41012_);
  and _48461_ (_41015_, _41008_, _40966_);
  not _48462_ (_41016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _48463_ (_41017_, _41008_, _41016_);
  or _48464_ (_43256_, _41017_, _41015_);
  and _48465_ (_41018_, _41008_, _40969_);
  not _48466_ (_41019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _48467_ (_41020_, _41008_, _41019_);
  or _48468_ (_43260_, _41020_, _41018_);
  and _48469_ (_41021_, _41008_, _40972_);
  not _48470_ (_41022_, _41008_);
  and _48471_ (_41023_, _41022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _48472_ (_43264_, _41023_, _41021_);
  and _48473_ (_41024_, _41008_, _40976_);
  and _48474_ (_41025_, _41022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _48475_ (_43268_, _41025_, _41024_);
  and _48476_ (_41026_, _41008_, _40980_);
  and _48477_ (_41027_, _41022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _48478_ (_43272_, _41027_, _41026_);
  and _48479_ (_41028_, _41008_, _40871_);
  nor _48480_ (_41029_, _41008_, _40758_);
  or _48481_ (_43275_, _41029_, _41028_);
  and _48482_ (_41030_, _40859_, _40720_);
  and _48483_ (_41031_, _41030_, _40876_);
  and _48484_ (_41032_, _41031_, _40957_);
  not _48485_ (_41033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _48486_ (_41034_, _41031_, _41033_);
  or _48487_ (_43283_, _41034_, _41032_);
  and _48488_ (_41035_, _41031_, _40963_);
  not _48489_ (_41036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _48490_ (_41037_, _41031_, _41036_);
  or _48491_ (_43287_, _41037_, _41035_);
  and _48492_ (_41038_, _41031_, _40966_);
  not _48493_ (_41039_, _41031_);
  and _48494_ (_41040_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _48495_ (_43291_, _41040_, _41038_);
  and _48496_ (_41041_, _41031_, _40969_);
  not _48497_ (_41042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _48498_ (_41043_, _41031_, _41042_);
  or _48499_ (_43295_, _41043_, _41041_);
  and _48500_ (_41044_, _41031_, _40972_);
  and _48501_ (_41045_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _48502_ (_43299_, _41045_, _41044_);
  and _48503_ (_41046_, _41031_, _40976_);
  and _48504_ (_41047_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _48505_ (_43303_, _41047_, _41046_);
  and _48506_ (_41048_, _41031_, _40980_);
  and _48507_ (_41049_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _48508_ (_43307_, _41049_, _41048_);
  and _48509_ (_41050_, _41031_, _40871_);
  and _48510_ (_41051_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _48511_ (_43310_, _41051_, _41050_);
  and _48512_ (_41052_, _41030_, _40958_);
  and _48513_ (_41053_, _41052_, _40957_);
  not _48514_ (_41054_, _41052_);
  and _48515_ (_41055_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _48516_ (_43315_, _41055_, _41053_);
  and _48517_ (_41056_, _41052_, _40963_);
  and _48518_ (_41057_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _48519_ (_43319_, _41057_, _41056_);
  and _48520_ (_41058_, _41052_, _40966_);
  and _48521_ (_41059_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _48522_ (_43322_, _41059_, _41058_);
  and _48523_ (_41060_, _41052_, _40969_);
  and _48524_ (_41061_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _48525_ (_43326_, _41061_, _41060_);
  and _48526_ (_41062_, _41052_, _40972_);
  not _48527_ (_41063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _48528_ (_41064_, _41052_, _41063_);
  or _48529_ (_43330_, _41064_, _41062_);
  and _48530_ (_41065_, _41052_, _40976_);
  not _48531_ (_41066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _48532_ (_41067_, _41052_, _41066_);
  or _48533_ (_43334_, _41067_, _41065_);
  and _48534_ (_41068_, _41052_, _40980_);
  not _48535_ (_41069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor _48536_ (_41070_, _41052_, _41069_);
  or _48537_ (_43338_, _41070_, _41068_);
  and _48538_ (_41071_, _41052_, _40871_);
  and _48539_ (_41072_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _48540_ (_43341_, _41072_, _41071_);
  and _48541_ (_41073_, _41030_, _40985_);
  and _48542_ (_41074_, _41073_, _40957_);
  not _48543_ (_41075_, _41073_);
  and _48544_ (_41076_, _41075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _48545_ (_43346_, _41076_, _41074_);
  and _48546_ (_41077_, _41073_, _40963_);
  and _48547_ (_41078_, _41075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _48548_ (_43350_, _41078_, _41077_);
  and _48549_ (_41079_, _41073_, _40966_);
  not _48550_ (_41080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _48551_ (_41081_, _41073_, _41080_);
  or _48552_ (_43354_, _41081_, _41079_);
  and _48553_ (_41082_, _41073_, _40969_);
  and _48554_ (_41083_, _41075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _48555_ (_43358_, _41083_, _41082_);
  and _48556_ (_41084_, _41073_, _40972_);
  not _48557_ (_41085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _48558_ (_41086_, _41073_, _41085_);
  or _48559_ (_43362_, _41086_, _41084_);
  and _48560_ (_41087_, _41073_, _40976_);
  not _48561_ (_41088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _48562_ (_41089_, _41073_, _41088_);
  or _48563_ (_43366_, _41089_, _41087_);
  and _48564_ (_41090_, _41073_, _40980_);
  not _48565_ (_41091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _48566_ (_41092_, _41073_, _41091_);
  or _48567_ (_43370_, _41092_, _41090_);
  and _48568_ (_41093_, _41073_, _40871_);
  not _48569_ (_41094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _48570_ (_41095_, _41073_, _41094_);
  or _48571_ (_43373_, _41095_, _41093_);
  and _48572_ (_41096_, _41030_, _40857_);
  and _48573_ (_41097_, _41096_, _40957_);
  not _48574_ (_41098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _48575_ (_41099_, _41096_, _41098_);
  or _48576_ (_43378_, _41099_, _41097_);
  and _48577_ (_41100_, _41096_, _40963_);
  not _48578_ (_41101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor _48579_ (_41102_, _41096_, _41101_);
  or _48580_ (_43382_, _41102_, _41100_);
  and _48581_ (_41103_, _41096_, _40966_);
  not _48582_ (_41104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _48583_ (_41105_, _41096_, _41104_);
  or _48584_ (_43386_, _41105_, _41103_);
  and _48585_ (_41106_, _41096_, _40969_);
  not _48586_ (_41107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor _48587_ (_41108_, _41096_, _41107_);
  or _48588_ (_43390_, _41108_, _41106_);
  and _48589_ (_41109_, _41096_, _40972_);
  not _48590_ (_41110_, _41096_);
  and _48591_ (_41111_, _41110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _48592_ (_43394_, _41111_, _41109_);
  and _48593_ (_41112_, _41096_, _40976_);
  and _48594_ (_41113_, _41110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _48595_ (_43398_, _41113_, _41112_);
  and _48596_ (_41114_, _41096_, _40980_);
  and _48597_ (_41115_, _41110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _48598_ (_43402_, _41115_, _41114_);
  and _48599_ (_41116_, _41096_, _40871_);
  nor _48600_ (_41117_, _41096_, _40794_);
  or _48601_ (_43405_, _41117_, _41116_);
  and _48602_ (_41118_, _40858_, _40505_);
  and _48603_ (_41119_, _41118_, _40876_);
  and _48604_ (_41120_, _41119_, _40957_);
  not _48605_ (_41121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _48606_ (_41122_, _41119_, _41121_);
  or _48607_ (_43413_, _41122_, _41120_);
  and _48608_ (_41123_, _41119_, _40963_);
  not _48609_ (_41124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _48610_ (_41125_, _41119_, _41124_);
  or _48611_ (_43417_, _41125_, _41123_);
  and _48612_ (_41126_, _41119_, _40966_);
  not _48613_ (_41127_, _41119_);
  and _48614_ (_41128_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _48615_ (_43421_, _41128_, _41126_);
  and _48616_ (_41129_, _41119_, _40969_);
  not _48617_ (_41130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _48618_ (_41131_, _41119_, _41130_);
  or _48619_ (_43425_, _41131_, _41129_);
  and _48620_ (_41132_, _41119_, _40972_);
  and _48621_ (_41133_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _48622_ (_43429_, _41133_, _41132_);
  and _48623_ (_41134_, _41119_, _40976_);
  and _48624_ (_41135_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _48625_ (_43433_, _41135_, _41134_);
  and _48626_ (_41136_, _41119_, _40980_);
  not _48627_ (_41137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _48628_ (_41138_, _41119_, _41137_);
  or _48629_ (_43437_, _41138_, _41136_);
  and _48630_ (_41139_, _41119_, _40871_);
  and _48631_ (_41140_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _48632_ (_43440_, _41140_, _41139_);
  and _48633_ (_41141_, _41118_, _40958_);
  and _48634_ (_41142_, _41141_, _40957_);
  not _48635_ (_41143_, _41141_);
  and _48636_ (_41144_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _48637_ (_43445_, _41144_, _41142_);
  and _48638_ (_41145_, _41141_, _40963_);
  and _48639_ (_41146_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _48640_ (_43449_, _41146_, _41145_);
  and _48641_ (_41147_, _41141_, _40966_);
  and _48642_ (_41148_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _48643_ (_43453_, _41148_, _41147_);
  and _48644_ (_41149_, _41141_, _40969_);
  and _48645_ (_41150_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _48646_ (_43457_, _41150_, _41149_);
  and _48647_ (_41151_, _41141_, _40972_);
  not _48648_ (_41152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _48649_ (_41153_, _41141_, _41152_);
  or _48650_ (_43461_, _41153_, _41151_);
  and _48651_ (_41154_, _41141_, _40976_);
  not _48652_ (_41155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor _48653_ (_41156_, _41141_, _41155_);
  or _48654_ (_43465_, _41156_, _41154_);
  and _48655_ (_41157_, _41141_, _40980_);
  and _48656_ (_41158_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _48657_ (_43469_, _41158_, _41157_);
  and _48658_ (_41159_, _41141_, _40871_);
  and _48659_ (_41160_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _48660_ (_43472_, _41160_, _41159_);
  and _48661_ (_41161_, _41118_, _40985_);
  and _48662_ (_41162_, _41161_, _40957_);
  not _48663_ (_41163_, _41161_);
  and _48664_ (_41164_, _41163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _48665_ (_43477_, _41164_, _41162_);
  and _48666_ (_41165_, _41161_, _40963_);
  and _48667_ (_41166_, _41163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _48668_ (_43484_, _41166_, _41165_);
  and _48669_ (_41167_, _41161_, _40966_);
  not _48670_ (_41168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor _48671_ (_41169_, _41161_, _41168_);
  or _48672_ (_43504_, _41169_, _41167_);
  and _48673_ (_41170_, _41161_, _40969_);
  not _48674_ (_41171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _48675_ (_41172_, _41161_, _41171_);
  or _48676_ (_43524_, _41172_, _41170_);
  and _48677_ (_41173_, _41161_, _40972_);
  not _48678_ (_41174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _48679_ (_41175_, _41161_, _41174_);
  or _48680_ (_43542_, _41175_, _41173_);
  and _48681_ (_41176_, _41161_, _40976_);
  not _48682_ (_41177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _48683_ (_41178_, _41161_, _41177_);
  or _48684_ (_43560_, _41178_, _41176_);
  and _48685_ (_41179_, _41161_, _40980_);
  not _48686_ (_41180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _48687_ (_41181_, _41161_, _41180_);
  or _48688_ (_43578_, _41181_, _41179_);
  and _48689_ (_41182_, _41161_, _40871_);
  nor _48690_ (_41183_, _41161_, _40831_);
  or _48691_ (_43593_, _41183_, _41182_);
  and _48692_ (_41184_, _41118_, _40857_);
  and _48693_ (_41185_, _41184_, _40957_);
  not _48694_ (_41186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _48695_ (_41187_, _41184_, _41186_);
  or _48696_ (_43617_, _41187_, _41185_);
  and _48697_ (_41188_, _41184_, _40963_);
  not _48698_ (_41189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _48699_ (_41190_, _41184_, _41189_);
  or _48700_ (_43637_, _41190_, _41188_);
  and _48701_ (_41191_, _41184_, _40966_);
  not _48702_ (_41192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _48703_ (_41193_, _41184_, _41192_);
  or _48704_ (_43657_, _41193_, _41191_);
  and _48705_ (_41194_, _41184_, _40969_);
  not _48706_ (_41195_, _41184_);
  and _48707_ (_41196_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _48708_ (_43669_, _41196_, _41194_);
  and _48709_ (_41197_, _41184_, _40972_);
  and _48710_ (_41198_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or _48711_ (_43694_, _41198_, _41197_);
  and _48712_ (_41199_, _41184_, _40976_);
  and _48713_ (_41200_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _48714_ (_43712_, _41200_, _41199_);
  and _48715_ (_41201_, _41184_, _40980_);
  and _48716_ (_41202_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _48717_ (_43723_, _41202_, _41201_);
  and _48718_ (_41203_, _41184_, _40871_);
  not _48719_ (_41204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _48720_ (_41205_, _41184_, _41204_);
  or _48721_ (_43726_, _41205_, _41203_);
  and _48722_ (_41206_, _40876_, _40860_);
  and _48723_ (_41208_, _41206_, _40957_);
  not _48724_ (_41210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _48725_ (_41212_, _41206_, _41210_);
  or _48726_ (_43732_, _41212_, _41208_);
  and _48727_ (_41215_, _41206_, _40963_);
  not _48728_ (_41217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _48729_ (_41219_, _41206_, _41217_);
  or _48730_ (_43736_, _41219_, _41215_);
  and _48731_ (_41222_, _41206_, _40966_);
  not _48732_ (_41224_, _41206_);
  and _48733_ (_41226_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _48734_ (_43740_, _41226_, _41222_);
  and _48735_ (_41229_, _41206_, _40969_);
  not _48736_ (_41231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _48737_ (_41233_, _41206_, _41231_);
  or _48738_ (_43744_, _41233_, _41229_);
  and _48739_ (_41236_, _41206_, _40972_);
  and _48740_ (_41238_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _48741_ (_43748_, _41238_, _41236_);
  and _48742_ (_41241_, _41206_, _40976_);
  and _48743_ (_41243_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _48744_ (_43752_, _41243_, _41241_);
  and _48745_ (_41246_, _41206_, _40980_);
  not _48746_ (_41248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _48747_ (_41250_, _41206_, _41248_);
  or _48748_ (_43756_, _41250_, _41246_);
  and _48749_ (_41253_, _41206_, _40871_);
  and _48750_ (_41255_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _48751_ (_43759_, _41255_, _41253_);
  and _48752_ (_41256_, _40958_, _40860_);
  and _48753_ (_41257_, _41256_, _40957_);
  not _48754_ (_41258_, _41256_);
  and _48755_ (_41259_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _48756_ (_43764_, _41259_, _41257_);
  and _48757_ (_41260_, _41256_, _40963_);
  and _48758_ (_41261_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _48759_ (_43768_, _41261_, _41260_);
  and _48760_ (_41262_, _41256_, _40966_);
  and _48761_ (_41263_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _48762_ (_43772_, _41263_, _41262_);
  and _48763_ (_41264_, _41256_, _40969_);
  and _48764_ (_41265_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _48765_ (_43776_, _41265_, _41264_);
  and _48766_ (_41266_, _41256_, _40972_);
  not _48767_ (_41267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _48768_ (_41268_, _41256_, _41267_);
  or _48769_ (_43780_, _41268_, _41266_);
  and _48770_ (_41269_, _41256_, _40976_);
  not _48771_ (_41270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor _48772_ (_41271_, _41256_, _41270_);
  or _48773_ (_43784_, _41271_, _41269_);
  and _48774_ (_41272_, _41256_, _40980_);
  and _48775_ (_41273_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _48776_ (_43788_, _41273_, _41272_);
  and _48777_ (_41274_, _41256_, _40871_);
  and _48778_ (_41275_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _48779_ (_43791_, _41275_, _41274_);
  and _48780_ (_41276_, _40985_, _40860_);
  and _48781_ (_41277_, _41276_, _40957_);
  not _48782_ (_41278_, _41276_);
  and _48783_ (_41279_, _41278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _48784_ (_43796_, _41279_, _41277_);
  and _48785_ (_41280_, _41276_, _40963_);
  and _48786_ (_41281_, _41278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _48787_ (_43800_, _41281_, _41280_);
  and _48788_ (_41282_, _41276_, _40966_);
  not _48789_ (_41283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _48790_ (_41284_, _41276_, _41283_);
  or _48791_ (_43804_, _41284_, _41282_);
  and _48792_ (_41285_, _41276_, _40969_);
  not _48793_ (_41286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _48794_ (_41287_, _41276_, _41286_);
  or _48795_ (_43808_, _41287_, _41285_);
  and _48796_ (_41288_, _41276_, _40972_);
  not _48797_ (_41289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _48798_ (_41290_, _41276_, _41289_);
  or _48799_ (_43812_, _41290_, _41288_);
  and _48800_ (_41291_, _41276_, _40976_);
  not _48801_ (_41292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _48802_ (_41293_, _41276_, _41292_);
  or _48803_ (_43816_, _41293_, _41291_);
  and _48804_ (_41294_, _41276_, _40980_);
  not _48805_ (_41295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _48806_ (_41296_, _41276_, _41295_);
  or _48807_ (_43820_, _41296_, _41294_);
  and _48808_ (_41297_, _41276_, _40871_);
  nor _48809_ (_41298_, _41276_, _40842_);
  or _48810_ (_43823_, _41298_, _41297_);
  and _48811_ (_41299_, _40957_, _40861_);
  not _48812_ (_41300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor _48813_ (_41301_, _40861_, _41300_);
  or _48814_ (_43826_, _41301_, _41299_);
  and _48815_ (_41302_, _40963_, _40861_);
  not _48816_ (_41303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor _48817_ (_41304_, _40861_, _41303_);
  or _48818_ (_43829_, _41304_, _41302_);
  and _48819_ (_41305_, _40966_, _40861_);
  not _48820_ (_41306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor _48821_ (_41307_, _40861_, _41306_);
  or _48822_ (_43833_, _41307_, _41305_);
  and _48823_ (_41308_, _40969_, _40861_);
  not _48824_ (_41309_, _40861_);
  and _48825_ (_41310_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _48826_ (_43837_, _41310_, _41308_);
  and _48827_ (_41311_, _40972_, _40861_);
  and _48828_ (_41312_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or _48829_ (_43841_, _41312_, _41311_);
  and _48830_ (_41313_, _40976_, _40861_);
  and _48831_ (_41314_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _48832_ (_43844_, _41314_, _41313_);
  and _48833_ (_41315_, _40980_, _40861_);
  and _48834_ (_41316_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _48835_ (_43847_, _41316_, _41315_);
  or _48836_ (_41317_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand _48837_ (_41318_, _40417_, _40890_);
  and _48838_ (_41319_, _41318_, _40613_);
  and _48839_ (_41320_, _41319_, _41317_);
  nor _48840_ (_41321_, _40417_, _41010_);
  and _48841_ (_41322_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _48842_ (_41323_, _41322_, _41321_);
  and _48843_ (_41324_, _41323_, _40757_);
  or _48844_ (_41325_, _41324_, _41320_);
  or _48845_ (_41326_, _41325_, _40740_);
  or _48846_ (_41327_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand _48847_ (_41328_, _40417_, _41033_);
  and _48848_ (_41329_, _41328_, _40613_);
  and _48849_ (_41330_, _41329_, _41327_);
  nor _48850_ (_41331_, _40417_, _41098_);
  and _48851_ (_41332_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _48852_ (_41333_, _41332_, _41331_);
  and _48853_ (_41334_, _41333_, _40757_);
  or _48854_ (_41335_, _41334_, _41330_);
  or _48855_ (_41336_, _41335_, _40502_);
  and _48856_ (_41337_, _41336_, _40781_);
  and _48857_ (_41338_, _41337_, _41326_);
  nand _48858_ (_41339_, _40417_, _41121_);
  or _48859_ (_41340_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _48860_ (_41341_, _41340_, _41339_);
  and _48861_ (_41342_, _41341_, _40613_);
  and _48862_ (_41343_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _48863_ (_41344_, _40417_, _41186_);
  or _48864_ (_41345_, _41344_, _41343_);
  and _48865_ (_41346_, _41345_, _40757_);
  or _48866_ (_41347_, _41346_, _41342_);
  or _48867_ (_41348_, _41347_, _40740_);
  nand _48868_ (_41349_, _40417_, _41210_);
  or _48869_ (_41350_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _48870_ (_41351_, _41350_, _41349_);
  and _48871_ (_41352_, _41351_, _40613_);
  and _48872_ (_41353_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _48873_ (_41354_, _40417_, _41300_);
  or _48874_ (_41355_, _41354_, _41353_);
  and _48875_ (_41356_, _41355_, _40757_);
  or _48876_ (_41357_, _41356_, _41352_);
  or _48877_ (_41358_, _41357_, _40502_);
  and _48878_ (_41359_, _41358_, _40708_);
  and _48879_ (_41360_, _41359_, _41348_);
  or _48880_ (_41361_, _41360_, _41338_);
  or _48881_ (_41362_, _41361_, _40734_);
  or _48882_ (_41363_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _48883_ (_41364_, _41363_, _41806_);
  and _48884_ (_01406_, _41364_, _41362_);
  or _48885_ (_41365_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand _48886_ (_41366_, _40417_, _40903_);
  and _48887_ (_41367_, _41366_, _40613_);
  and _48888_ (_41368_, _41367_, _41365_);
  nor _48889_ (_41369_, _40417_, _41013_);
  and _48890_ (_41370_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _48891_ (_41371_, _41370_, _41369_);
  and _48892_ (_41372_, _41371_, _40757_);
  or _48893_ (_41373_, _41372_, _41368_);
  or _48894_ (_41374_, _41373_, _40740_);
  or _48895_ (_41375_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand _48896_ (_41376_, _40417_, _41036_);
  and _48897_ (_41377_, _41376_, _40613_);
  and _48898_ (_41378_, _41377_, _41375_);
  nor _48899_ (_41379_, _40417_, _41101_);
  and _48900_ (_41380_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _48901_ (_41381_, _41380_, _41379_);
  and _48902_ (_41382_, _41381_, _40757_);
  or _48903_ (_41383_, _41382_, _41378_);
  or _48904_ (_41384_, _41383_, _40502_);
  and _48905_ (_41385_, _41384_, _40781_);
  and _48906_ (_41386_, _41385_, _41374_);
  nand _48907_ (_41387_, _40417_, _41124_);
  or _48908_ (_41388_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _48909_ (_41389_, _41388_, _41387_);
  and _48910_ (_41390_, _41389_, _40613_);
  and _48911_ (_41391_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _48912_ (_41392_, _40417_, _41189_);
  or _48913_ (_41393_, _41392_, _41391_);
  and _48914_ (_41394_, _41393_, _40757_);
  or _48915_ (_41395_, _41394_, _41390_);
  or _48916_ (_41396_, _41395_, _40740_);
  nand _48917_ (_41397_, _40417_, _41217_);
  or _48918_ (_41398_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _48919_ (_41399_, _41398_, _41397_);
  and _48920_ (_41400_, _41399_, _40613_);
  and _48921_ (_41401_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _48922_ (_41402_, _40417_, _41303_);
  or _48923_ (_41403_, _41402_, _41401_);
  and _48924_ (_41404_, _41403_, _40757_);
  or _48925_ (_41405_, _41404_, _41400_);
  or _48926_ (_41406_, _41405_, _40502_);
  and _48927_ (_41407_, _41406_, _40708_);
  and _48928_ (_41408_, _41407_, _41396_);
  or _48929_ (_41409_, _41408_, _41386_);
  or _48930_ (_41410_, _41409_, _40734_);
  or _48931_ (_41411_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _48932_ (_41412_, _41411_, _41806_);
  and _48933_ (_01408_, _41412_, _41410_);
  and _48934_ (_41413_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _48935_ (_41414_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _48936_ (_41415_, _41414_, _41413_);
  and _48937_ (_41416_, _41415_, _40613_);
  nor _48938_ (_41417_, _40417_, _41016_);
  and _48939_ (_41418_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _48940_ (_41419_, _41418_, _41417_);
  and _48941_ (_41420_, _41419_, _40757_);
  or _48942_ (_41421_, _41420_, _41416_);
  or _48943_ (_41422_, _41421_, _40740_);
  and _48944_ (_41423_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and _48945_ (_41424_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _48946_ (_41425_, _41424_, _41423_);
  and _48947_ (_41426_, _41425_, _40613_);
  nor _48948_ (_41427_, _40417_, _41104_);
  and _48949_ (_41428_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _48950_ (_41429_, _41428_, _41427_);
  and _48951_ (_41430_, _41429_, _40757_);
  or _48952_ (_41431_, _41430_, _41426_);
  or _48953_ (_41432_, _41431_, _40502_);
  and _48954_ (_41433_, _41432_, _40781_);
  and _48955_ (_41434_, _41433_, _41422_);
  or _48956_ (_41435_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _48957_ (_41436_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _48958_ (_41437_, _41436_, _41435_);
  and _48959_ (_41438_, _41437_, _40613_);
  or _48960_ (_41439_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand _48961_ (_41440_, _40417_, _41168_);
  and _48962_ (_41441_, _41440_, _41439_);
  and _48963_ (_41442_, _41441_, _40757_);
  or _48964_ (_41443_, _41442_, _41438_);
  or _48965_ (_41444_, _41443_, _40740_);
  or _48966_ (_41445_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _48967_ (_41446_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _48968_ (_41447_, _41446_, _41445_);
  and _48969_ (_41448_, _41447_, _40613_);
  or _48970_ (_41449_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand _48971_ (_41450_, _40417_, _41283_);
  and _48972_ (_41451_, _41450_, _41449_);
  and _48973_ (_41452_, _41451_, _40757_);
  or _48974_ (_41453_, _41452_, _41448_);
  or _48975_ (_41454_, _41453_, _40502_);
  and _48976_ (_41455_, _41454_, _40708_);
  and _48977_ (_41456_, _41455_, _41444_);
  or _48978_ (_41457_, _41456_, _41434_);
  or _48979_ (_41458_, _41457_, _40734_);
  or _48980_ (_41459_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _48981_ (_41460_, _41459_, _41806_);
  and _48982_ (_01410_, _41460_, _41458_);
  and _48983_ (_41461_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _48984_ (_41462_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _48985_ (_41463_, _41462_, _41461_);
  and _48986_ (_41464_, _41463_, _40613_);
  nor _48987_ (_41465_, _40417_, _41019_);
  and _48988_ (_41466_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _48989_ (_41467_, _41466_, _41465_);
  and _48990_ (_41468_, _41467_, _40757_);
  or _48991_ (_41469_, _41468_, _41464_);
  or _48992_ (_41470_, _41469_, _40740_);
  or _48993_ (_41471_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand _48994_ (_41472_, _40417_, _41042_);
  and _48995_ (_41473_, _41472_, _40613_);
  and _48996_ (_41474_, _41473_, _41471_);
  nor _48997_ (_41475_, _40417_, _41107_);
  and _48998_ (_41476_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _48999_ (_41477_, _41476_, _41475_);
  and _49000_ (_41478_, _41477_, _40757_);
  or _49001_ (_41479_, _41478_, _41474_);
  or _49002_ (_41480_, _41479_, _40502_);
  and _49003_ (_41481_, _41480_, _40781_);
  and _49004_ (_41482_, _41481_, _41470_);
  nand _49005_ (_41483_, _40417_, _41130_);
  or _49006_ (_41484_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _49007_ (_41485_, _41484_, _41483_);
  and _49008_ (_41486_, _41485_, _40613_);
  or _49009_ (_41487_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand _49010_ (_41488_, _40417_, _41171_);
  and _49011_ (_41489_, _41488_, _41487_);
  and _49012_ (_41490_, _41489_, _40757_);
  or _49013_ (_41491_, _41490_, _41486_);
  or _49014_ (_41492_, _41491_, _40740_);
  nand _49015_ (_41493_, _40417_, _41231_);
  or _49016_ (_41494_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _49017_ (_41495_, _41494_, _41493_);
  and _49018_ (_41496_, _41495_, _40613_);
  or _49019_ (_41497_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand _49020_ (_41498_, _40417_, _41286_);
  and _49021_ (_41499_, _41498_, _41497_);
  and _49022_ (_41500_, _41499_, _40757_);
  or _49023_ (_41501_, _41500_, _41496_);
  or _49024_ (_41502_, _41501_, _40502_);
  and _49025_ (_41503_, _41502_, _40708_);
  and _49026_ (_41504_, _41503_, _41492_);
  or _49027_ (_41505_, _41504_, _41482_);
  or _49028_ (_41506_, _41505_, _40734_);
  or _49029_ (_41507_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _49030_ (_41508_, _41507_, _41806_);
  and _49031_ (_01412_, _41508_, _41506_);
  and _49032_ (_41509_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _49033_ (_41510_, _40417_, _40974_);
  or _49034_ (_41511_, _41510_, _41509_);
  and _49035_ (_41512_, _41511_, _40613_);
  or _49036_ (_41513_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand _49037_ (_41514_, _40417_, _40998_);
  and _49038_ (_41515_, _41514_, _41513_);
  and _49039_ (_41516_, _41515_, _40757_);
  or _49040_ (_41517_, _41516_, _41512_);
  or _49041_ (_41518_, _41517_, _40740_);
  and _49042_ (_41519_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _49043_ (_41520_, _40417_, _41063_);
  or _49044_ (_41521_, _41520_, _41519_);
  and _49045_ (_41522_, _41521_, _40613_);
  or _49046_ (_41523_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand _49047_ (_41524_, _40417_, _41085_);
  and _49048_ (_41525_, _41524_, _41523_);
  and _49049_ (_41526_, _41525_, _40757_);
  or _49050_ (_41527_, _41526_, _41522_);
  or _49051_ (_41528_, _41527_, _40502_);
  and _49052_ (_41529_, _41528_, _40781_);
  and _49053_ (_41530_, _41529_, _41518_);
  and _49054_ (_41531_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _49055_ (_41532_, _40417_, _41152_);
  or _49056_ (_41533_, _41532_, _41531_);
  and _49057_ (_41534_, _41533_, _40613_);
  or _49058_ (_41535_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand _49059_ (_41536_, _40417_, _41174_);
  and _49060_ (_41537_, _41536_, _41535_);
  and _49061_ (_41538_, _41537_, _40757_);
  or _49062_ (_41539_, _41538_, _41534_);
  or _49063_ (_41540_, _41539_, _40740_);
  and _49064_ (_41541_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _49065_ (_41542_, _40417_, _41267_);
  or _49066_ (_41543_, _41542_, _41541_);
  and _49067_ (_41544_, _41543_, _40613_);
  or _49068_ (_41545_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand _49069_ (_41546_, _40417_, _41289_);
  and _49070_ (_41547_, _41546_, _41545_);
  and _49071_ (_41548_, _41547_, _40757_);
  or _49072_ (_41549_, _41548_, _41544_);
  or _49073_ (_41550_, _41549_, _40502_);
  and _49074_ (_41551_, _41550_, _40708_);
  and _49075_ (_41552_, _41551_, _41540_);
  or _49076_ (_41553_, _41552_, _41530_);
  or _49077_ (_41554_, _41553_, _40734_);
  or _49078_ (_41555_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and _49079_ (_41556_, _41555_, _41806_);
  and _49080_ (_01414_, _41556_, _41554_);
  and _49081_ (_41557_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _49082_ (_41558_, _40417_, _40978_);
  or _49083_ (_41559_, _41558_, _41557_);
  and _49084_ (_41560_, _41559_, _40613_);
  or _49085_ (_41561_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand _49086_ (_41562_, _40417_, _41001_);
  and _49087_ (_41563_, _41562_, _41561_);
  and _49088_ (_41564_, _41563_, _40757_);
  or _49089_ (_41565_, _41564_, _41560_);
  or _49090_ (_41566_, _41565_, _40740_);
  and _49091_ (_41567_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _49092_ (_41568_, _40417_, _41066_);
  or _49093_ (_41569_, _41568_, _41567_);
  and _49094_ (_41570_, _41569_, _40613_);
  or _49095_ (_41571_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand _49096_ (_41572_, _40417_, _41088_);
  and _49097_ (_41573_, _41572_, _41571_);
  and _49098_ (_41574_, _41573_, _40757_);
  or _49099_ (_41575_, _41574_, _41570_);
  or _49100_ (_41576_, _41575_, _40502_);
  and _49101_ (_41577_, _41576_, _40781_);
  and _49102_ (_41578_, _41577_, _41566_);
  and _49103_ (_41579_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _49104_ (_41580_, _40417_, _41155_);
  or _49105_ (_41581_, _41580_, _41579_);
  and _49106_ (_41582_, _41581_, _40613_);
  or _49107_ (_41583_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand _49108_ (_41584_, _40417_, _41177_);
  and _49109_ (_41585_, _41584_, _41583_);
  and _49110_ (_41586_, _41585_, _40757_);
  or _49111_ (_41587_, _41586_, _41582_);
  or _49112_ (_41588_, _41587_, _40740_);
  and _49113_ (_41589_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor _49114_ (_41590_, _40417_, _41270_);
  or _49115_ (_41591_, _41590_, _41589_);
  and _49116_ (_41592_, _41591_, _40613_);
  or _49117_ (_41593_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand _49118_ (_41594_, _40417_, _41292_);
  and _49119_ (_41595_, _41594_, _41593_);
  and _49120_ (_41596_, _41595_, _40757_);
  or _49121_ (_41597_, _41596_, _41592_);
  or _49122_ (_41598_, _41597_, _40502_);
  and _49123_ (_41599_, _41598_, _40708_);
  and _49124_ (_41600_, _41599_, _41588_);
  or _49125_ (_41601_, _41600_, _41578_);
  or _49126_ (_41602_, _41601_, _40734_);
  or _49127_ (_41603_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _49128_ (_41604_, _41603_, _41806_);
  and _49129_ (_01416_, _41604_, _41602_);
  and _49130_ (_41605_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and _49131_ (_41606_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _49132_ (_41607_, _41606_, _41605_);
  and _49133_ (_41608_, _41607_, _40613_);
  and _49134_ (_41609_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and _49135_ (_41610_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _49136_ (_41611_, _41610_, _41609_);
  and _49137_ (_41612_, _41611_, _40757_);
  or _49138_ (_41613_, _41612_, _41608_);
  or _49139_ (_41614_, _41613_, _40740_);
  and _49140_ (_41615_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _49141_ (_41616_, _40417_, _41069_);
  or _49142_ (_41617_, _41616_, _41615_);
  and _49143_ (_41618_, _41617_, _40613_);
  or _49144_ (_41619_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nand _49145_ (_41620_, _40417_, _41091_);
  and _49146_ (_41621_, _41620_, _41619_);
  and _49147_ (_41622_, _41621_, _40757_);
  or _49148_ (_41623_, _41622_, _41618_);
  or _49149_ (_41624_, _41623_, _40502_);
  and _49150_ (_41625_, _41624_, _40781_);
  and _49151_ (_41626_, _41625_, _41614_);
  nand _49152_ (_41627_, _40417_, _41137_);
  or _49153_ (_41628_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _49154_ (_41629_, _41628_, _41627_);
  and _49155_ (_41630_, _41629_, _40613_);
  or _49156_ (_41631_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand _49157_ (_41632_, _40417_, _41180_);
  and _49158_ (_41633_, _41632_, _41631_);
  and _49159_ (_41634_, _41633_, _40757_);
  or _49160_ (_41635_, _41634_, _41630_);
  or _49161_ (_41636_, _41635_, _40740_);
  nand _49162_ (_41637_, _40417_, _41248_);
  or _49163_ (_41638_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _49164_ (_41639_, _41638_, _41637_);
  and _49165_ (_41640_, _41639_, _40613_);
  or _49166_ (_41641_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand _49167_ (_41642_, _40417_, _41295_);
  and _49168_ (_41643_, _41642_, _41641_);
  and _49169_ (_41644_, _41643_, _40757_);
  or _49170_ (_41645_, _41644_, _41640_);
  or _49171_ (_41646_, _41645_, _40502_);
  and _49172_ (_41647_, _41646_, _40708_);
  and _49173_ (_41648_, _41647_, _41636_);
  or _49174_ (_41649_, _41648_, _41626_);
  or _49175_ (_41650_, _41649_, _40734_);
  or _49176_ (_41651_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _49177_ (_41652_, _41651_, _41806_);
  and _49178_ (_01418_, _41652_, _41650_);
  or _49179_ (_41653_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not _49180_ (_41654_, \oc8051_gm_cxrom_1.cell0.valid );
  or _49181_ (_41655_, _41654_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand _49182_ (_41656_, _41655_, _41653_);
  nand _49183_ (_41657_, _41656_, _41806_);
  or _49184_ (_41658_, \oc8051_gm_cxrom_1.cell0.data [7], _41806_);
  and _49185_ (_01426_, _41658_, _41657_);
  or _49186_ (_41659_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or _49187_ (_41660_, \oc8051_gm_cxrom_1.cell0.data [0], _41654_);
  nand _49188_ (_41661_, _41660_, _41659_);
  nand _49189_ (_41662_, _41661_, _41806_);
  or _49190_ (_41663_, \oc8051_gm_cxrom_1.cell0.data [0], _41806_);
  and _49191_ (_01433_, _41663_, _41662_);
  or _49192_ (_41664_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or _49193_ (_41665_, \oc8051_gm_cxrom_1.cell0.data [1], _41654_);
  nand _49194_ (_41666_, _41665_, _41664_);
  nand _49195_ (_41667_, _41666_, _41806_);
  or _49196_ (_41668_, \oc8051_gm_cxrom_1.cell0.data [1], _41806_);
  and _49197_ (_01437_, _41668_, _41667_);
  or _49198_ (_41669_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or _49199_ (_41670_, \oc8051_gm_cxrom_1.cell0.data [2], _41654_);
  nand _49200_ (_41671_, _41670_, _41669_);
  nand _49201_ (_41672_, _41671_, _41806_);
  or _49202_ (_41673_, \oc8051_gm_cxrom_1.cell0.data [2], _41806_);
  and _49203_ (_01441_, _41673_, _41672_);
  or _49204_ (_41674_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or _49205_ (_41675_, \oc8051_gm_cxrom_1.cell0.data [3], _41654_);
  nand _49206_ (_41676_, _41675_, _41674_);
  nand _49207_ (_41677_, _41676_, _41806_);
  or _49208_ (_41678_, \oc8051_gm_cxrom_1.cell0.data [3], _41806_);
  and _49209_ (_01444_, _41678_, _41677_);
  or _49210_ (_41679_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or _49211_ (_41680_, \oc8051_gm_cxrom_1.cell0.data [4], _41654_);
  nand _49212_ (_41681_, _41680_, _41679_);
  nand _49213_ (_41682_, _41681_, _41806_);
  or _49214_ (_41683_, \oc8051_gm_cxrom_1.cell0.data [4], _41806_);
  and _49215_ (_01448_, _41683_, _41682_);
  or _49216_ (_41684_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or _49217_ (_41685_, \oc8051_gm_cxrom_1.cell0.data [5], _41654_);
  nand _49218_ (_41686_, _41685_, _41684_);
  nand _49219_ (_41687_, _41686_, _41806_);
  or _49220_ (_41688_, \oc8051_gm_cxrom_1.cell0.data [5], _41806_);
  and _49221_ (_01452_, _41688_, _41687_);
  or _49222_ (_41689_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or _49223_ (_41690_, \oc8051_gm_cxrom_1.cell0.data [6], _41654_);
  nand _49224_ (_41691_, _41690_, _41689_);
  nand _49225_ (_41692_, _41691_, _41806_);
  or _49226_ (_41693_, \oc8051_gm_cxrom_1.cell0.data [6], _41806_);
  and _49227_ (_01456_, _41693_, _41692_);
  or _49228_ (_41694_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not _49229_ (_41695_, \oc8051_gm_cxrom_1.cell1.valid );
  or _49230_ (_41696_, _41695_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand _49231_ (_41697_, _41696_, _41694_);
  nand _49232_ (_41698_, _41697_, _41806_);
  or _49233_ (_41699_, \oc8051_gm_cxrom_1.cell1.data [7], _41806_);
  and _49234_ (_01477_, _41699_, _41698_);
  or _49235_ (_41700_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or _49236_ (_41701_, \oc8051_gm_cxrom_1.cell1.data [0], _41695_);
  nand _49237_ (_41702_, _41701_, _41700_);
  nand _49238_ (_41703_, _41702_, _41806_);
  or _49239_ (_41704_, \oc8051_gm_cxrom_1.cell1.data [0], _41806_);
  and _49240_ (_01484_, _41704_, _41703_);
  or _49241_ (_41705_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or _49242_ (_41706_, \oc8051_gm_cxrom_1.cell1.data [1], _41695_);
  nand _49243_ (_41707_, _41706_, _41705_);
  nand _49244_ (_41708_, _41707_, _41806_);
  or _49245_ (_41709_, \oc8051_gm_cxrom_1.cell1.data [1], _41806_);
  and _49246_ (_01488_, _41709_, _41708_);
  or _49247_ (_41710_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or _49248_ (_41711_, \oc8051_gm_cxrom_1.cell1.data [2], _41695_);
  nand _49249_ (_41712_, _41711_, _41710_);
  nand _49250_ (_41713_, _41712_, _41806_);
  or _49251_ (_41714_, \oc8051_gm_cxrom_1.cell1.data [2], _41806_);
  and _49252_ (_01492_, _41714_, _41713_);
  or _49253_ (_41715_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or _49254_ (_41716_, \oc8051_gm_cxrom_1.cell1.data [3], _41695_);
  nand _49255_ (_41717_, _41716_, _41715_);
  nand _49256_ (_41718_, _41717_, _41806_);
  or _49257_ (_41719_, \oc8051_gm_cxrom_1.cell1.data [3], _41806_);
  and _49258_ (_01496_, _41719_, _41718_);
  or _49259_ (_41720_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or _49260_ (_41721_, \oc8051_gm_cxrom_1.cell1.data [4], _41695_);
  nand _49261_ (_41722_, _41721_, _41720_);
  nand _49262_ (_41723_, _41722_, _41806_);
  or _49263_ (_41724_, \oc8051_gm_cxrom_1.cell1.data [4], _41806_);
  and _49264_ (_01500_, _41724_, _41723_);
  or _49265_ (_41725_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or _49266_ (_41726_, \oc8051_gm_cxrom_1.cell1.data [5], _41695_);
  nand _49267_ (_41727_, _41726_, _41725_);
  nand _49268_ (_41728_, _41727_, _41806_);
  or _49269_ (_41729_, \oc8051_gm_cxrom_1.cell1.data [5], _41806_);
  and _49270_ (_01504_, _41729_, _41728_);
  or _49271_ (_41730_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or _49272_ (_41731_, \oc8051_gm_cxrom_1.cell1.data [6], _41695_);
  nand _49273_ (_41732_, _41731_, _41730_);
  nand _49274_ (_41733_, _41732_, _41806_);
  or _49275_ (_41734_, \oc8051_gm_cxrom_1.cell1.data [6], _41806_);
  and _49276_ (_01508_, _41734_, _41733_);
  or _49277_ (_41735_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not _49278_ (_41736_, \oc8051_gm_cxrom_1.cell2.valid );
  or _49279_ (_41737_, _41736_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand _49280_ (_41738_, _41737_, _41735_);
  nand _49281_ (_41739_, _41738_, _41806_);
  or _49282_ (_41740_, \oc8051_gm_cxrom_1.cell2.data [7], _41806_);
  and _49283_ (_01529_, _41740_, _41739_);
  or _49284_ (_41741_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or _49285_ (_41742_, \oc8051_gm_cxrom_1.cell2.data [0], _41736_);
  nand _49286_ (_41743_, _41742_, _41741_);
  nand _49287_ (_41744_, _41743_, _41806_);
  or _49288_ (_41745_, \oc8051_gm_cxrom_1.cell2.data [0], _41806_);
  and _49289_ (_01536_, _41745_, _41744_);
  or _49290_ (_41746_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or _49291_ (_41747_, \oc8051_gm_cxrom_1.cell2.data [1], _41736_);
  nand _49292_ (_41749_, _41747_, _41746_);
  nand _49293_ (_41750_, _41749_, _41806_);
  or _49294_ (_41752_, \oc8051_gm_cxrom_1.cell2.data [1], _41806_);
  and _49295_ (_01540_, _41752_, _41750_);
  or _49296_ (_41754_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or _49297_ (_41756_, \oc8051_gm_cxrom_1.cell2.data [2], _41736_);
  nand _49298_ (_41758_, _41756_, _41754_);
  nand _49299_ (_41760_, _41758_, _41806_);
  or _49300_ (_41762_, \oc8051_gm_cxrom_1.cell2.data [2], _41806_);
  and _49301_ (_01544_, _41762_, _41760_);
  or _49302_ (_41763_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or _49303_ (_41764_, \oc8051_gm_cxrom_1.cell2.data [3], _41736_);
  nand _49304_ (_41765_, _41764_, _41763_);
  nand _49305_ (_41766_, _41765_, _41806_);
  or _49306_ (_41767_, \oc8051_gm_cxrom_1.cell2.data [3], _41806_);
  and _49307_ (_01548_, _41767_, _41766_);
  or _49308_ (_41768_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or _49309_ (_41769_, \oc8051_gm_cxrom_1.cell2.data [4], _41736_);
  nand _49310_ (_41770_, _41769_, _41768_);
  nand _49311_ (_41771_, _41770_, _41806_);
  or _49312_ (_41772_, \oc8051_gm_cxrom_1.cell2.data [4], _41806_);
  and _49313_ (_01552_, _41772_, _41771_);
  or _49314_ (_41773_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or _49315_ (_41774_, \oc8051_gm_cxrom_1.cell2.data [5], _41736_);
  nand _49316_ (_41775_, _41774_, _41773_);
  nand _49317_ (_41776_, _41775_, _41806_);
  or _49318_ (_41777_, \oc8051_gm_cxrom_1.cell2.data [5], _41806_);
  and _49319_ (_01555_, _41777_, _41776_);
  or _49320_ (_41778_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or _49321_ (_41779_, \oc8051_gm_cxrom_1.cell2.data [6], _41736_);
  nand _49322_ (_41780_, _41779_, _41778_);
  nand _49323_ (_41781_, _41780_, _41806_);
  or _49324_ (_41782_, \oc8051_gm_cxrom_1.cell2.data [6], _41806_);
  and _49325_ (_01559_, _41782_, _41781_);
  or _49326_ (_41783_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not _49327_ (_41784_, \oc8051_gm_cxrom_1.cell3.valid );
  or _49328_ (_41785_, _41784_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand _49329_ (_41786_, _41785_, _41783_);
  nand _49330_ (_41787_, _41786_, _41806_);
  or _49331_ (_41788_, \oc8051_gm_cxrom_1.cell3.data [7], _41806_);
  and _49332_ (_01581_, _41788_, _41787_);
  or _49333_ (_41789_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or _49334_ (_41790_, \oc8051_gm_cxrom_1.cell3.data [0], _41784_);
  nand _49335_ (_41791_, _41790_, _41789_);
  nand _49336_ (_41792_, _41791_, _41806_);
  or _49337_ (_41794_, \oc8051_gm_cxrom_1.cell3.data [0], _41806_);
  and _49338_ (_01588_, _41794_, _41792_);
  or _49339_ (_41797_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or _49340_ (_41799_, \oc8051_gm_cxrom_1.cell3.data [1], _41784_);
  nand _49341_ (_41801_, _41799_, _41797_);
  nand _49342_ (_41803_, _41801_, _41806_);
  or _49343_ (_41805_, \oc8051_gm_cxrom_1.cell3.data [1], _41806_);
  and _49344_ (_01591_, _41805_, _41803_);
  or _49345_ (_41807_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or _49346_ (_41808_, \oc8051_gm_cxrom_1.cell3.data [2], _41784_);
  nand _49347_ (_41809_, _41808_, _41807_);
  nand _49348_ (_41810_, _41809_, _41806_);
  or _49349_ (_41811_, \oc8051_gm_cxrom_1.cell3.data [2], _41806_);
  and _49350_ (_01595_, _41811_, _41810_);
  or _49351_ (_41812_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or _49352_ (_41813_, \oc8051_gm_cxrom_1.cell3.data [3], _41784_);
  nand _49353_ (_41814_, _41813_, _41812_);
  nand _49354_ (_41815_, _41814_, _41806_);
  or _49355_ (_41816_, \oc8051_gm_cxrom_1.cell3.data [3], _41806_);
  and _49356_ (_01599_, _41816_, _41815_);
  or _49357_ (_41817_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or _49358_ (_41818_, \oc8051_gm_cxrom_1.cell3.data [4], _41784_);
  nand _49359_ (_41819_, _41818_, _41817_);
  nand _49360_ (_41820_, _41819_, _41806_);
  or _49361_ (_41821_, \oc8051_gm_cxrom_1.cell3.data [4], _41806_);
  and _49362_ (_01603_, _41821_, _41820_);
  or _49363_ (_41822_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or _49364_ (_41823_, \oc8051_gm_cxrom_1.cell3.data [5], _41784_);
  nand _49365_ (_41824_, _41823_, _41822_);
  nand _49366_ (_41825_, _41824_, _41806_);
  or _49367_ (_41826_, \oc8051_gm_cxrom_1.cell3.data [5], _41806_);
  and _49368_ (_01607_, _41826_, _41825_);
  or _49369_ (_41827_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or _49370_ (_41828_, \oc8051_gm_cxrom_1.cell3.data [6], _41784_);
  nand _49371_ (_41829_, _41828_, _41827_);
  nand _49372_ (_41830_, _41829_, _41806_);
  or _49373_ (_41831_, \oc8051_gm_cxrom_1.cell3.data [6], _41806_);
  and _49374_ (_01611_, _41831_, _41830_);
  or _49375_ (_41832_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not _49376_ (_41833_, \oc8051_gm_cxrom_1.cell4.valid );
  or _49377_ (_41834_, _41833_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand _49378_ (_41835_, _41834_, _41832_);
  nand _49379_ (_41836_, _41835_, _41806_);
  or _49380_ (_41837_, \oc8051_gm_cxrom_1.cell4.data [7], _41806_);
  and _49381_ (_01628_, _41837_, _41836_);
  or _49382_ (_41838_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or _49383_ (_41839_, \oc8051_gm_cxrom_1.cell4.data [0], _41833_);
  nand _49384_ (_41840_, _41839_, _41838_);
  nand _49385_ (_41841_, _41840_, _41806_);
  or _49386_ (_41842_, \oc8051_gm_cxrom_1.cell4.data [0], _41806_);
  and _49387_ (_01630_, _41842_, _41841_);
  or _49388_ (_41843_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or _49389_ (_41844_, \oc8051_gm_cxrom_1.cell4.data [1], _41833_);
  nand _49390_ (_41845_, _41844_, _41843_);
  nand _49391_ (_41846_, _41845_, _41806_);
  or _49392_ (_41847_, \oc8051_gm_cxrom_1.cell4.data [1], _41806_);
  and _49393_ (_01631_, _41847_, _41846_);
  or _49394_ (_41848_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or _49395_ (_41849_, \oc8051_gm_cxrom_1.cell4.data [2], _41833_);
  nand _49396_ (_41850_, _41849_, _41848_);
  nand _49397_ (_41851_, _41850_, _41806_);
  or _49398_ (_41852_, \oc8051_gm_cxrom_1.cell4.data [2], _41806_);
  and _49399_ (_01634_, _41852_, _41851_);
  or _49400_ (_41853_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or _49401_ (_41854_, \oc8051_gm_cxrom_1.cell4.data [3], _41833_);
  nand _49402_ (_41855_, _41854_, _41853_);
  nand _49403_ (_41856_, _41855_, _41806_);
  or _49404_ (_41857_, \oc8051_gm_cxrom_1.cell4.data [3], _41806_);
  and _49405_ (_01638_, _41857_, _41856_);
  or _49406_ (_41858_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or _49407_ (_41859_, \oc8051_gm_cxrom_1.cell4.data [4], _41833_);
  nand _49408_ (_41860_, _41859_, _41858_);
  nand _49409_ (_41861_, _41860_, _41806_);
  or _49410_ (_41862_, \oc8051_gm_cxrom_1.cell4.data [4], _41806_);
  and _49411_ (_01642_, _41862_, _41861_);
  or _49412_ (_41863_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or _49413_ (_41864_, \oc8051_gm_cxrom_1.cell4.data [5], _41833_);
  nand _49414_ (_41865_, _41864_, _41863_);
  nand _49415_ (_41866_, _41865_, _41806_);
  or _49416_ (_41867_, \oc8051_gm_cxrom_1.cell4.data [5], _41806_);
  and _49417_ (_01646_, _41867_, _41866_);
  or _49418_ (_41868_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or _49419_ (_41869_, \oc8051_gm_cxrom_1.cell4.data [6], _41833_);
  nand _49420_ (_41870_, _41869_, _41868_);
  nand _49421_ (_41871_, _41870_, _41806_);
  or _49422_ (_41872_, \oc8051_gm_cxrom_1.cell4.data [6], _41806_);
  and _49423_ (_01650_, _41872_, _41871_);
  or _49424_ (_41873_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not _49425_ (_41874_, \oc8051_gm_cxrom_1.cell5.valid );
  or _49426_ (_41875_, _41874_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand _49427_ (_41876_, _41875_, _41873_);
  nand _49428_ (_41877_, _41876_, _41806_);
  or _49429_ (_41878_, \oc8051_gm_cxrom_1.cell5.data [7], _41806_);
  and _49430_ (_01672_, _41878_, _41877_);
  or _49431_ (_41879_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or _49432_ (_41880_, \oc8051_gm_cxrom_1.cell5.data [0], _41874_);
  nand _49433_ (_41881_, _41880_, _41879_);
  nand _49434_ (_41882_, _41881_, _41806_);
  or _49435_ (_41883_, \oc8051_gm_cxrom_1.cell5.data [0], _41806_);
  and _49436_ (_01679_, _41883_, _41882_);
  or _49437_ (_41884_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or _49438_ (_41885_, \oc8051_gm_cxrom_1.cell5.data [1], _41874_);
  nand _49439_ (_41886_, _41885_, _41884_);
  nand _49440_ (_41887_, _41886_, _41806_);
  or _49441_ (_41888_, \oc8051_gm_cxrom_1.cell5.data [1], _41806_);
  and _49442_ (_01683_, _41888_, _41887_);
  or _49443_ (_41889_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or _49444_ (_41890_, \oc8051_gm_cxrom_1.cell5.data [2], _41874_);
  nand _49445_ (_41891_, _41890_, _41889_);
  nand _49446_ (_41892_, _41891_, _41806_);
  or _49447_ (_41893_, \oc8051_gm_cxrom_1.cell5.data [2], _41806_);
  and _49448_ (_01687_, _41893_, _41892_);
  or _49449_ (_41894_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or _49450_ (_41895_, \oc8051_gm_cxrom_1.cell5.data [3], _41874_);
  nand _49451_ (_41896_, _41895_, _41894_);
  nand _49452_ (_41897_, _41896_, _41806_);
  or _49453_ (_41898_, \oc8051_gm_cxrom_1.cell5.data [3], _41806_);
  and _49454_ (_01691_, _41898_, _41897_);
  or _49455_ (_41899_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or _49456_ (_41900_, \oc8051_gm_cxrom_1.cell5.data [4], _41874_);
  nand _49457_ (_41901_, _41900_, _41899_);
  nand _49458_ (_41902_, _41901_, _41806_);
  or _49459_ (_41903_, \oc8051_gm_cxrom_1.cell5.data [4], _41806_);
  and _49460_ (_01695_, _41903_, _41902_);
  or _49461_ (_41904_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or _49462_ (_41905_, \oc8051_gm_cxrom_1.cell5.data [5], _41874_);
  nand _49463_ (_41906_, _41905_, _41904_);
  nand _49464_ (_41907_, _41906_, _41806_);
  or _49465_ (_41908_, \oc8051_gm_cxrom_1.cell5.data [5], _41806_);
  and _49466_ (_01699_, _41908_, _41907_);
  or _49467_ (_41909_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or _49468_ (_41910_, \oc8051_gm_cxrom_1.cell5.data [6], _41874_);
  nand _49469_ (_41911_, _41910_, _41909_);
  nand _49470_ (_41912_, _41911_, _41806_);
  or _49471_ (_41913_, \oc8051_gm_cxrom_1.cell5.data [6], _41806_);
  and _49472_ (_01703_, _41913_, _41912_);
  or _49473_ (_41914_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not _49474_ (_41915_, \oc8051_gm_cxrom_1.cell6.valid );
  or _49475_ (_41916_, _41915_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand _49476_ (_41917_, _41916_, _41914_);
  nand _49477_ (_41918_, _41917_, _41806_);
  or _49478_ (_41919_, \oc8051_gm_cxrom_1.cell6.data [7], _41806_);
  and _49479_ (_01725_, _41919_, _41918_);
  or _49480_ (_41920_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or _49481_ (_41921_, \oc8051_gm_cxrom_1.cell6.data [0], _41915_);
  nand _49482_ (_41922_, _41921_, _41920_);
  nand _49483_ (_41923_, _41922_, _41806_);
  or _49484_ (_41924_, \oc8051_gm_cxrom_1.cell6.data [0], _41806_);
  and _49485_ (_01732_, _41924_, _41923_);
  or _49486_ (_41925_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or _49487_ (_41926_, \oc8051_gm_cxrom_1.cell6.data [1], _41915_);
  nand _49488_ (_41927_, _41926_, _41925_);
  nand _49489_ (_41928_, _41927_, _41806_);
  or _49490_ (_41929_, \oc8051_gm_cxrom_1.cell6.data [1], _41806_);
  and _49491_ (_01736_, _41929_, _41928_);
  or _49492_ (_41930_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or _49493_ (_41931_, \oc8051_gm_cxrom_1.cell6.data [2], _41915_);
  nand _49494_ (_41932_, _41931_, _41930_);
  nand _49495_ (_41933_, _41932_, _41806_);
  or _49496_ (_41934_, \oc8051_gm_cxrom_1.cell6.data [2], _41806_);
  and _49497_ (_01740_, _41934_, _41933_);
  or _49498_ (_41935_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or _49499_ (_41936_, \oc8051_gm_cxrom_1.cell6.data [3], _41915_);
  nand _49500_ (_41937_, _41936_, _41935_);
  nand _49501_ (_41938_, _41937_, _41806_);
  or _49502_ (_41939_, \oc8051_gm_cxrom_1.cell6.data [3], _41806_);
  and _49503_ (_01743_, _41939_, _41938_);
  or _49504_ (_41940_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or _49505_ (_41941_, \oc8051_gm_cxrom_1.cell6.data [4], _41915_);
  nand _49506_ (_41942_, _41941_, _41940_);
  nand _49507_ (_41943_, _41942_, _41806_);
  or _49508_ (_41944_, \oc8051_gm_cxrom_1.cell6.data [4], _41806_);
  and _49509_ (_01747_, _41944_, _41943_);
  or _49510_ (_41945_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or _49511_ (_41946_, \oc8051_gm_cxrom_1.cell6.data [5], _41915_);
  nand _49512_ (_41947_, _41946_, _41945_);
  nand _49513_ (_41948_, _41947_, _41806_);
  or _49514_ (_41949_, \oc8051_gm_cxrom_1.cell6.data [5], _41806_);
  and _49515_ (_01751_, _41949_, _41948_);
  or _49516_ (_41950_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or _49517_ (_41951_, \oc8051_gm_cxrom_1.cell6.data [6], _41915_);
  nand _49518_ (_41952_, _41951_, _41950_);
  nand _49519_ (_41953_, _41952_, _41806_);
  or _49520_ (_41954_, \oc8051_gm_cxrom_1.cell6.data [6], _41806_);
  and _49521_ (_01755_, _41954_, _41953_);
  or _49522_ (_41955_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not _49523_ (_41956_, \oc8051_gm_cxrom_1.cell7.valid );
  or _49524_ (_41957_, _41956_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand _49525_ (_41958_, _41957_, _41955_);
  nand _49526_ (_41959_, _41958_, _41806_);
  or _49527_ (_41960_, \oc8051_gm_cxrom_1.cell7.data [7], _41806_);
  and _49528_ (_01777_, _41960_, _41959_);
  or _49529_ (_41961_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or _49530_ (_41962_, \oc8051_gm_cxrom_1.cell7.data [0], _41956_);
  nand _49531_ (_41963_, _41962_, _41961_);
  nand _49532_ (_41964_, _41963_, _41806_);
  or _49533_ (_41965_, \oc8051_gm_cxrom_1.cell7.data [0], _41806_);
  and _49534_ (_01783_, _41965_, _41964_);
  or _49535_ (_41966_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or _49536_ (_41967_, \oc8051_gm_cxrom_1.cell7.data [1], _41956_);
  nand _49537_ (_41968_, _41967_, _41966_);
  nand _49538_ (_41969_, _41968_, _41806_);
  or _49539_ (_41970_, \oc8051_gm_cxrom_1.cell7.data [1], _41806_);
  and _49540_ (_01787_, _41970_, _41969_);
  or _49541_ (_41971_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or _49542_ (_41972_, \oc8051_gm_cxrom_1.cell7.data [2], _41956_);
  nand _49543_ (_41973_, _41972_, _41971_);
  nand _49544_ (_41974_, _41973_, _41806_);
  or _49545_ (_41975_, \oc8051_gm_cxrom_1.cell7.data [2], _41806_);
  and _49546_ (_01791_, _41975_, _41974_);
  or _49547_ (_41976_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or _49548_ (_41977_, \oc8051_gm_cxrom_1.cell7.data [3], _41956_);
  nand _49549_ (_41978_, _41977_, _41976_);
  nand _49550_ (_41979_, _41978_, _41806_);
  or _49551_ (_41980_, \oc8051_gm_cxrom_1.cell7.data [3], _41806_);
  and _49552_ (_01795_, _41980_, _41979_);
  or _49553_ (_41981_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or _49554_ (_41982_, \oc8051_gm_cxrom_1.cell7.data [4], _41956_);
  nand _49555_ (_41983_, _41982_, _41981_);
  nand _49556_ (_41984_, _41983_, _41806_);
  or _49557_ (_41985_, \oc8051_gm_cxrom_1.cell7.data [4], _41806_);
  and _49558_ (_01799_, _41985_, _41984_);
  or _49559_ (_41986_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or _49560_ (_41987_, \oc8051_gm_cxrom_1.cell7.data [5], _41956_);
  nand _49561_ (_41988_, _41987_, _41986_);
  nand _49562_ (_41989_, _41988_, _41806_);
  or _49563_ (_41990_, \oc8051_gm_cxrom_1.cell7.data [5], _41806_);
  and _49564_ (_01803_, _41990_, _41989_);
  or _49565_ (_41991_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or _49566_ (_41992_, \oc8051_gm_cxrom_1.cell7.data [6], _41956_);
  nand _49567_ (_41993_, _41992_, _41991_);
  nand _49568_ (_41994_, _41993_, _41806_);
  or _49569_ (_41995_, \oc8051_gm_cxrom_1.cell7.data [6], _41806_);
  and _49570_ (_01807_, _41995_, _41994_);
  or _49571_ (_41996_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not _49572_ (_41997_, \oc8051_gm_cxrom_1.cell8.valid );
  or _49573_ (_41998_, _41997_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand _49574_ (_41999_, _41998_, _41996_);
  nand _49575_ (_42000_, _41999_, _41806_);
  or _49576_ (_42001_, \oc8051_gm_cxrom_1.cell8.data [7], _41806_);
  and _49577_ (_01828_, _42001_, _42000_);
  or _49578_ (_42002_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or _49579_ (_42003_, \oc8051_gm_cxrom_1.cell8.data [0], _41997_);
  nand _49580_ (_42004_, _42003_, _42002_);
  nand _49581_ (_42005_, _42004_, _41806_);
  or _49582_ (_42006_, \oc8051_gm_cxrom_1.cell8.data [0], _41806_);
  and _49583_ (_01835_, _42006_, _42005_);
  or _49584_ (_42007_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or _49585_ (_42008_, \oc8051_gm_cxrom_1.cell8.data [1], _41997_);
  nand _49586_ (_42009_, _42008_, _42007_);
  nand _49587_ (_42010_, _42009_, _41806_);
  or _49588_ (_42011_, \oc8051_gm_cxrom_1.cell8.data [1], _41806_);
  and _49589_ (_01839_, _42011_, _42010_);
  or _49590_ (_42012_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or _49591_ (_42013_, \oc8051_gm_cxrom_1.cell8.data [2], _41997_);
  nand _49592_ (_42014_, _42013_, _42012_);
  nand _49593_ (_42015_, _42014_, _41806_);
  or _49594_ (_42016_, \oc8051_gm_cxrom_1.cell8.data [2], _41806_);
  and _49595_ (_01843_, _42016_, _42015_);
  or _49596_ (_42017_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or _49597_ (_42018_, \oc8051_gm_cxrom_1.cell8.data [3], _41997_);
  nand _49598_ (_42019_, _42018_, _42017_);
  nand _49599_ (_42020_, _42019_, _41806_);
  or _49600_ (_42021_, \oc8051_gm_cxrom_1.cell8.data [3], _41806_);
  and _49601_ (_01847_, _42021_, _42020_);
  or _49602_ (_42022_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or _49603_ (_42023_, \oc8051_gm_cxrom_1.cell8.data [4], _41997_);
  nand _49604_ (_42024_, _42023_, _42022_);
  nand _49605_ (_42025_, _42024_, _41806_);
  or _49606_ (_42026_, \oc8051_gm_cxrom_1.cell8.data [4], _41806_);
  and _49607_ (_01851_, _42026_, _42025_);
  or _49608_ (_42027_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or _49609_ (_42028_, \oc8051_gm_cxrom_1.cell8.data [5], _41997_);
  nand _49610_ (_42029_, _42028_, _42027_);
  nand _49611_ (_42030_, _42029_, _41806_);
  or _49612_ (_42031_, \oc8051_gm_cxrom_1.cell8.data [5], _41806_);
  and _49613_ (_01854_, _42031_, _42030_);
  or _49614_ (_42032_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or _49615_ (_42033_, \oc8051_gm_cxrom_1.cell8.data [6], _41997_);
  nand _49616_ (_42034_, _42033_, _42032_);
  nand _49617_ (_42035_, _42034_, _41806_);
  or _49618_ (_42036_, \oc8051_gm_cxrom_1.cell8.data [6], _41806_);
  and _49619_ (_01858_, _42036_, _42035_);
  or _49620_ (_42037_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not _49621_ (_42038_, \oc8051_gm_cxrom_1.cell9.valid );
  or _49622_ (_42039_, _42038_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand _49623_ (_42040_, _42039_, _42037_);
  nand _49624_ (_42041_, _42040_, _41806_);
  or _49625_ (_42042_, \oc8051_gm_cxrom_1.cell9.data [7], _41806_);
  and _49626_ (_01880_, _42042_, _42041_);
  or _49627_ (_42043_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or _49628_ (_42044_, \oc8051_gm_cxrom_1.cell9.data [0], _42038_);
  nand _49629_ (_42045_, _42044_, _42043_);
  nand _49630_ (_42046_, _42045_, _41806_);
  or _49631_ (_42047_, \oc8051_gm_cxrom_1.cell9.data [0], _41806_);
  and _49632_ (_01887_, _42047_, _42046_);
  or _49633_ (_42048_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or _49634_ (_42049_, \oc8051_gm_cxrom_1.cell9.data [1], _42038_);
  nand _49635_ (_42050_, _42049_, _42048_);
  nand _49636_ (_42051_, _42050_, _41806_);
  or _49637_ (_42052_, \oc8051_gm_cxrom_1.cell9.data [1], _41806_);
  and _49638_ (_01891_, _42052_, _42051_);
  or _49639_ (_42053_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or _49640_ (_42054_, \oc8051_gm_cxrom_1.cell9.data [2], _42038_);
  nand _49641_ (_42055_, _42054_, _42053_);
  nand _49642_ (_42056_, _42055_, _41806_);
  or _49643_ (_42057_, \oc8051_gm_cxrom_1.cell9.data [2], _41806_);
  and _49644_ (_01895_, _42057_, _42056_);
  or _49645_ (_42058_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or _49646_ (_42059_, \oc8051_gm_cxrom_1.cell9.data [3], _42038_);
  nand _49647_ (_42060_, _42059_, _42058_);
  nand _49648_ (_42061_, _42060_, _41806_);
  or _49649_ (_42062_, \oc8051_gm_cxrom_1.cell9.data [3], _41806_);
  and _49650_ (_01899_, _42062_, _42061_);
  or _49651_ (_42063_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or _49652_ (_42064_, \oc8051_gm_cxrom_1.cell9.data [4], _42038_);
  nand _49653_ (_42065_, _42064_, _42063_);
  nand _49654_ (_42066_, _42065_, _41806_);
  or _49655_ (_42067_, \oc8051_gm_cxrom_1.cell9.data [4], _41806_);
  and _49656_ (_01903_, _42067_, _42066_);
  or _49657_ (_42068_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or _49658_ (_42069_, \oc8051_gm_cxrom_1.cell9.data [5], _42038_);
  nand _49659_ (_42070_, _42069_, _42068_);
  nand _49660_ (_42071_, _42070_, _41806_);
  or _49661_ (_42072_, \oc8051_gm_cxrom_1.cell9.data [5], _41806_);
  and _49662_ (_01907_, _42072_, _42071_);
  or _49663_ (_42073_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or _49664_ (_42074_, \oc8051_gm_cxrom_1.cell9.data [6], _42038_);
  nand _49665_ (_42075_, _42074_, _42073_);
  nand _49666_ (_42076_, _42075_, _41806_);
  or _49667_ (_42077_, \oc8051_gm_cxrom_1.cell9.data [6], _41806_);
  and _49668_ (_01910_, _42077_, _42076_);
  or _49669_ (_42078_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not _49670_ (_42079_, \oc8051_gm_cxrom_1.cell10.valid );
  or _49671_ (_42080_, _42079_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand _49672_ (_42081_, _42080_, _42078_);
  nand _49673_ (_42082_, _42081_, _41806_);
  or _49674_ (_42083_, \oc8051_gm_cxrom_1.cell10.data [7], _41806_);
  and _49675_ (_01932_, _42083_, _42082_);
  or _49676_ (_42084_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or _49677_ (_42085_, \oc8051_gm_cxrom_1.cell10.data [0], _42079_);
  nand _49678_ (_42086_, _42085_, _42084_);
  nand _49679_ (_42087_, _42086_, _41806_);
  or _49680_ (_42088_, \oc8051_gm_cxrom_1.cell10.data [0], _41806_);
  and _49681_ (_01939_, _42088_, _42087_);
  or _49682_ (_42089_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or _49683_ (_42090_, \oc8051_gm_cxrom_1.cell10.data [1], _42079_);
  nand _49684_ (_42091_, _42090_, _42089_);
  nand _49685_ (_42092_, _42091_, _41806_);
  or _49686_ (_42093_, \oc8051_gm_cxrom_1.cell10.data [1], _41806_);
  and _49687_ (_01943_, _42093_, _42092_);
  or _49688_ (_42094_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or _49689_ (_42095_, \oc8051_gm_cxrom_1.cell10.data [2], _42079_);
  nand _49690_ (_42096_, _42095_, _42094_);
  nand _49691_ (_42097_, _42096_, _41806_);
  or _49692_ (_42098_, \oc8051_gm_cxrom_1.cell10.data [2], _41806_);
  and _49693_ (_01947_, _42098_, _42097_);
  or _49694_ (_42099_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or _49695_ (_42100_, \oc8051_gm_cxrom_1.cell10.data [3], _42079_);
  nand _49696_ (_42101_, _42100_, _42099_);
  nand _49697_ (_42102_, _42101_, _41806_);
  or _49698_ (_42103_, \oc8051_gm_cxrom_1.cell10.data [3], _41806_);
  and _49699_ (_01951_, _42103_, _42102_);
  or _49700_ (_42104_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or _49701_ (_42105_, \oc8051_gm_cxrom_1.cell10.data [4], _42079_);
  nand _49702_ (_42106_, _42105_, _42104_);
  nand _49703_ (_42107_, _42106_, _41806_);
  or _49704_ (_42108_, \oc8051_gm_cxrom_1.cell10.data [4], _41806_);
  and _49705_ (_01955_, _42108_, _42107_);
  or _49706_ (_42109_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or _49707_ (_42110_, \oc8051_gm_cxrom_1.cell10.data [5], _42079_);
  nand _49708_ (_42111_, _42110_, _42109_);
  nand _49709_ (_42112_, _42111_, _41806_);
  or _49710_ (_42113_, \oc8051_gm_cxrom_1.cell10.data [5], _41806_);
  and _49711_ (_01959_, _42113_, _42112_);
  or _49712_ (_42114_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or _49713_ (_42115_, \oc8051_gm_cxrom_1.cell10.data [6], _42079_);
  nand _49714_ (_42116_, _42115_, _42114_);
  nand _49715_ (_42117_, _42116_, _41806_);
  or _49716_ (_42118_, \oc8051_gm_cxrom_1.cell10.data [6], _41806_);
  and _49717_ (_01963_, _42118_, _42117_);
  or _49718_ (_42119_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not _49719_ (_42120_, \oc8051_gm_cxrom_1.cell11.valid );
  or _49720_ (_42121_, _42120_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand _49721_ (_42122_, _42121_, _42119_);
  nand _49722_ (_42123_, _42122_, _41806_);
  or _49723_ (_42124_, \oc8051_gm_cxrom_1.cell11.data [7], _41806_);
  and _49724_ (_01984_, _42124_, _42123_);
  or _49725_ (_42125_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or _49726_ (_42126_, \oc8051_gm_cxrom_1.cell11.data [0], _42120_);
  nand _49727_ (_42127_, _42126_, _42125_);
  nand _49728_ (_42128_, _42127_, _41806_);
  or _49729_ (_42129_, \oc8051_gm_cxrom_1.cell11.data [0], _41806_);
  and _49730_ (_01991_, _42129_, _42128_);
  or _49731_ (_42130_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or _49732_ (_42131_, \oc8051_gm_cxrom_1.cell11.data [1], _42120_);
  nand _49733_ (_42132_, _42131_, _42130_);
  nand _49734_ (_42133_, _42132_, _41806_);
  or _49735_ (_42134_, \oc8051_gm_cxrom_1.cell11.data [1], _41806_);
  and _49736_ (_01995_, _42134_, _42133_);
  or _49737_ (_42135_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or _49738_ (_42136_, \oc8051_gm_cxrom_1.cell11.data [2], _42120_);
  nand _49739_ (_42137_, _42136_, _42135_);
  nand _49740_ (_42138_, _42137_, _41806_);
  or _49741_ (_42139_, \oc8051_gm_cxrom_1.cell11.data [2], _41806_);
  and _49742_ (_01999_, _42139_, _42138_);
  or _49743_ (_42140_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or _49744_ (_42141_, \oc8051_gm_cxrom_1.cell11.data [3], _42120_);
  nand _49745_ (_42142_, _42141_, _42140_);
  nand _49746_ (_42143_, _42142_, _41806_);
  or _49747_ (_42144_, \oc8051_gm_cxrom_1.cell11.data [3], _41806_);
  and _49748_ (_02003_, _42144_, _42143_);
  or _49749_ (_42145_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or _49750_ (_42146_, \oc8051_gm_cxrom_1.cell11.data [4], _42120_);
  nand _49751_ (_42147_, _42146_, _42145_);
  nand _49752_ (_42148_, _42147_, _41806_);
  or _49753_ (_42149_, \oc8051_gm_cxrom_1.cell11.data [4], _41806_);
  and _49754_ (_02007_, _42149_, _42148_);
  or _49755_ (_42150_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or _49756_ (_42151_, \oc8051_gm_cxrom_1.cell11.data [5], _42120_);
  nand _49757_ (_42152_, _42151_, _42150_);
  nand _49758_ (_42153_, _42152_, _41806_);
  or _49759_ (_42154_, \oc8051_gm_cxrom_1.cell11.data [5], _41806_);
  and _49760_ (_02011_, _42154_, _42153_);
  or _49761_ (_42155_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or _49762_ (_42156_, \oc8051_gm_cxrom_1.cell11.data [6], _42120_);
  nand _49763_ (_42157_, _42156_, _42155_);
  nand _49764_ (_42158_, _42157_, _41806_);
  or _49765_ (_42159_, \oc8051_gm_cxrom_1.cell11.data [6], _41806_);
  and _49766_ (_02015_, _42159_, _42158_);
  or _49767_ (_42160_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not _49768_ (_42161_, \oc8051_gm_cxrom_1.cell12.valid );
  or _49769_ (_42162_, _42161_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand _49770_ (_42163_, _42162_, _42160_);
  nand _49771_ (_42164_, _42163_, _41806_);
  or _49772_ (_42165_, \oc8051_gm_cxrom_1.cell12.data [7], _41806_);
  and _49773_ (_02036_, _42165_, _42164_);
  or _49774_ (_42166_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or _49775_ (_42167_, \oc8051_gm_cxrom_1.cell12.data [0], _42161_);
  nand _49776_ (_42168_, _42167_, _42166_);
  nand _49777_ (_42169_, _42168_, _41806_);
  or _49778_ (_42170_, \oc8051_gm_cxrom_1.cell12.data [0], _41806_);
  and _49779_ (_02043_, _42170_, _42169_);
  or _49780_ (_42171_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or _49781_ (_42172_, \oc8051_gm_cxrom_1.cell12.data [1], _42161_);
  nand _49782_ (_42173_, _42172_, _42171_);
  nand _49783_ (_42174_, _42173_, _41806_);
  or _49784_ (_42175_, \oc8051_gm_cxrom_1.cell12.data [1], _41806_);
  and _49785_ (_02047_, _42175_, _42174_);
  or _49786_ (_42176_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or _49787_ (_42177_, \oc8051_gm_cxrom_1.cell12.data [2], _42161_);
  nand _49788_ (_42178_, _42177_, _42176_);
  nand _49789_ (_42179_, _42178_, _41806_);
  or _49790_ (_42180_, \oc8051_gm_cxrom_1.cell12.data [2], _41806_);
  and _49791_ (_02051_, _42180_, _42179_);
  or _49792_ (_42181_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or _49793_ (_42182_, \oc8051_gm_cxrom_1.cell12.data [3], _42161_);
  nand _49794_ (_42183_, _42182_, _42181_);
  nand _49795_ (_42184_, _42183_, _41806_);
  or _49796_ (_42185_, \oc8051_gm_cxrom_1.cell12.data [3], _41806_);
  and _49797_ (_02055_, _42185_, _42184_);
  or _49798_ (_42186_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or _49799_ (_42187_, \oc8051_gm_cxrom_1.cell12.data [4], _42161_);
  nand _49800_ (_42188_, _42187_, _42186_);
  nand _49801_ (_42189_, _42188_, _41806_);
  or _49802_ (_42190_, \oc8051_gm_cxrom_1.cell12.data [4], _41806_);
  and _49803_ (_02059_, _42190_, _42189_);
  or _49804_ (_42191_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or _49805_ (_42192_, \oc8051_gm_cxrom_1.cell12.data [5], _42161_);
  nand _49806_ (_42193_, _42192_, _42191_);
  nand _49807_ (_42194_, _42193_, _41806_);
  or _49808_ (_42195_, \oc8051_gm_cxrom_1.cell12.data [5], _41806_);
  and _49809_ (_02063_, _42195_, _42194_);
  or _49810_ (_42196_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or _49811_ (_42197_, \oc8051_gm_cxrom_1.cell12.data [6], _42161_);
  nand _49812_ (_42198_, _42197_, _42196_);
  nand _49813_ (_42199_, _42198_, _41806_);
  or _49814_ (_42200_, \oc8051_gm_cxrom_1.cell12.data [6], _41806_);
  and _49815_ (_02067_, _42200_, _42199_);
  or _49816_ (_42201_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not _49817_ (_42202_, \oc8051_gm_cxrom_1.cell13.valid );
  or _49818_ (_42203_, _42202_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand _49819_ (_42204_, _42203_, _42201_);
  nand _49820_ (_42205_, _42204_, _41806_);
  or _49821_ (_42206_, \oc8051_gm_cxrom_1.cell13.data [7], _41806_);
  and _49822_ (_02088_, _42206_, _42205_);
  or _49823_ (_42207_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or _49824_ (_42208_, \oc8051_gm_cxrom_1.cell13.data [0], _42202_);
  nand _49825_ (_42209_, _42208_, _42207_);
  nand _49826_ (_42210_, _42209_, _41806_);
  or _49827_ (_42211_, \oc8051_gm_cxrom_1.cell13.data [0], _41806_);
  and _49828_ (_02095_, _42211_, _42210_);
  or _49829_ (_42212_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or _49830_ (_42213_, \oc8051_gm_cxrom_1.cell13.data [1], _42202_);
  nand _49831_ (_42214_, _42213_, _42212_);
  nand _49832_ (_42215_, _42214_, _41806_);
  or _49833_ (_42216_, \oc8051_gm_cxrom_1.cell13.data [1], _41806_);
  and _49834_ (_02099_, _42216_, _42215_);
  or _49835_ (_42217_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or _49836_ (_42218_, \oc8051_gm_cxrom_1.cell13.data [2], _42202_);
  nand _49837_ (_42219_, _42218_, _42217_);
  nand _49838_ (_42220_, _42219_, _41806_);
  or _49839_ (_42221_, \oc8051_gm_cxrom_1.cell13.data [2], _41806_);
  and _49840_ (_02103_, _42221_, _42220_);
  or _49841_ (_42222_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or _49842_ (_42223_, \oc8051_gm_cxrom_1.cell13.data [3], _42202_);
  nand _49843_ (_42224_, _42223_, _42222_);
  nand _49844_ (_42225_, _42224_, _41806_);
  or _49845_ (_42226_, \oc8051_gm_cxrom_1.cell13.data [3], _41806_);
  and _49846_ (_02107_, _42226_, _42225_);
  or _49847_ (_42227_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or _49848_ (_42228_, \oc8051_gm_cxrom_1.cell13.data [4], _42202_);
  nand _49849_ (_42229_, _42228_, _42227_);
  nand _49850_ (_42230_, _42229_, _41806_);
  or _49851_ (_42231_, \oc8051_gm_cxrom_1.cell13.data [4], _41806_);
  and _49852_ (_02111_, _42231_, _42230_);
  or _49853_ (_42232_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or _49854_ (_42233_, \oc8051_gm_cxrom_1.cell13.data [5], _42202_);
  nand _49855_ (_42234_, _42233_, _42232_);
  nand _49856_ (_42235_, _42234_, _41806_);
  or _49857_ (_42236_, \oc8051_gm_cxrom_1.cell13.data [5], _41806_);
  and _49858_ (_02115_, _42236_, _42235_);
  or _49859_ (_42237_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or _49860_ (_42238_, \oc8051_gm_cxrom_1.cell13.data [6], _42202_);
  nand _49861_ (_42239_, _42238_, _42237_);
  nand _49862_ (_42240_, _42239_, _41806_);
  or _49863_ (_42241_, \oc8051_gm_cxrom_1.cell13.data [6], _41806_);
  and _49864_ (_02119_, _42241_, _42240_);
  or _49865_ (_42242_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not _49866_ (_42243_, \oc8051_gm_cxrom_1.cell14.valid );
  or _49867_ (_42244_, _42243_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand _49868_ (_42245_, _42244_, _42242_);
  nand _49869_ (_42246_, _42245_, _41806_);
  or _49870_ (_42247_, \oc8051_gm_cxrom_1.cell14.data [7], _41806_);
  and _49871_ (_02140_, _42247_, _42246_);
  or _49872_ (_42248_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or _49873_ (_42249_, \oc8051_gm_cxrom_1.cell14.data [0], _42243_);
  nand _49874_ (_42250_, _42249_, _42248_);
  nand _49875_ (_42251_, _42250_, _41806_);
  or _49876_ (_42252_, \oc8051_gm_cxrom_1.cell14.data [0], _41806_);
  and _49877_ (_02147_, _42252_, _42251_);
  or _49878_ (_42253_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or _49879_ (_42254_, \oc8051_gm_cxrom_1.cell14.data [1], _42243_);
  nand _49880_ (_42255_, _42254_, _42253_);
  nand _49881_ (_42256_, _42255_, _41806_);
  or _49882_ (_42257_, \oc8051_gm_cxrom_1.cell14.data [1], _41806_);
  and _49883_ (_02151_, _42257_, _42256_);
  or _49884_ (_42258_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or _49885_ (_42259_, \oc8051_gm_cxrom_1.cell14.data [2], _42243_);
  nand _49886_ (_42260_, _42259_, _42258_);
  nand _49887_ (_42261_, _42260_, _41806_);
  or _49888_ (_42262_, \oc8051_gm_cxrom_1.cell14.data [2], _41806_);
  and _49889_ (_02155_, _42262_, _42261_);
  or _49890_ (_42263_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or _49891_ (_42264_, \oc8051_gm_cxrom_1.cell14.data [3], _42243_);
  nand _49892_ (_42265_, _42264_, _42263_);
  nand _49893_ (_42266_, _42265_, _41806_);
  or _49894_ (_42267_, \oc8051_gm_cxrom_1.cell14.data [3], _41806_);
  and _49895_ (_02159_, _42267_, _42266_);
  or _49896_ (_42268_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or _49897_ (_42269_, \oc8051_gm_cxrom_1.cell14.data [4], _42243_);
  nand _49898_ (_42270_, _42269_, _42268_);
  nand _49899_ (_42271_, _42270_, _41806_);
  or _49900_ (_42272_, \oc8051_gm_cxrom_1.cell14.data [4], _41806_);
  and _49901_ (_02163_, _42272_, _42271_);
  or _49902_ (_42273_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or _49903_ (_42274_, \oc8051_gm_cxrom_1.cell14.data [5], _42243_);
  nand _49904_ (_42275_, _42274_, _42273_);
  nand _49905_ (_42276_, _42275_, _41806_);
  or _49906_ (_42277_, \oc8051_gm_cxrom_1.cell14.data [5], _41806_);
  and _49907_ (_02167_, _42277_, _42276_);
  or _49908_ (_42278_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or _49909_ (_42279_, \oc8051_gm_cxrom_1.cell14.data [6], _42243_);
  nand _49910_ (_42280_, _42279_, _42278_);
  nand _49911_ (_42281_, _42280_, _41806_);
  or _49912_ (_42282_, \oc8051_gm_cxrom_1.cell14.data [6], _41806_);
  and _49913_ (_02171_, _42282_, _42281_);
  or _49914_ (_42283_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not _49915_ (_42284_, \oc8051_gm_cxrom_1.cell15.valid );
  or _49916_ (_42285_, _42284_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand _49917_ (_42286_, _42285_, _42283_);
  nand _49918_ (_42287_, _42286_, _41806_);
  or _49919_ (_42288_, \oc8051_gm_cxrom_1.cell15.data [7], _41806_);
  and _49920_ (_02192_, _42288_, _42287_);
  or _49921_ (_42289_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or _49922_ (_42290_, \oc8051_gm_cxrom_1.cell15.data [0], _42284_);
  nand _49923_ (_42291_, _42290_, _42289_);
  nand _49924_ (_42292_, _42291_, _41806_);
  or _49925_ (_42293_, \oc8051_gm_cxrom_1.cell15.data [0], _41806_);
  and _49926_ (_02199_, _42293_, _42292_);
  or _49927_ (_42294_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or _49928_ (_42295_, \oc8051_gm_cxrom_1.cell15.data [1], _42284_);
  nand _49929_ (_42296_, _42295_, _42294_);
  nand _49930_ (_42297_, _42296_, _41806_);
  or _49931_ (_42298_, \oc8051_gm_cxrom_1.cell15.data [1], _41806_);
  and _49932_ (_02203_, _42298_, _42297_);
  or _49933_ (_42299_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or _49934_ (_42300_, \oc8051_gm_cxrom_1.cell15.data [2], _42284_);
  nand _49935_ (_42301_, _42300_, _42299_);
  nand _49936_ (_42302_, _42301_, _41806_);
  or _49937_ (_42303_, \oc8051_gm_cxrom_1.cell15.data [2], _41806_);
  and _49938_ (_02207_, _42303_, _42302_);
  or _49939_ (_42304_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or _49940_ (_42305_, \oc8051_gm_cxrom_1.cell15.data [3], _42284_);
  nand _49941_ (_42306_, _42305_, _42304_);
  nand _49942_ (_42307_, _42306_, _41806_);
  or _49943_ (_42308_, \oc8051_gm_cxrom_1.cell15.data [3], _41806_);
  and _49944_ (_02211_, _42308_, _42307_);
  or _49945_ (_42309_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or _49946_ (_42310_, \oc8051_gm_cxrom_1.cell15.data [4], _42284_);
  nand _49947_ (_42311_, _42310_, _42309_);
  nand _49948_ (_42312_, _42311_, _41806_);
  or _49949_ (_42313_, \oc8051_gm_cxrom_1.cell15.data [4], _41806_);
  and _49950_ (_02215_, _42313_, _42312_);
  or _49951_ (_42314_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or _49952_ (_42315_, \oc8051_gm_cxrom_1.cell15.data [5], _42284_);
  nand _49953_ (_42316_, _42315_, _42314_);
  nand _49954_ (_42317_, _42316_, _41806_);
  or _49955_ (_42318_, \oc8051_gm_cxrom_1.cell15.data [5], _41806_);
  and _49956_ (_02219_, _42318_, _42317_);
  or _49957_ (_42319_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or _49958_ (_42320_, \oc8051_gm_cxrom_1.cell15.data [6], _42284_);
  nand _49959_ (_42321_, _42320_, _42319_);
  nand _49960_ (_42322_, _42321_, _41806_);
  or _49961_ (_42323_, \oc8051_gm_cxrom_1.cell15.data [6], _41806_);
  and _49962_ (_02223_, _42323_, _42322_);
  nor _49963_ (_05996_, _37932_, rst);
  and _49964_ (_42324_, _33860_, _41806_);
  nand _49965_ (_42325_, _42324_, _36091_);
  nor _49966_ (_42326_, _36584_, _36453_);
  or _49967_ (_05999_, _42326_, _42325_);
  and _49968_ (_42327_, _35242_, _35012_);
  and _49969_ (_42328_, _42327_, _35496_);
  not _49970_ (_42329_, _34486_);
  nor _49971_ (_42330_, _34727_, _34233_);
  and _49972_ (_42331_, _42330_, _42329_);
  and _49973_ (_42332_, _42331_, _42328_);
  not _49974_ (_42333_, _34233_);
  and _49975_ (_42334_, _34727_, _42333_);
  not _49976_ (_42335_, _35751_);
  not _49977_ (_42336_, _35242_);
  and _49978_ (_42337_, _35496_, _42336_);
  not _49979_ (_42338_, _35012_);
  and _49980_ (_42339_, _36365_, _42338_);
  and _49981_ (_42340_, _42339_, _42337_);
  and _49982_ (_42341_, _42340_, _42335_);
  and _49983_ (_42342_, _42341_, _42334_);
  and _49984_ (_42343_, _42335_, _34486_);
  nor _49985_ (_42344_, _42335_, _34486_);
  nor _49986_ (_42345_, _42344_, _42343_);
  and _49987_ (_42346_, _35496_, _35242_);
  and _49988_ (_42347_, _42346_, _42339_);
  and _49989_ (_42348_, _34727_, _34233_);
  and _49990_ (_42349_, _42348_, _42347_);
  and _49991_ (_42350_, _42349_, _42345_);
  or _49992_ (_42351_, _42350_, _42342_);
  or _49993_ (_42352_, _42351_, _42332_);
  not _49994_ (_42353_, _34727_);
  and _49995_ (_42354_, _42353_, _34233_);
  and _49996_ (_42355_, _42354_, _42344_);
  not _49997_ (_42356_, _36365_);
  and _49998_ (_42357_, _42328_, _42356_);
  and _49999_ (_42358_, _42357_, _42355_);
  and _50000_ (_42359_, _42344_, _42334_);
  not _50001_ (_42360_, _35496_);
  and _50002_ (_42361_, _42336_, _35012_);
  nor _50003_ (_42362_, _42361_, _42360_);
  not _50004_ (_42363_, _42362_);
  and _50005_ (_42364_, _42363_, _42359_);
  or _50006_ (_42365_, _42364_, _42358_);
  and _50007_ (_42366_, _35751_, _34486_);
  and _50008_ (_42367_, _42366_, _42330_);
  and _50009_ (_42368_, _42337_, _42338_);
  and _50010_ (_42369_, _42368_, _42356_);
  and _50011_ (_42370_, _42369_, _42367_);
  and _50012_ (_42371_, _42348_, _42329_);
  and _50013_ (_42372_, _42328_, _36365_);
  and _50014_ (_42373_, _42372_, _42371_);
  or _50015_ (_42374_, _42373_, _42370_);
  or _50016_ (_42375_, _42374_, _42365_);
  and _50017_ (_42376_, _42343_, _42334_);
  and _50018_ (_42377_, _42347_, _42376_);
  and _50019_ (_42378_, _42367_, _42360_);
  nor _50020_ (_42379_, _42378_, _42377_);
  and _50021_ (_42380_, _42354_, _35751_);
  and _50022_ (_42381_, _42380_, _42347_);
  and _50023_ (_42382_, _42348_, _34486_);
  and _50024_ (_42383_, _42382_, _42372_);
  nor _50025_ (_42384_, _42383_, _42381_);
  nand _50026_ (_42385_, _42384_, _42379_);
  or _50027_ (_42386_, _42385_, _42375_);
  nor _50028_ (_42387_, _35751_, _34486_);
  and _50029_ (_42388_, _42354_, _42387_);
  nor _50030_ (_42389_, _42388_, _42356_);
  and _50031_ (_42390_, _42346_, _42338_);
  not _50032_ (_42391_, _42390_);
  nor _50033_ (_42392_, _42391_, _42389_);
  not _50034_ (_42393_, _42392_);
  and _50035_ (_42394_, _42348_, _42344_);
  and _50036_ (_42395_, _42394_, _42347_);
  and _50037_ (_42396_, _42354_, _42343_);
  and _50038_ (_42397_, _42396_, _42347_);
  nor _50039_ (_42398_, _42397_, _42395_);
  and _50040_ (_42399_, _42398_, _42393_);
  and _50041_ (_42400_, _42359_, _42368_);
  and _50042_ (_42401_, _42334_, _34486_);
  and _50043_ (_42402_, _42357_, _42401_);
  and _50044_ (_42403_, _42347_, _42331_);
  or _50045_ (_42404_, _42403_, _42402_);
  nor _50046_ (_42405_, _42404_, _42400_);
  nand _50047_ (_42406_, _42405_, _42399_);
  or _50048_ (_42407_, _42406_, _42386_);
  or _50049_ (_42408_, _42407_, _42352_);
  and _50050_ (_42409_, _42408_, _33881_);
  not _50051_ (_42410_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _50052_ (_42411_, _33849_, _15636_);
  and _50053_ (_42412_, _42411_, _36727_);
  nor _50054_ (_42413_, _42412_, _42410_);
  or _50055_ (_42414_, _42413_, rst);
  or _50056_ (_06002_, _42414_, _42409_);
  nand _50057_ (_42415_, _34233_, _33806_);
  or _50058_ (_42416_, _33806_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _50059_ (_42417_, _42416_, _41806_);
  and _50060_ (_06005_, _42417_, _42415_);
  and _50061_ (_42418_, \oc8051_top_1.oc8051_sfr1.wait_data , _41806_);
  and _50062_ (_42419_, _42418_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _50063_ (_42420_, _36464_, _36124_);
  and _50064_ (_42421_, _37833_, _36935_);
  or _50065_ (_42422_, _42421_, _42420_);
  and _50066_ (_42423_, _36584_, _36124_);
  or _50067_ (_42424_, _42423_, _37657_);
  or _50068_ (_42425_, _42424_, _37340_);
  and _50069_ (_42426_, _37102_, _36464_);
  and _50070_ (_42427_, _36595_, _36453_);
  or _50071_ (_42428_, _42427_, _42426_);
  or _50072_ (_42429_, _42428_, _42425_);
  or _50073_ (_42430_, _42429_, _37550_);
  or _50074_ (_42431_, _42430_, _42422_);
  and _50075_ (_42432_, _42431_, _42324_);
  or _50076_ (_06008_, _42432_, _42419_);
  and _50077_ (_42433_, _36584_, _36003_);
  or _50078_ (_42434_, _42433_, _36485_);
  and _50079_ (_42435_, _37023_, _36025_);
  or _50080_ (_42436_, _42435_, _36036_);
  and _50081_ (_42437_, _36880_, _35056_);
  and _50082_ (_42438_, _42437_, _37102_);
  or _50083_ (_42439_, _42438_, _42436_);
  or _50084_ (_42440_, _42439_, _42434_);
  and _50085_ (_42441_, _42440_, _33860_);
  and _50086_ (_42442_, \oc8051_top_1.oc8051_decoder1.state [0], _15636_);
  and _50087_ (_42443_, _42442_, _42410_);
  not _50088_ (_42444_, _37866_);
  and _50089_ (_42445_, _42444_, _42443_);
  and _50090_ (_42446_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50091_ (_42447_, _42446_, _42445_);
  or _50092_ (_42448_, _42447_, _42441_);
  and _50093_ (_06011_, _42448_, _41806_);
  and _50094_ (_42449_, _42418_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _50095_ (_42450_, _37833_, _37045_);
  not _50096_ (_42451_, _36902_);
  nor _50097_ (_42452_, _37045_, _36595_);
  nor _50098_ (_42453_, _42452_, _42451_);
  or _50099_ (_42454_, _42453_, _42450_);
  and _50100_ (_42455_, _42437_, _37186_);
  or _50101_ (_42456_, _42455_, _42454_);
  nor _50102_ (_42457_, _42452_, _35542_);
  not _50103_ (_42458_, _35542_);
  and _50104_ (_42459_, _37186_, _42458_);
  or _50105_ (_42460_, _42459_, _42457_);
  nor _50106_ (_42461_, _35795_, _35542_);
  and _50107_ (_42462_, _42461_, _35959_);
  and _50108_ (_42463_, _37833_, _36913_);
  nor _50109_ (_42464_, _42463_, _42462_);
  nand _50110_ (_42465_, _42464_, _35981_);
  or _50111_ (_42466_, _42465_, _42434_);
  or _50112_ (_42467_, _42466_, _42460_);
  or _50113_ (_42468_, _42467_, _42456_);
  and _50114_ (_42469_, _42468_, _42324_);
  or _50115_ (_06014_, _42469_, _42449_);
  and _50116_ (_42470_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _50117_ (_42471_, _37394_, _33860_);
  or _50118_ (_42472_, _42471_, _42470_);
  or _50119_ (_42473_, _42472_, _42445_);
  and _50120_ (_06017_, _42473_, _41806_);
  and _50121_ (_42474_, _36464_, _35992_);
  not _50122_ (_42475_, _36935_);
  nor _50123_ (_42476_, _42326_, _42475_);
  nor _50124_ (_42477_, _42476_, _42474_);
  not _50125_ (_42478_, _42477_);
  and _50126_ (_42479_, _42478_, _42443_);
  and _50127_ (_42480_, _37186_, _36628_);
  and _50128_ (_42481_, _36891_, _36442_);
  and _50129_ (_42482_, _42481_, _35806_);
  or _50130_ (_42483_, _42482_, _42480_);
  or _50131_ (_42484_, _42483_, _42420_);
  and _50132_ (_42485_, _42484_, _36858_);
  or _50133_ (_42486_, _42485_, _42479_);
  and _50134_ (_42487_, _42483_, _36749_);
  or _50135_ (_42488_, _42487_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50136_ (_42489_, _42488_, _42486_);
  or _50137_ (_42490_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _15636_);
  and _50138_ (_42491_, _42490_, _41806_);
  and _50139_ (_06020_, _42491_, _42489_);
  and _50140_ (_42492_, _42418_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _50141_ (_42493_, _42459_, _36485_);
  and _50142_ (_42494_, _36595_, _42458_);
  or _50143_ (_42495_, _42494_, _37263_);
  or _50144_ (_42496_, _42495_, _42493_);
  and _50145_ (_42497_, _36628_, _35959_);
  or _50146_ (_42498_, _42455_, _42427_);
  or _50147_ (_42499_, _42498_, _42497_);
  or _50148_ (_42500_, _37186_, _37102_);
  and _50149_ (_42501_, _42500_, _35850_);
  or _50150_ (_42502_, _42435_, _37110_);
  or _50151_ (_42503_, _42502_, _42501_);
  or _50152_ (_42504_, _42503_, _42499_);
  or _50153_ (_42505_, _42504_, _42496_);
  and _50154_ (_42506_, _42505_, _42324_);
  or _50155_ (_06023_, _42506_, _42492_);
  and _50156_ (_42507_, _42418_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or _50157_ (_42508_, _42438_, _37219_);
  and _50158_ (_42509_, _36464_, _35860_);
  and _50159_ (_42510_, _42437_, _36650_);
  or _50160_ (_42511_, _42510_, _42509_);
  or _50161_ (_42512_, _42511_, _42508_);
  or _50162_ (_42513_, _42512_, _42460_);
  and _50163_ (_42514_, _37833_, _37164_);
  or _50164_ (_42515_, _37252_, _37175_);
  or _50165_ (_42516_, _42515_, _42514_);
  and _50166_ (_42517_, _36069_, _34782_);
  or _50167_ (_42518_, _42517_, _36661_);
  and _50168_ (_42519_, _36595_, _35850_);
  or _50169_ (_42520_, _42519_, _42518_);
  or _50170_ (_42521_, _42520_, _42516_);
  or _50171_ (_42522_, _42521_, _42513_);
  and _50172_ (_42523_, _37023_, _34782_);
  and _50173_ (_42524_, _37023_, _36507_);
  or _50174_ (_42525_, _42524_, _42523_);
  nor _50175_ (_42526_, _37421_, _35926_);
  nand _50176_ (_42527_, _42526_, _37318_);
  or _50177_ (_42528_, _42527_, _42525_);
  or _50178_ (_42529_, _42528_, _42456_);
  or _50179_ (_42530_, _42529_, _42522_);
  and _50180_ (_42531_, _42530_, _42324_);
  or _50181_ (_06026_, _42531_, _42507_);
  and _50182_ (_42532_, _42461_, _35992_);
  or _50183_ (_42533_, _42532_, _35882_);
  and _50184_ (_42534_, _42437_, _35871_);
  and _50185_ (_42535_, _35871_, _42458_);
  or _50186_ (_42536_, _42535_, _36014_);
  or _50187_ (_42537_, _42536_, _42534_);
  or _50188_ (_42538_, _42537_, _42533_);
  and _50189_ (_42539_, _42437_, _36003_);
  or _50190_ (_42540_, _42539_, _42538_);
  and _50191_ (_42541_, _42540_, _33860_);
  and _50192_ (_42542_, _37855_, _15636_);
  and _50193_ (_42543_, _37844_, _15636_);
  or _50194_ (_42544_, _42543_, _42542_);
  and _50195_ (_42545_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _50196_ (_42546_, _42545_, _42544_);
  or _50197_ (_42547_, _42546_, _42541_);
  and _50198_ (_06029_, _42547_, _41806_);
  or _50199_ (_42548_, _37133_, _37110_);
  not _50200_ (_42549_, _37351_);
  or _50201_ (_42550_, _42453_, _42549_);
  or _50202_ (_42551_, _42550_, _42548_);
  and _50203_ (_42552_, _36080_, _35806_);
  and _50204_ (_42553_, _42552_, _36902_);
  or _50205_ (_42554_, _42553_, _37197_);
  or _50206_ (_42555_, _42554_, _37175_);
  or _50207_ (_42556_, _42555_, _42480_);
  or _50208_ (_42557_, _42556_, _37443_);
  or _50209_ (_42558_, _42557_, _42551_);
  or _50210_ (_42559_, _37034_, _36135_);
  or _50211_ (_42560_, _42559_, _37464_);
  or _50212_ (_42561_, _42560_, _42436_);
  and _50213_ (_42562_, _42552_, _35850_);
  or _50214_ (_42563_, _42562_, _35926_);
  or _50215_ (_42564_, _42563_, _36957_);
  and _50216_ (_42565_, _36124_, _42458_);
  and _50217_ (_42566_, _42461_, _36080_);
  or _50218_ (_42567_, _42566_, _42482_);
  or _50219_ (_42568_, _42567_, _42565_);
  or _50220_ (_42569_, _42568_, _42564_);
  or _50221_ (_42570_, _42569_, _42561_);
  or _50222_ (_42571_, _42570_, _42460_);
  or _50223_ (_42572_, _42571_, _42558_);
  and _50224_ (_42573_, _42572_, _33860_);
  and _50225_ (_42574_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50226_ (_42575_, _42487_, _42445_);
  and _50227_ (_42576_, _37712_, _36749_);
  or _50228_ (_42577_, _42576_, _42575_);
  or _50229_ (_42578_, _42577_, _42574_);
  or _50230_ (_42579_, _42578_, _42573_);
  and _50231_ (_06032_, _42579_, _41806_);
  nor _50232_ (_06091_, _36814_, rst);
  nor _50233_ (_06093_, _37778_, rst);
  nand _50234_ (_06096_, _42478_, _42324_);
  and _50235_ (_42580_, _36584_, _36091_);
  or _50236_ (_42581_, _42580_, _42474_);
  nand _50237_ (_06099_, _42581_, _42324_);
  or _50238_ (_42582_, _42373_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _50239_ (_42583_, _42582_, _42402_);
  or _50240_ (_42584_, _42583_, _42342_);
  and _50241_ (_42585_, _42584_, _42412_);
  nor _50242_ (_42586_, _42411_, _36727_);
  or _50243_ (_42587_, _42586_, rst);
  or _50244_ (_06102_, _42587_, _42585_);
  nand _50245_ (_42588_, _36365_, _33806_);
  or _50246_ (_42589_, _33806_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _50247_ (_42590_, _42589_, _41806_);
  and _50248_ (_06105_, _42590_, _42588_);
  not _50249_ (_42591_, _33806_);
  or _50250_ (_42592_, _35012_, _42591_);
  or _50251_ (_42593_, _33806_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _50252_ (_42594_, _42593_, _41806_);
  and _50253_ (_06108_, _42594_, _42592_);
  nand _50254_ (_42595_, _35242_, _33806_);
  or _50255_ (_42596_, _33806_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _50256_ (_42597_, _42596_, _41806_);
  and _50257_ (_06111_, _42597_, _42595_);
  nand _50258_ (_42598_, _35496_, _33806_);
  or _50259_ (_42599_, _33806_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _50260_ (_42600_, _42599_, _41806_);
  and _50261_ (_06114_, _42600_, _42598_);
  or _50262_ (_42601_, _35751_, _42591_);
  or _50263_ (_42602_, _33806_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _50264_ (_42603_, _42602_, _41806_);
  and _50265_ (_06117_, _42603_, _42601_);
  nand _50266_ (_42604_, _34486_, _33806_);
  or _50267_ (_42605_, _33806_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _50268_ (_42606_, _42605_, _41806_);
  and _50269_ (_06120_, _42606_, _42604_);
  nand _50270_ (_42607_, _34727_, _33806_);
  or _50271_ (_42608_, _33806_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _50272_ (_42609_, _42608_, _41806_);
  and _50273_ (_06123_, _42609_, _42607_);
  and _50274_ (_42610_, _37023_, _34793_);
  or _50275_ (_42611_, _42534_, _36014_);
  or _50276_ (_42612_, _42611_, _42610_);
  or _50277_ (_42613_, _36485_, _36113_);
  or _50278_ (_42614_, _42613_, _42612_);
  and _50279_ (_42615_, _42437_, _37164_);
  or _50280_ (_42616_, _42615_, _42433_);
  or _50281_ (_42617_, _36595_, _35915_);
  and _50282_ (_42618_, _42617_, _37833_);
  or _50283_ (_42619_, _42618_, _42616_);
  or _50284_ (_42620_, _42619_, _42614_);
  or _50285_ (_42621_, _42524_, _42509_);
  and _50286_ (_42622_, _42437_, _36990_);
  or _50287_ (_42623_, _42622_, _42533_);
  or _50288_ (_42624_, _42623_, _42621_);
  or _50289_ (_42625_, _36946_, _36661_);
  or _50290_ (_42626_, _42510_, _42421_);
  or _50291_ (_42627_, _42626_, _42625_);
  or _50292_ (_42628_, _42627_, _42624_);
  and _50293_ (_42629_, _37001_, _42458_);
  or _50294_ (_42630_, _42629_, _42539_);
  and _50295_ (_42631_, _36091_, _35806_);
  and _50296_ (_42632_, _42631_, _37833_);
  or _50297_ (_42633_, _42632_, _35839_);
  and _50298_ (_42634_, _37833_, _36518_);
  and _50299_ (_42635_, _37023_, _36091_);
  or _50300_ (_42636_, _42635_, _42634_);
  or _50301_ (_42637_, _42636_, _42633_);
  or _50302_ (_42638_, _42637_, _42630_);
  or _50303_ (_42639_, _42638_, _42628_);
  or _50304_ (_42640_, _42639_, _42620_);
  and _50305_ (_42641_, _42640_, _33860_);
  and _50306_ (_42642_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50307_ (_42643_, _42642_, _42479_);
  or _50308_ (_42644_, _42643_, _42641_);
  and _50309_ (_30468_, _42644_, _41806_);
  and _50310_ (_42645_, _42418_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _50311_ (_42646_, _37164_, _36650_);
  and _50312_ (_42647_, _42646_, _36628_);
  or _50313_ (_42648_, _42616_, _42525_);
  or _50314_ (_42649_, _42648_, _42647_);
  nor _50315_ (_42650_, _42462_, _35970_);
  not _50316_ (_42651_, _42650_);
  or _50317_ (_42652_, _42651_, _42463_);
  or _50318_ (_42653_, _42652_, _37118_);
  or _50319_ (_42654_, _42653_, _42422_);
  or _50320_ (_42655_, _36650_, _37001_);
  and _50321_ (_42656_, _42655_, _37833_);
  or _50322_ (_42657_, _42656_, _42520_);
  or _50323_ (_42658_, _42657_, _42654_);
  or _50324_ (_42659_, _42658_, _42649_);
  and _50325_ (_42660_, _42659_, _42324_);
  or _50326_ (_30471_, _42660_, _42645_);
  or _50327_ (_42661_, _42482_, _36135_);
  or _50328_ (_42662_, _42661_, _42565_);
  or _50329_ (_42663_, _42662_, _37464_);
  or _50330_ (_42664_, _42663_, _42558_);
  and _50331_ (_42665_, _42664_, _33860_);
  and _50332_ (_42666_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50333_ (_42667_, _42666_, _42577_);
  or _50334_ (_42668_, _42667_, _42665_);
  and _50335_ (_30473_, _42668_, _41806_);
  and _50336_ (_42669_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _50337_ (_42670_, _37416_, _35795_);
  or _50338_ (_42671_, _42670_, _36036_);
  or _50339_ (_42672_, _42671_, _42564_);
  or _50340_ (_42673_, _42672_, _42483_);
  and _50341_ (_42674_, _42673_, _33860_);
  or _50342_ (_42675_, _42674_, _42669_);
  or _50343_ (_42676_, _42675_, _42575_);
  and _50344_ (_30475_, _42676_, _41806_);
  and _50345_ (_42677_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50346_ (_42678_, _42479_, _37910_);
  or _50347_ (_42679_, _42678_, _42677_);
  and _50348_ (_42680_, _42679_, _41806_);
  or _50349_ (_42681_, _42474_, _37855_);
  and _50350_ (_42682_, _42534_, _35806_);
  or _50351_ (_42683_, _42682_, _42622_);
  or _50352_ (_42684_, _42683_, _42681_);
  or _50353_ (_42685_, _42684_, _42483_);
  or _50354_ (_42686_, _42533_, _35839_);
  or _50355_ (_42687_, _42646_, _36518_);
  and _50356_ (_42688_, _42687_, _37833_);
  or _50357_ (_42689_, _42688_, _42686_);
  or _50358_ (_42690_, _42689_, _42685_);
  and _50359_ (_42691_, _37833_, _37102_);
  or _50360_ (_42692_, _42509_, _42691_);
  or _50361_ (_42693_, _42692_, _42630_);
  and _50362_ (_42694_, _42437_, _37208_);
  or _50363_ (_42695_, _42694_, _42421_);
  or _50364_ (_42696_, _42632_, _37844_);
  or _50365_ (_42697_, _42696_, _42618_);
  or _50366_ (_42698_, _42697_, _42695_);
  and _50367_ (_42699_, _42631_, _36902_);
  or _50368_ (_42700_, _42562_, _36014_);
  or _50369_ (_42701_, _42700_, _42566_);
  or _50370_ (_42702_, _42701_, _42699_);
  and _50371_ (_42703_, _42534_, _35795_);
  or _50372_ (_42704_, _42703_, _36529_);
  and _50373_ (_42705_, _37464_, _36409_);
  or _50374_ (_42706_, _42705_, _42704_);
  or _50375_ (_42707_, _42706_, _42702_);
  or _50376_ (_42708_, _42707_, _42698_);
  or _50377_ (_42709_, _42708_, _42693_);
  or _50378_ (_42710_, _42709_, _42690_);
  and _50379_ (_42711_, _42710_, _42324_);
  or _50380_ (_30477_, _42711_, _42680_);
  or _50381_ (_42712_, _37855_, _36014_);
  or _50382_ (_42713_, _42553_, _42433_);
  or _50383_ (_42714_, _42713_, _42712_);
  or _50384_ (_42715_, _35297_, _42458_);
  and _50385_ (_42716_, _42715_, _42631_);
  or _50386_ (_42717_, _42716_, _37464_);
  or _50387_ (_42718_, _42717_, _42714_);
  or _50388_ (_42719_, _37012_, _36551_);
  or _50389_ (_42720_, _42719_, _42718_);
  or _50390_ (_42721_, _37421_, _37175_);
  and _50391_ (_42722_, _42721_, _36420_);
  or _50392_ (_42723_, _42722_, _42686_);
  or _50393_ (_42724_, _42723_, _42720_);
  or _50394_ (_42725_, _42698_, _42693_);
  or _50395_ (_42726_, _42725_, _42724_);
  and _50396_ (_42727_, _42726_, _33860_);
  and _50397_ (_42728_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50398_ (_42730_, _42728_, _42678_);
  or _50399_ (_42732_, _42730_, _42727_);
  and _50400_ (_30479_, _42732_, _41806_);
  and _50401_ (_42735_, _42418_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not _50402_ (_42737_, _40330_);
  or _50403_ (_42739_, _42539_, _42737_);
  and _50404_ (_42741_, _36464_, _35915_);
  and _50405_ (_42743_, _42741_, _35806_);
  and _50406_ (_42745_, _42427_, _36420_);
  or _50407_ (_42747_, _42745_, _42743_);
  or _50408_ (_42749_, _42747_, _42496_);
  or _50409_ (_42751_, _42749_, _42739_);
  not _50410_ (_42753_, _40329_);
  or _50411_ (_42755_, _42501_, _42753_);
  and _50412_ (_42757_, _37833_, _36595_);
  or _50413_ (_42759_, _42757_, _42455_);
  or _50414_ (_42761_, _42759_, _42548_);
  or _50415_ (_42763_, _42761_, _42755_);
  and _50416_ (_42765_, _36464_, _37208_);
  or _50417_ (_42767_, _42532_, _42435_);
  and _50418_ (_42769_, _35882_, _35806_);
  or _50419_ (_42771_, _42769_, _42767_);
  or _50420_ (_42773_, _42771_, _42765_);
  and _50421_ (_42775_, _37507_, _42458_);
  or _50422_ (_42777_, _42775_, _36014_);
  or _50423_ (_42779_, _42777_, _37384_);
  and _50424_ (_42781_, _37507_, _36464_);
  or _50425_ (_42783_, _42682_, _42781_);
  or _50426_ (_42785_, _42783_, _42779_);
  or _50427_ (_42787_, _42785_, _42773_);
  or _50428_ (_42789_, _42787_, _42763_);
  or _50429_ (_42790_, _42789_, _42751_);
  and _50430_ (_42791_, _42790_, _42324_);
  or _50431_ (_30481_, _42791_, _42735_);
  or _50432_ (_42792_, _42438_, _37307_);
  or _50433_ (_42793_, _42519_, _42517_);
  or _50434_ (_42794_, _42793_, _42792_);
  or _50435_ (_42795_, _42794_, _42516_);
  or _50436_ (_42796_, _42795_, _42684_);
  or _50437_ (_42797_, _42757_, _42781_);
  or _50438_ (_42798_, _42743_, _42704_);
  or _50439_ (_42799_, _42798_, _42797_);
  or _50440_ (_42800_, _42523_, _36485_);
  or _50441_ (_42801_, _42800_, _35893_);
  or _50442_ (_42802_, _42629_, _37475_);
  or _50443_ (_42803_, _42802_, _42801_);
  or _50444_ (_42804_, _42803_, _42799_);
  or _50445_ (_42805_, _42804_, _42796_);
  and _50446_ (_42806_, _42805_, _42324_);
  and _50447_ (_42807_, _33817_, _41806_);
  and _50448_ (_42808_, _42807_, _37855_);
  and _50449_ (_42809_, _42418_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _50450_ (_42810_, _42809_, _42808_);
  or _50451_ (_30483_, _42810_, _42806_);
  and _50452_ (_42811_, _36464_, _35871_);
  or _50453_ (_42812_, _42767_, _42438_);
  or _50454_ (_42813_, _42812_, _42811_);
  or _50455_ (_42814_, _42462_, _37296_);
  nor _50456_ (_42815_, _42814_, _42539_);
  nand _50457_ (_42816_, _42815_, _36058_);
  or _50458_ (_42817_, _42816_, _42813_);
  not _50459_ (_42818_, _37454_);
  nor _50460_ (_42819_, _42622_, _37464_);
  and _50461_ (_42820_, _42819_, _42818_);
  not _50462_ (_42821_, _42820_);
  or _50463_ (_42822_, _42821_, _42460_);
  or _50464_ (_42823_, _42822_, _42817_);
  and _50465_ (_42824_, _36453_, _37208_);
  or _50466_ (_42825_, _42824_, _42632_);
  and _50467_ (_42826_, _42461_, _34793_);
  or _50468_ (_42827_, _42826_, _35839_);
  or _50469_ (_42828_, _42827_, _42695_);
  or _50470_ (_42829_, _42828_, _42825_);
  or _50471_ (_42830_, _42829_, _42456_);
  or _50472_ (_42831_, _42830_, _42823_);
  and _50473_ (_42832_, _42831_, _33860_);
  and _50474_ (_42833_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50475_ (_42834_, _42833_, _42542_);
  or _50476_ (_42835_, _42834_, _42832_);
  and _50477_ (_30485_, _42835_, _41806_);
  nor _50478_ (_42836_, _42827_, _42825_);
  nand _50479_ (_42837_, _42836_, _42819_);
  or _50480_ (_42838_, _36036_, _35926_);
  nor _50481_ (_42839_, _42838_, _42741_);
  nand _50482_ (_42840_, _42839_, _40330_);
  or _50483_ (_42841_, _42759_, _42502_);
  or _50484_ (_42842_, _42841_, _42840_);
  or _50485_ (_42843_, _42460_, _42454_);
  or _50486_ (_42844_, _42843_, _42842_);
  or _50487_ (_42845_, _42844_, _42837_);
  and _50488_ (_42846_, _42845_, _33860_);
  and _50489_ (_42847_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50490_ (_42848_, _42847_, _42543_);
  or _50491_ (_42849_, _42848_, _42846_);
  and _50492_ (_30487_, _42849_, _41806_);
  and _50493_ (_42850_, _42418_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _50494_ (_42851_, _36442_);
  and _50495_ (_42852_, _42851_, _37208_);
  or _50496_ (_42853_, _42852_, _37125_);
  or _50497_ (_42854_, _42765_, _42426_);
  or _50498_ (_42855_, _42854_, _42853_);
  or _50499_ (_42856_, _42797_, _42753_);
  or _50500_ (_42857_, _42856_, _42855_);
  or _50501_ (_42858_, _42747_, _42538_);
  or _50502_ (_42859_, _42858_, _42739_);
  or _50503_ (_42860_, _42859_, _42857_);
  and _50504_ (_42861_, _42860_, _42324_);
  or _50505_ (_30489_, _42861_, _42850_);
  nor _50506_ (_38811_, _34233_, rst);
  nor _50507_ (_38813_, _40321_, rst);
  and _50508_ (_42862_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _50509_ (_42864_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _50510_ (_42865_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _50511_ (_42866_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _50512_ (_42867_, _42866_, _42865_);
  and _50513_ (_42868_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _50514_ (_42869_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _50515_ (_42870_, _42869_, _42868_);
  and _50516_ (_42871_, _42870_, _42867_);
  and _50517_ (_42872_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _50518_ (_42873_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _50519_ (_42874_, _42873_, _42872_);
  and _50520_ (_42876_, _42874_, _42871_);
  nor _50521_ (_42877_, _42876_, _33915_);
  nor _50522_ (_42878_, _42877_, _42864_);
  nor _50523_ (_42879_, _42878_, _40305_);
  nor _50524_ (_42880_, _42879_, _42862_);
  nor _50525_ (_38814_, _42880_, rst);
  nor _50526_ (_38825_, _36365_, rst);
  and _50527_ (_38826_, _35012_, _41806_);
  nor _50528_ (_38827_, _35242_, rst);
  nor _50529_ (_38828_, _35496_, rst);
  and _50530_ (_38829_, _35751_, _41806_);
  nor _50531_ (_38830_, _34486_, rst);
  nor _50532_ (_38831_, _34727_, rst);
  nor _50533_ (_38832_, _40396_, rst);
  nor _50534_ (_38834_, _40606_, rst);
  nor _50535_ (_38835_, _40479_, rst);
  nor _50536_ (_38836_, _40356_, rst);
  nor _50537_ (_38837_, _40527_, rst);
  nor _50538_ (_38838_, _40458_, rst);
  nor _50539_ (_38840_, _40682_, rst);
  and _50540_ (_42881_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _50541_ (_42882_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _50542_ (_42883_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _50543_ (_42884_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _50544_ (_42885_, _42884_, _42883_);
  and _50545_ (_42886_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _50546_ (_42887_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _50547_ (_42888_, _42887_, _42886_);
  and _50548_ (_42889_, _42888_, _42885_);
  and _50549_ (_42890_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _50550_ (_42891_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _50551_ (_42892_, _42891_, _42890_);
  and _50552_ (_42893_, _42892_, _42889_);
  nor _50553_ (_42894_, _42893_, _33915_);
  nor _50554_ (_42895_, _42894_, _42882_);
  nor _50555_ (_42896_, _42895_, _40305_);
  nor _50556_ (_42897_, _42896_, _42881_);
  nor _50557_ (_38841_, _42897_, rst);
  and _50558_ (_42898_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _50559_ (_42899_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _50560_ (_42900_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _50561_ (_42901_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _50562_ (_42902_, _42901_, _42900_);
  and _50563_ (_42903_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _50564_ (_42904_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _50565_ (_42905_, _42904_, _42903_);
  and _50566_ (_42906_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _50567_ (_42907_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _50568_ (_42908_, _42907_, _42906_);
  and _50569_ (_42909_, _42908_, _42905_);
  and _50570_ (_42910_, _42909_, _42902_);
  nor _50571_ (_42911_, _42910_, _33915_);
  nor _50572_ (_42912_, _42911_, _42899_);
  nor _50573_ (_42913_, _42912_, _40305_);
  nor _50574_ (_42914_, _42913_, _42898_);
  nor _50575_ (_38842_, _42914_, rst);
  and _50576_ (_42915_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _50577_ (_42916_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _50578_ (_42917_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _50579_ (_42918_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _50580_ (_42919_, _42918_, _42917_);
  and _50581_ (_42920_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _50582_ (_42921_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _50583_ (_42922_, _42921_, _42920_);
  and _50584_ (_42923_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _50585_ (_42924_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _50586_ (_42925_, _42924_, _42923_);
  and _50587_ (_42926_, _42925_, _42922_);
  and _50588_ (_42927_, _42926_, _42919_);
  nor _50589_ (_42928_, _42927_, _33915_);
  nor _50590_ (_42929_, _42928_, _42916_);
  nor _50591_ (_42930_, _42929_, _40305_);
  nor _50592_ (_42931_, _42930_, _42915_);
  nor _50593_ (_38843_, _42931_, rst);
  and _50594_ (_42932_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _50595_ (_42933_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _50596_ (_42934_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _50597_ (_42935_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _50598_ (_42936_, _42935_, _42934_);
  and _50599_ (_42937_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _50600_ (_42938_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _50601_ (_42939_, _42938_, _42937_);
  and _50602_ (_42940_, _42939_, _42936_);
  and _50603_ (_42941_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _50604_ (_42942_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _50605_ (_42943_, _42942_, _42941_);
  and _50606_ (_42944_, _42943_, _42940_);
  nor _50607_ (_42945_, _42944_, _33915_);
  nor _50608_ (_42946_, _42945_, _42933_);
  nor _50609_ (_42947_, _42946_, _40305_);
  nor _50610_ (_42948_, _42947_, _42932_);
  nor _50611_ (_38844_, _42948_, rst);
  and _50612_ (_42949_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _50613_ (_42950_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _50614_ (_42951_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _50615_ (_42952_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _50616_ (_42953_, _42952_, _42951_);
  and _50617_ (_42954_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _50618_ (_42955_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _50619_ (_42956_, _42955_, _42954_);
  and _50620_ (_42957_, _42956_, _42953_);
  and _50621_ (_42958_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _50622_ (_42959_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _50623_ (_42960_, _42959_, _42958_);
  and _50624_ (_42961_, _42960_, _42957_);
  nor _50625_ (_42962_, _42961_, _33915_);
  nor _50626_ (_42963_, _42962_, _42950_);
  nor _50627_ (_42964_, _42963_, _40305_);
  nor _50628_ (_42965_, _42964_, _42949_);
  nor _50629_ (_38846_, _42965_, rst);
  and _50630_ (_42966_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _50631_ (_42967_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _50632_ (_42968_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _50633_ (_42969_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _50634_ (_42970_, _42969_, _42968_);
  and _50635_ (_42971_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _50636_ (_42972_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _50637_ (_42973_, _42972_, _42971_);
  and _50638_ (_42974_, _42973_, _42970_);
  and _50639_ (_42975_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _50640_ (_42976_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _50641_ (_42977_, _42976_, _42975_);
  and _50642_ (_42978_, _42977_, _42974_);
  nor _50643_ (_42979_, _42978_, _33915_);
  nor _50644_ (_42980_, _42979_, _42967_);
  nor _50645_ (_42981_, _42980_, _40305_);
  nor _50646_ (_42982_, _42981_, _42966_);
  nor _50647_ (_38847_, _42982_, rst);
  and _50648_ (_42983_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _50649_ (_42984_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _50650_ (_42985_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _50651_ (_42986_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _50652_ (_42987_, _42986_, _42985_);
  and _50653_ (_42988_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _50654_ (_42989_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _50655_ (_42990_, _42989_, _42988_);
  and _50656_ (_42991_, _42990_, _42987_);
  and _50657_ (_42992_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _50658_ (_42993_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _50659_ (_42994_, _42993_, _42992_);
  and _50660_ (_42995_, _42994_, _42991_);
  nor _50661_ (_42996_, _42995_, _33915_);
  nor _50662_ (_42997_, _42996_, _42984_);
  nor _50663_ (_42998_, _42997_, _40305_);
  nor _50664_ (_42999_, _42998_, _42983_);
  nor _50665_ (_38848_, _42999_, rst);
  and _50666_ (_43000_, _33881_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _50667_ (_43001_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _50668_ (_43002_, _43000_, _38571_);
  and _50669_ (_43003_, _43002_, _41806_);
  and _50670_ (_38872_, _43003_, _43001_);
  not _50671_ (_43004_, _43000_);
  or _50672_ (_43005_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _50673_ (_00000_, _43000_, _41806_);
  and _50674_ (_43006_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _41806_);
  or _50675_ (_43007_, _43006_, _00000_);
  and _50676_ (_38874_, _43007_, _43005_);
  nor _50677_ (_38911_, _40327_, rst);
  and _50678_ (_38913_, _40544_, _41806_);
  nor _50679_ (_38914_, _40300_, rst);
  nor _50680_ (_43008_, _40327_, _24949_);
  and _50681_ (_43009_, _40327_, _24949_);
  nor _50682_ (_43010_, _43009_, _43008_);
  nor _50683_ (_43011_, _40703_, _24665_);
  and _50684_ (_43012_, _40703_, _24665_);
  nor _50685_ (_43013_, _43012_, _43011_);
  nor _50686_ (_43014_, _43013_, _43010_);
  nor _50687_ (_43015_, _40380_, _25112_);
  and _50688_ (_43016_, _40380_, _25112_);
  nor _50689_ (_43017_, _43016_, _43015_);
  not _50690_ (_43018_, _43017_);
  and _50691_ (_43019_, _40547_, _40614_);
  nor _50692_ (_43020_, _40547_, _40614_);
  nor _50693_ (_43021_, _43020_, _43019_);
  nor _50694_ (_43022_, _40463_, _24796_);
  and _50695_ (_43023_, _40463_, _24796_);
  nor _50696_ (_43024_, _43023_, _43022_);
  nor _50697_ (_43025_, _43024_, _43021_);
  and _50698_ (_43026_, _43025_, _43018_);
  and _50699_ (_43027_, _43026_, _43014_);
  nor _50700_ (_43028_, _37539_, _42442_);
  and _50701_ (_43029_, _38853_, _28087_);
  and _50702_ (_43030_, _43029_, _43028_);
  and _50703_ (_43031_, _43030_, _43027_);
  nor _50704_ (_43032_, _25984_, _25593_);
  and _50705_ (_43033_, _43032_, _28872_);
  and _50706_ (_43034_, _43033_, _30240_);
  nand _50707_ (_43035_, _43034_, _30914_);
  nor _50708_ (_43036_, _43035_, _31652_);
  and _50709_ (_43037_, _43036_, _32393_);
  nor _50710_ (_43038_, _43028_, _37668_);
  and _50711_ (_43039_, _43038_, _43037_);
  and _50712_ (_43040_, _43039_, _26604_);
  and _50713_ (_43041_, _43028_, _26354_);
  not _50714_ (_43042_, _37668_);
  nor _50715_ (_43043_, _43028_, _34530_);
  nor _50716_ (_43044_, _43043_, _43042_);
  and _50717_ (_43045_, _43044_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _50718_ (_43046_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _50719_ (_43047_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _50720_ (_43048_, _43047_, _43046_);
  nor _50721_ (_43049_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _50722_ (_43050_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _50723_ (_43051_, _43050_, _43049_);
  and _50724_ (_43052_, _43051_, _43048_);
  and _50725_ (_43053_, _43052_, _36771_);
  or _50726_ (_43054_, _43053_, _43045_);
  or _50727_ (_43055_, _43054_, _43041_);
  nor _50728_ (_43056_, _43055_, _43040_);
  not _50729_ (_43057_, _42494_);
  nor _50730_ (_43058_, _42694_, _37263_);
  and _50731_ (_43059_, _43058_, _43057_);
  or _50732_ (_43060_, _37507_, _36518_);
  or _50733_ (_43061_, _43060_, _36990_);
  and _50734_ (_43062_, _43061_, _36584_);
  nor _50735_ (_43063_, _43062_, _42651_);
  nand _50736_ (_43064_, _43063_, _43059_);
  and _50737_ (_43065_, _43064_, _43056_);
  nand _50738_ (_43066_, _37657_, _35795_);
  and _50739_ (_43067_, _43066_, _37723_);
  or _50740_ (_43068_, _43067_, _43056_);
  nor _50741_ (_43069_, _42423_, _36529_);
  nand _50742_ (_43070_, _43069_, _43068_);
  or _50743_ (_43071_, _43070_, _43065_);
  and _50744_ (_43072_, _43071_, _36749_);
  and _50745_ (_43073_, _36628_, _35915_);
  nor _50746_ (_43074_, _43073_, _42481_);
  nor _50747_ (_43075_, _43074_, _33817_);
  nor _50748_ (_43076_, _43075_, _36781_);
  not _50749_ (_43077_, _43076_);
  nor _50750_ (_43078_, _43077_, _43072_);
  nor _50751_ (_43079_, _38955_, _38823_);
  and _50752_ (_43080_, _43079_, _38860_);
  not _50753_ (_43081_, _43080_);
  and _50754_ (_43082_, _43081_, _43044_);
  not _50755_ (_43083_, _39080_);
  and _50756_ (_43084_, _43083_, _36771_);
  nor _50757_ (_43085_, _43084_, _43082_);
  not _50758_ (_43086_, _43085_);
  nor _50759_ (_43087_, _43086_, _43078_);
  not _50760_ (_43088_, _43087_);
  nor _50761_ (_43089_, _43088_, _43031_);
  and _50762_ (_43090_, _40611_, _30686_);
  nor _50763_ (_43091_, _40611_, _30686_);
  or _50764_ (_43092_, _43091_, _43090_);
  nand _50765_ (_43093_, _43018_, _28076_);
  nor _50766_ (_43094_, _40415_, _24434_);
  and _50767_ (_43095_, _40415_, _24434_);
  nor _50768_ (_43096_, _43095_, _43094_);
  nor _50769_ (_43097_, _40500_, _24197_);
  and _50770_ (_43098_, _40500_, _24197_);
  nor _50771_ (_43099_, _43098_, _43097_);
  or _50772_ (_43100_, _43099_, _43096_);
  or _50773_ (_43101_, _43100_, _43093_);
  nor _50774_ (_43102_, _43101_, _43092_);
  and _50775_ (_43103_, _43102_, _43025_);
  and _50776_ (_43104_, _43103_, _43014_);
  nor _50777_ (_43105_, _24949_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _50778_ (_43106_, _43105_, _43104_);
  not _50779_ (_43107_, _43106_);
  and _50780_ (_43108_, _43107_, _43089_);
  and _50781_ (_43109_, _43108_, _37635_);
  and _50782_ (_38918_, _43109_, _41806_);
  and _50783_ (_38919_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _41806_);
  and _50784_ (_38920_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _41806_);
  nor _50785_ (_43110_, _37635_, _28011_);
  and _50786_ (_43111_, _36749_, _36529_);
  not _50787_ (_43112_, _43111_);
  nor _50788_ (_43113_, _43112_, _38582_);
  and _50789_ (_43114_, _43073_, _36858_);
  and _50790_ (_43115_, _43114_, _40322_);
  and _50791_ (_43116_, _42650_, _37539_);
  and _50792_ (_43117_, _43116_, _43058_);
  nor _50793_ (_43118_, _43117_, _37679_);
  nor _50794_ (_43119_, _43114_, _37624_);
  not _50795_ (_43120_, _43119_);
  nor _50796_ (_43121_, _43120_, _43118_);
  nor _50797_ (_43122_, _43111_, _43075_);
  and _50798_ (_43123_, _43122_, _43121_);
  and _50799_ (_43124_, _36584_, _36858_);
  and _50800_ (_43125_, _43124_, _35871_);
  not _50801_ (_43126_, _37657_);
  and _50802_ (_43127_, _43069_, _43126_);
  and _50803_ (_43128_, _43127_, _43059_);
  and _50804_ (_43129_, _43128_, _43116_);
  nor _50805_ (_43130_, _43129_, _37679_);
  nor _50806_ (_43131_, _43130_, _43125_);
  and _50807_ (_43132_, _43131_, _43123_);
  and _50808_ (_43134_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _50809_ (_43135_, _43134_, _43115_);
  or _50810_ (_43136_, _43135_, _43113_);
  or _50811_ (_43137_, _43136_, _43110_);
  not _50812_ (_43138_, _42880_);
  and _50813_ (_43140_, _37485_, _36858_);
  not _50814_ (_43141_, _43140_);
  and _50815_ (_43142_, _43141_, _43121_);
  nor _50816_ (_43143_, _43142_, _43138_);
  and _50817_ (_43144_, _43142_, _40321_);
  nor _50818_ (_43146_, _43144_, _43143_);
  and _50819_ (_43147_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _50820_ (_43148_, _43147_);
  nor _50821_ (_43149_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _50822_ (_43150_, _43149_, _43147_);
  not _50823_ (_43152_, _42999_);
  nor _50824_ (_43153_, _43142_, _43152_);
  and _50825_ (_43154_, _43142_, _40682_);
  nor _50826_ (_43155_, _43154_, _43153_);
  and _50827_ (_43156_, _43155_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _50828_ (_43158_, _43155_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _50829_ (_43159_, _43158_, _43156_);
  not _50830_ (_43160_, _42982_);
  nor _50831_ (_43161_, _43142_, _43160_);
  and _50832_ (_43162_, _43142_, _40458_);
  nor _50833_ (_43164_, _43162_, _43161_);
  and _50834_ (_43165_, _43164_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _50835_ (_43166_, _43164_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _50836_ (_43167_, _42965_);
  nor _50837_ (_43168_, _43142_, _43167_);
  and _50838_ (_43170_, _43142_, _40527_);
  nor _50839_ (_43171_, _43170_, _43168_);
  nand _50840_ (_43173_, _43171_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _50841_ (_43174_, _42948_);
  nor _50842_ (_43175_, _43142_, _43174_);
  and _50843_ (_43176_, _43142_, _40356_);
  nor _50844_ (_43177_, _43176_, _43175_);
  and _50845_ (_43178_, _43177_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _50846_ (_43179_, _43177_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _50847_ (_43181_, _42931_);
  nor _50848_ (_43182_, _43142_, _43181_);
  and _50849_ (_43183_, _43142_, _40479_);
  nor _50850_ (_43185_, _43183_, _43182_);
  and _50851_ (_43186_, _43185_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _50852_ (_43187_, _42914_);
  nor _50853_ (_43189_, _43142_, _43187_);
  and _50854_ (_43190_, _43142_, _40606_);
  nor _50855_ (_43191_, _43190_, _43189_);
  and _50856_ (_43193_, _43191_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _50857_ (_43194_, _42897_);
  nor _50858_ (_43195_, _43142_, _43194_);
  and _50859_ (_43197_, _43142_, _40396_);
  nor _50860_ (_43198_, _43197_, _43195_);
  and _50861_ (_43199_, _43198_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _50862_ (_43201_, _43191_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _50863_ (_43202_, _43201_, _43193_);
  and _50864_ (_43203_, _43202_, _43199_);
  nor _50865_ (_43205_, _43203_, _43193_);
  not _50866_ (_43206_, _43205_);
  nor _50867_ (_43208_, _43185_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _50868_ (_43209_, _43208_, _43186_);
  and _50869_ (_43210_, _43209_, _43206_);
  nor _50870_ (_43211_, _43210_, _43186_);
  nor _50871_ (_43212_, _43211_, _43179_);
  or _50872_ (_43213_, _43212_, _43178_);
  or _50873_ (_43214_, _43171_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _50874_ (_43216_, _43214_, _43173_);
  nand _50875_ (_43217_, _43216_, _43213_);
  and _50876_ (_43218_, _43217_, _43173_);
  nor _50877_ (_43220_, _43218_, _43166_);
  or _50878_ (_43221_, _43220_, _43165_);
  and _50879_ (_43222_, _43221_, _43159_);
  nor _50880_ (_43224_, _43222_, _43156_);
  not _50881_ (_43225_, _43224_);
  nand _50882_ (_43226_, _43225_, _43150_);
  and _50883_ (_43228_, _43226_, _43148_);
  nor _50884_ (_43229_, _43228_, _38543_);
  and _50885_ (_43230_, _43229_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _50886_ (_43232_, _43230_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _50887_ (_43233_, _43232_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _50888_ (_43234_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _50889_ (_43236_, _43234_, _43233_);
  nor _50890_ (_43237_, _43236_, _43146_);
  not _50891_ (_43238_, _43146_);
  and _50892_ (_43240_, _43228_, _38543_);
  and _50893_ (_43241_, _43240_, _38549_);
  and _50894_ (_43243_, _43241_, _38554_);
  and _50895_ (_43244_, _43243_, _38539_);
  nor _50896_ (_43245_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _50897_ (_43246_, _43245_, _43244_);
  nor _50898_ (_43247_, _43246_, _43238_);
  nor _50899_ (_43249_, _43247_, _43237_);
  or _50900_ (_43250_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _50901_ (_43251_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _50902_ (_43253_, _43251_, _43250_);
  and _50903_ (_43254_, _43253_, _43249_);
  or _50904_ (_43255_, _43254_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _50905_ (_43257_, _43254_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _50906_ (_43258_, _43122_);
  and _50907_ (_43259_, _43258_, _43142_);
  nor _50908_ (_43261_, _43131_, _43259_);
  and _50909_ (_43262_, _43261_, _43257_);
  and _50910_ (_43263_, _43262_, _43255_);
  or _50911_ (_43265_, _43263_, _43137_);
  and _50912_ (_43266_, _43121_, _43075_);
  and _50913_ (_43267_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _50914_ (_43269_, _43267_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _50915_ (_43270_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _50916_ (_43271_, _43270_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _50917_ (_43273_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _50918_ (_43274_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _50919_ (_43276_, _43274_, _43273_);
  and _50920_ (_43277_, _43276_, _43271_);
  and _50921_ (_43278_, _43277_, _43269_);
  and _50922_ (_43279_, _43278_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _50923_ (_43280_, _43279_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _50924_ (_43281_, _43280_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _50925_ (_43282_, _43281_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _50926_ (_43284_, _43282_, _38571_);
  or _50927_ (_43285_, _43282_, _38571_);
  and _50928_ (_43286_, _43285_, _43284_);
  nand _50929_ (_43288_, _43286_, _43266_);
  nand _50930_ (_43289_, _43288_, _43108_);
  or _50931_ (_43290_, _43289_, _43265_);
  not _50932_ (_43292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _50933_ (_43293_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _50934_ (_43294_, _43293_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _50935_ (_43296_, _43294_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _50936_ (_43297_, _43296_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _50937_ (_43298_, _43297_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _50938_ (_43300_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _50939_ (_43301_, _43300_, _43298_);
  and _50940_ (_43302_, _43301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _50941_ (_43304_, _43302_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _50942_ (_43305_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _50943_ (_43306_, _34036_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _50944_ (_43308_, _43306_, _40305_);
  nor _50945_ (_43309_, _43308_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _50946_ (_43311_, _43309_);
  and _50947_ (_43312_, _43311_, _43305_);
  and _50948_ (_43313_, _43312_, _43304_);
  nand _50949_ (_43314_, _43313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _50950_ (_43316_, _43314_, _43292_);
  or _50951_ (_43317_, _43314_, _43292_);
  and _50952_ (_43318_, _43317_, _43316_);
  or _50953_ (_43320_, _43318_, _43108_);
  and _50954_ (_43321_, _43320_, _41806_);
  and _50955_ (_38922_, _43321_, _43290_);
  and _50956_ (_43323_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _41806_);
  and _50957_ (_43324_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _50958_ (_43325_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _50959_ (_43327_, _33860_, _43325_);
  not _50960_ (_43328_, _43327_);
  not _50961_ (_43329_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _50962_ (_43331_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _50963_ (_43332_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _50964_ (_43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _50965_ (_43335_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _50966_ (_43336_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _50967_ (_43337_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _50968_ (_43339_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _50969_ (_43340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _50970_ (_43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _50971_ (_43343_, _43342_, _43340_);
  and _50972_ (_43344_, _43343_, _43339_);
  and _50973_ (_43345_, _43344_, _43337_);
  and _50974_ (_43347_, _43345_, _43336_);
  and _50975_ (_43348_, _43347_, _43335_);
  and _50976_ (_43349_, _43348_, _43333_);
  and _50977_ (_43351_, _43349_, _43332_);
  and _50978_ (_43352_, _43351_, _43331_);
  and _50979_ (_43353_, _43352_, _43329_);
  nor _50980_ (_43355_, _43353_, _43292_);
  and _50981_ (_43356_, _43353_, _43292_);
  nor _50982_ (_43357_, _43356_, _43355_);
  nor _50983_ (_43359_, _43352_, _43329_);
  or _50984_ (_43360_, _43359_, _43353_);
  and _50985_ (_43361_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _50986_ (_43363_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _50987_ (_43364_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _50988_ (_43365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _50989_ (_43367_, _43365_, _43363_);
  and _50990_ (_43368_, _43367_, _43364_);
  nor _50991_ (_43369_, _43368_, _43363_);
  nor _50992_ (_43371_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _50993_ (_43372_, _43371_, _43361_);
  not _50994_ (_43374_, _43372_);
  nor _50995_ (_43375_, _43374_, _43369_);
  nor _50996_ (_43376_, _43375_, _43361_);
  not _50997_ (_43377_, _43376_);
  and _50998_ (_43379_, _43377_, _43349_);
  and _50999_ (_43380_, _43379_, _43332_);
  and _51000_ (_43381_, _43380_, _43331_);
  and _51001_ (_43383_, _43381_, _43360_);
  nor _51002_ (_43384_, _43381_, _43360_);
  or _51003_ (_43385_, _43384_, _43383_);
  not _51004_ (_43387_, _43385_);
  and _51005_ (_43388_, _43376_, _43352_);
  and _51006_ (_43389_, _43376_, _43351_);
  nor _51007_ (_43391_, _43389_, _43331_);
  nor _51008_ (_43392_, _43391_, _43388_);
  not _51009_ (_43393_, _43392_);
  and _51010_ (_43395_, _43376_, _43349_);
  nor _51011_ (_43396_, _43395_, _43332_);
  nor _51012_ (_43397_, _43396_, _43389_);
  not _51013_ (_43399_, _43397_);
  and _51014_ (_43400_, _43376_, _43347_);
  and _51015_ (_43401_, _43400_, _43335_);
  nor _51016_ (_43403_, _43401_, _43333_);
  nor _51017_ (_43404_, _43403_, _43395_);
  not _51018_ (_43406_, _43404_);
  nor _51019_ (_43407_, _43400_, _43335_);
  nor _51020_ (_43408_, _43407_, _43401_);
  not _51021_ (_43409_, _43408_);
  not _51022_ (_43410_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _51023_ (_43411_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _51024_ (_43412_, _43376_, _43345_);
  and _51025_ (_43414_, _43412_, _43411_);
  nor _51026_ (_43415_, _43414_, _43410_);
  nor _51027_ (_43416_, _43415_, _43400_);
  not _51028_ (_43418_, _43416_);
  and _51029_ (_43419_, _43376_, _43343_);
  and _51030_ (_43420_, _43419_, _43339_);
  nor _51031_ (_43422_, _43420_, _43337_);
  nor _51032_ (_43423_, _43422_, _43412_);
  not _51033_ (_43424_, _43423_);
  nor _51034_ (_43426_, _43419_, _43339_);
  nor _51035_ (_43427_, _43426_, _43420_);
  not _51036_ (_43428_, _43427_);
  and _51037_ (_43430_, _43376_, _43342_);
  nor _51038_ (_43431_, _43430_, _43340_);
  nor _51039_ (_43432_, _43431_, _43419_);
  not _51040_ (_43434_, _43432_);
  not _51041_ (_43435_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _51042_ (_43436_, _43376_, _43435_);
  nor _51043_ (_43438_, _43376_, _43435_);
  nor _51044_ (_43439_, _43438_, _43436_);
  not _51045_ (_43441_, _43439_);
  nor _51046_ (_43442_, _42372_, _42340_);
  not _51047_ (_43443_, _42372_);
  nor _51048_ (_43444_, _42367_, _42355_);
  nor _51049_ (_43446_, _43444_, _43443_);
  nor _51050_ (_43447_, _43446_, _42396_);
  or _51051_ (_43448_, _43447_, _43442_);
  and _51052_ (_43450_, _42354_, _42366_);
  not _51053_ (_43451_, _43450_);
  nor _51054_ (_43452_, _42372_, _42368_);
  nor _51055_ (_43454_, _43452_, _43451_);
  not _51056_ (_43455_, _42369_);
  and _51057_ (_43456_, _42387_, _42330_);
  nor _51058_ (_43458_, _43456_, _42348_);
  nor _51059_ (_43459_, _43458_, _43455_);
  nor _51060_ (_43460_, _43459_, _43454_);
  and _51061_ (_43462_, _43460_, _43448_);
  and _51062_ (_43463_, _42343_, _42330_);
  nor _51063_ (_43464_, _43463_, _42359_);
  nor _51064_ (_43466_, _43464_, _43443_);
  and _51065_ (_43467_, _42372_, _42334_);
  and _51066_ (_43468_, _43467_, _42345_);
  nor _51067_ (_43470_, _43468_, _43466_);
  and _51068_ (_43471_, _42396_, _42357_);
  nor _51069_ (_43473_, _43471_, _42364_);
  not _51070_ (_43474_, _43473_);
  not _51071_ (_43475_, _42361_);
  and _51072_ (_43476_, _42335_, _35496_);
  and _51073_ (_43478_, _43476_, _42334_);
  and _51074_ (_43479_, _42354_, _42329_);
  and _51075_ (_43483_, _35751_, _35496_);
  and _51076_ (_43489_, _43483_, _43479_);
  nor _51077_ (_43490_, _43489_, _43478_);
  nor _51078_ (_43503_, _43490_, _43475_);
  nor _51079_ (_43508_, _43503_, _43474_);
  and _51080_ (_43509_, _43508_, _43470_);
  and _51081_ (_43523_, _43509_, _43462_);
  and _51082_ (_43528_, _42359_, _42340_);
  not _51083_ (_43529_, _43528_);
  nor _51084_ (_43541_, _42370_, _42350_);
  and _51085_ (_43548_, _43541_, _43529_);
  nor _51086_ (_43549_, _42355_, _42376_);
  nor _51087_ (_43559_, _43549_, _43455_);
  not _51088_ (_43568_, _43559_);
  not _51089_ (_43569_, _42368_);
  and _51090_ (_43577_, _42366_, _42334_);
  nor _51091_ (_43586_, _43577_, _42388_);
  nor _51092_ (_43587_, _43586_, _43569_);
  not _51093_ (_43597_, _42347_);
  and _51094_ (_43598_, _42387_, _42334_);
  and _51095_ (_43605_, _42330_, _34486_);
  nor _51096_ (_43616_, _43605_, _43598_);
  nor _51097_ (_43622_, _43616_, _43597_);
  nor _51098_ (_43623_, _43622_, _43587_);
  and _51099_ (_43636_, _43623_, _43568_);
  and _51100_ (_43641_, _43636_, _43548_);
  and _51101_ (_43642_, _43641_, _43523_);
  not _51102_ (_43656_, _43598_);
  and _51103_ (_43661_, _43549_, _43656_);
  nor _51104_ (_43662_, _43661_, _35496_);
  not _51105_ (_43668_, _43662_);
  and _51106_ (_43680_, _42344_, _42330_);
  not _51107_ (_43681_, _43680_);
  nor _51108_ (_43693_, _43463_, _42396_);
  and _51109_ (_43700_, _43693_, _43681_);
  nor _51110_ (_43701_, _43700_, _43455_);
  not _51111_ (_43711_, _43701_);
  and _51112_ (_43720_, _43711_, _42399_);
  and _51113_ (_43721_, _43720_, _43668_);
  and _51114_ (_43722_, _43467_, _42343_);
  not _51115_ (_43724_, _43722_);
  and _51116_ (_43725_, _43724_, _42379_);
  and _51117_ (_43727_, _42369_, _42359_);
  and _51118_ (_43728_, _43450_, _42357_);
  nor _51119_ (_43729_, _43728_, _43727_);
  and _51120_ (_43730_, _42371_, _42341_);
  not _51121_ (_43731_, _43730_);
  and _51122_ (_43733_, _43731_, _43729_);
  and _51123_ (_43734_, _43733_, _43725_);
  and _51124_ (_43735_, _42394_, _42340_);
  not _51125_ (_43737_, _43735_);
  and _51126_ (_43738_, _42388_, _42328_);
  and _51127_ (_43739_, _42355_, _42340_);
  nor _51128_ (_43741_, _43739_, _43738_);
  and _51129_ (_43742_, _43741_, _43737_);
  and _51130_ (_43743_, _43577_, _42347_);
  and _51131_ (_43745_, _42359_, _42347_);
  nor _51132_ (_43746_, _43745_, _43743_);
  and _51133_ (_43747_, _43746_, _42384_);
  and _51134_ (_43749_, _43747_, _43742_);
  and _51135_ (_43750_, _43749_, _43734_);
  and _51136_ (_43751_, _43750_, _43721_);
  and _51137_ (_43753_, _43751_, _43642_);
  nor _51138_ (_43754_, _43367_, _43364_);
  nor _51139_ (_43755_, _43754_, _43368_);
  not _51140_ (_43757_, _43755_);
  nor _51141_ (_43758_, _43757_, _43753_);
  and _51142_ (_43760_, _43729_, _43548_);
  nor _51143_ (_43761_, _42383_, _42364_);
  and _51144_ (_43762_, _43761_, _43568_);
  nor _51145_ (_43763_, _43471_, _42395_);
  and _51146_ (_43765_, _42388_, _42357_);
  nor _51147_ (_43766_, _43765_, _43743_);
  and _51148_ (_43767_, _43766_, _43763_);
  and _51149_ (_43769_, _43767_, _43762_);
  and _51150_ (_43770_, _43769_, _43760_);
  not _51151_ (_43771_, _43770_);
  nor _51152_ (_43773_, _43771_, _43753_);
  not _51153_ (_43774_, _43773_);
  nor _51154_ (_43775_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _51155_ (_43777_, _43775_, _43364_);
  and _51156_ (_43778_, _43777_, _43774_);
  and _51157_ (_43779_, _43757_, _43753_);
  nor _51158_ (_43781_, _43779_, _43758_);
  and _51159_ (_43782_, _43781_, _43778_);
  nor _51160_ (_43783_, _43782_, _43758_);
  not _51161_ (_43785_, _43783_);
  and _51162_ (_43786_, _43374_, _43369_);
  nor _51163_ (_43787_, _43786_, _43375_);
  and _51164_ (_43789_, _43787_, _43785_);
  and _51165_ (_43790_, _43789_, _43441_);
  not _51166_ (_43792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _51167_ (_43793_, _43436_, _43792_);
  or _51168_ (_43794_, _43793_, _43430_);
  and _51169_ (_43795_, _43794_, _43790_);
  and _51170_ (_43797_, _43795_, _43434_);
  and _51171_ (_43798_, _43797_, _43428_);
  and _51172_ (_43799_, _43798_, _43424_);
  nor _51173_ (_43801_, _43412_, _43411_);
  or _51174_ (_43802_, _43801_, _43414_);
  and _51175_ (_43803_, _43802_, _43799_);
  and _51176_ (_43805_, _43803_, _43418_);
  and _51177_ (_43806_, _43805_, _43409_);
  and _51178_ (_43807_, _43806_, _43406_);
  and _51179_ (_43809_, _43807_, _43399_);
  and _51180_ (_43810_, _43809_, _43393_);
  and _51181_ (_43811_, _43810_, _43387_);
  or _51182_ (_43813_, _43811_, _43383_);
  nor _51183_ (_43814_, _43813_, _43357_);
  and _51184_ (_43815_, _43813_, _43357_);
  or _51185_ (_43817_, _43815_, _43814_);
  or _51186_ (_43818_, _43817_, _43328_);
  or _51187_ (_43819_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _51188_ (_43821_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _51189_ (_43822_, _43821_, _43819_);
  and _51190_ (_43824_, _43822_, _43818_);
  or _51191_ (_38923_, _43824_, _43324_);
  nor _51192_ (_43825_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _51193_ (_38924_, _43825_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _51194_ (_38925_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _41806_);
  nor _51195_ (_43827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _51196_ (_43828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _51197_ (_43830_, _43828_, _43827_);
  nor _51198_ (_43831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _51199_ (_43832_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _51200_ (_43834_, _43832_, _43831_);
  and _51201_ (_43835_, _43834_, _43830_);
  nor _51202_ (_43836_, _43835_, rst);
  and _51203_ (_43838_, \oc8051_top_1.oc8051_rom1.ea_int , _33828_);
  nand _51204_ (_43839_, _43838_, _33860_);
  and _51205_ (_43840_, _43839_, _38925_);
  or _51206_ (_38927_, _43840_, _43836_);
  and _51207_ (_43842_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _51208_ (_43843_, _43842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _51209_ (_38928_, _43843_, _41806_);
  nor _51210_ (_43845_, _43309_, _40305_);
  nor _51211_ (_43846_, _43753_, _33981_);
  nor _51212_ (_43848_, _43773_, _34069_);
  and _51213_ (_43849_, _43753_, _33981_);
  nor _51214_ (_43850_, _43849_, _43846_);
  and _51215_ (_43851_, _43850_, _43848_);
  nor _51216_ (_43852_, _43851_, _43846_);
  nor _51217_ (_43853_, _43852_, _40305_);
  and _51218_ (_43854_, _43853_, _33937_);
  nor _51219_ (_43855_, _43853_, _33937_);
  nor _51220_ (_43856_, _43855_, _43854_);
  nor _51221_ (_43857_, _43856_, _43845_);
  and _51222_ (_43858_, _33992_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _51223_ (_43859_, _43858_, _43845_);
  nor _51224_ (_43860_, _43859_, _43770_);
  or _51225_ (_43861_, _43860_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _51226_ (_43862_, _43861_, _43857_);
  and _51227_ (_38929_, _43862_, _41806_);
  not _51228_ (_43863_, _34935_);
  and _51229_ (_43864_, _34190_, _43863_);
  not _51230_ (_43865_, _35685_);
  and _51231_ (_43866_, _43865_, _34683_);
  and _51232_ (_43867_, _43866_, _43864_);
  and _51233_ (_43868_, _33881_, _41806_);
  nand _51234_ (_43869_, _43868_, _35199_);
  nor _51235_ (_43870_, _43869_, _35451_);
  not _51236_ (_43871_, _34442_);
  nor _51237_ (_43872_, _36321_, _43871_);
  and _51238_ (_43873_, _43872_, _43870_);
  and _51239_ (_38932_, _43873_, _43867_);
  nor _51240_ (_43874_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _51241_ (_43875_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _51242_ (_43876_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _51243_ (_38935_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _41806_);
  and _51244_ (_43877_, _38935_, _43876_);
  or _51245_ (_38934_, _43877_, _43875_);
  not _51246_ (_43878_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _51247_ (_43879_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _51248_ (_43880_, _43879_, _43878_);
  and _51249_ (_43881_, _43879_, _43878_);
  nor _51250_ (_43882_, _43881_, _43880_);
  not _51251_ (_43883_, _43882_);
  and _51252_ (_43884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _51253_ (_43885_, _43884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _51254_ (_43886_, _43884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _51255_ (_43887_, _43886_, _43885_);
  or _51256_ (_43888_, _43887_, _43879_);
  and _51257_ (_43889_, _43888_, _43883_);
  nor _51258_ (_43890_, _43880_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _51259_ (_43891_, _43880_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _51260_ (_43892_, _43891_, _43890_);
  or _51261_ (_43893_, _43885_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _51262_ (_38937_, _43893_, _41806_);
  and _51263_ (_43894_, _38937_, _43892_);
  and _51264_ (_38936_, _43894_, _43889_);
  not _51265_ (_43895_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _51266_ (_43896_, _43309_, _43895_);
  and _51267_ (_43897_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _51268_ (_43898_, _43896_);
  and _51269_ (_43899_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _51270_ (_43900_, _43899_, _43897_);
  and _51271_ (_38938_, _43900_, _41806_);
  and _51272_ (_43901_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _51273_ (_43902_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _51274_ (_43903_, _43902_, _43901_);
  and _51275_ (_38939_, _43903_, _41806_);
  and _51276_ (_43904_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _51277_ (_43905_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _51278_ (_43906_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _43905_);
  and _51279_ (_43907_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _51280_ (_43908_, _43907_, _43904_);
  and _51281_ (_38940_, _43908_, _41806_);
  and _51282_ (_43909_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _51283_ (_43910_, _43909_, _43906_);
  and _51284_ (_38941_, _43910_, _41806_);
  or _51285_ (_43911_, _43905_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _51286_ (_38942_, _43911_, _41806_);
  not _51287_ (_43912_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _51288_ (_43913_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _51289_ (_43914_, _43913_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _51290_ (_43915_, _43905_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _51291_ (_43916_, _43915_, _41806_);
  and _51292_ (_38943_, _43916_, _43914_);
  or _51293_ (_43917_, _43905_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _51294_ (_38944_, _43917_, _41806_);
  nor _51295_ (_43918_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _51296_ (_43919_, _43918_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _51297_ (_43920_, _43919_, _41806_);
  and _51298_ (_43921_, _38935_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _51299_ (_38945_, _43921_, _43920_);
  and _51300_ (_43922_, _43895_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _51301_ (_43923_, _43922_, _43919_);
  and _51302_ (_38946_, _43923_, _41806_);
  nand _51303_ (_43924_, _43919_, _38582_);
  or _51304_ (_43925_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _51305_ (_43926_, _43925_, _41806_);
  and _51306_ (_38947_, _43926_, _43924_);
  and _51307_ (_38948_, _37965_, _40269_);
  or _51308_ (_43927_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _51309_ (_43928_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _41806_);
  or _51310_ (_43929_, _43928_, _00000_);
  and _51311_ (_38985_, _43929_, _43927_);
  or _51312_ (_43930_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _51313_ (_43931_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _51314_ (_43932_, _43000_, _43931_);
  and _51315_ (_43933_, _43932_, _41806_);
  and _51316_ (_38986_, _43933_, _43930_);
  or _51317_ (_43934_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _51318_ (_43935_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _51319_ (_43936_, _43000_, _43935_);
  and _51320_ (_43937_, _43936_, _41806_);
  and _51321_ (_38987_, _43937_, _43934_);
  or _51322_ (_43938_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _51323_ (_43939_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _51324_ (_43940_, _43000_, _43939_);
  and _51325_ (_43941_, _43940_, _41806_);
  and _51326_ (_38989_, _43941_, _43938_);
  or _51327_ (_43942_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not _51328_ (_43943_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _51329_ (_43944_, _43000_, _43943_);
  and _51330_ (_43945_, _43944_, _41806_);
  and _51331_ (_38990_, _43945_, _43942_);
  or _51332_ (_43946_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _51333_ (_43947_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _51334_ (_43948_, _43000_, _43947_);
  and _51335_ (_43949_, _43948_, _41806_);
  and _51336_ (_38991_, _43949_, _43946_);
  or _51337_ (_43950_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not _51338_ (_43951_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand _51339_ (_43952_, _43000_, _43951_);
  and _51340_ (_43953_, _43952_, _41806_);
  and _51341_ (_38992_, _43953_, _43950_);
  or _51342_ (_43954_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _51343_ (_43955_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand _51344_ (_43956_, _43000_, _43955_);
  and _51345_ (_43957_, _43956_, _41806_);
  and _51346_ (_38993_, _43957_, _43954_);
  or _51347_ (_43958_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _51348_ (_43959_, _43000_, _38543_);
  and _51349_ (_43960_, _43959_, _41806_);
  and _51350_ (_38994_, _43960_, _43958_);
  or _51351_ (_43961_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _51352_ (_43962_, _43000_, _38549_);
  and _51353_ (_43963_, _43962_, _41806_);
  and _51354_ (_38995_, _43963_, _43961_);
  or _51355_ (_43964_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _51356_ (_43965_, _43000_, _38554_);
  and _51357_ (_43966_, _43965_, _41806_);
  and _51358_ (_38996_, _43966_, _43964_);
  or _51359_ (_43967_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _51360_ (_43968_, _43000_, _38539_);
  and _51361_ (_43969_, _43968_, _41806_);
  and _51362_ (_38997_, _43969_, _43967_);
  or _51363_ (_43970_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _51364_ (_43971_, _43000_, _38560_);
  and _51365_ (_43972_, _43971_, _41806_);
  and _51366_ (_38998_, _43972_, _43970_);
  or _51367_ (_43973_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _51368_ (_43974_, _43000_, _38535_);
  and _51369_ (_43975_, _43974_, _41806_);
  and _51370_ (_39000_, _43975_, _43973_);
  or _51371_ (_43976_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _51372_ (_43977_, _43000_, _38566_);
  and _51373_ (_43978_, _43977_, _41806_);
  and _51374_ (_39001_, _43978_, _43976_);
  or _51375_ (_43979_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _51376_ (_43980_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _41806_);
  or _51377_ (_43981_, _43980_, _00000_);
  and _51378_ (_39005_, _43981_, _43979_);
  or _51379_ (_43982_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _51380_ (_43983_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _41806_);
  or _51381_ (_43984_, _43983_, _00000_);
  and _51382_ (_39006_, _43984_, _43982_);
  or _51383_ (_43985_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _51384_ (_43986_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _41806_);
  or _51385_ (_43987_, _43986_, _00000_);
  and _51386_ (_39007_, _43987_, _43985_);
  or _51387_ (_43988_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _51388_ (_43989_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _41806_);
  or _51389_ (_43990_, _43989_, _00000_);
  and _51390_ (_39008_, _43990_, _43988_);
  or _51391_ (_43991_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _51392_ (_43992_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _41806_);
  or _51393_ (_43993_, _43992_, _00000_);
  and _51394_ (_39009_, _43993_, _43991_);
  or _51395_ (_43994_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _51396_ (_43995_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _41806_);
  or _51397_ (_43996_, _43995_, _00000_);
  and _51398_ (_39010_, _43996_, _43994_);
  or _51399_ (_43997_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _51400_ (_43998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _41806_);
  or _51401_ (_43999_, _43998_, _00000_);
  and _51402_ (_39011_, _43999_, _43997_);
  or _51403_ (_44000_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _51404_ (_44001_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _41806_);
  or _51405_ (_44002_, _44001_, _00000_);
  and _51406_ (_39012_, _44002_, _44000_);
  or _51407_ (_44003_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _51408_ (_44004_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _41806_);
  or _51409_ (_44005_, _44004_, _00000_);
  and _51410_ (_39013_, _44005_, _44003_);
  or _51411_ (_44006_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _51412_ (_44007_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _41806_);
  or _51413_ (_44008_, _44007_, _00000_);
  and _51414_ (_39014_, _44008_, _44006_);
  or _51415_ (_44009_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _51416_ (_44010_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _41806_);
  or _51417_ (_44011_, _44010_, _00000_);
  and _51418_ (_39015_, _44011_, _44009_);
  or _51419_ (_44012_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _51420_ (_44013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _41806_);
  or _51421_ (_44014_, _44013_, _00000_);
  and _51422_ (_39016_, _44014_, _44012_);
  or _51423_ (_44015_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _51424_ (_44016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _41806_);
  or _51425_ (_44017_, _44016_, _00000_);
  and _51426_ (_39017_, _44017_, _44015_);
  or _51427_ (_44018_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _51428_ (_44019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _41806_);
  or _51429_ (_44020_, _44019_, _00000_);
  and _51430_ (_39018_, _44020_, _44018_);
  or _51431_ (_44021_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _51432_ (_44022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _41806_);
  or _51433_ (_44023_, _44022_, _00000_);
  and _51434_ (_39019_, _44023_, _44021_);
  and _51435_ (_44024_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _51436_ (_44025_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _51437_ (_44026_, _44025_, _44024_);
  and _51438_ (_39197_, _44026_, _41806_);
  and _51439_ (_44027_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _51440_ (_44028_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or _51441_ (_44029_, _44028_, _44027_);
  and _51442_ (_39198_, _44029_, _41806_);
  and _51443_ (_44030_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _51444_ (_44031_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _51445_ (_44032_, _44031_, _44030_);
  and _51446_ (_39199_, _44032_, _41806_);
  and _51447_ (_44033_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _51448_ (_44034_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _51449_ (_44035_, _44034_, _43896_);
  or _51450_ (_44036_, _44035_, _44033_);
  and _51451_ (_39200_, _44036_, _41806_);
  and _51452_ (_44037_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _51453_ (_44038_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _51454_ (_44039_, _44038_, _44037_);
  and _51455_ (_39201_, _44039_, _41806_);
  and _51456_ (_44040_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _51457_ (_44041_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or _51458_ (_44042_, _44041_, _44040_);
  and _51459_ (_39202_, _44042_, _41806_);
  and _51460_ (_44043_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _51461_ (_44044_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _51462_ (_44045_, _44044_, _43896_);
  or _51463_ (_44046_, _44045_, _44043_);
  and _51464_ (_39204_, _44046_, _41806_);
  and _51465_ (_44047_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _51466_ (_44048_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _51467_ (_44049_, _44048_, _44047_);
  and _51468_ (_39205_, _44049_, _41806_);
  and _51469_ (_44050_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _51470_ (_44051_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _51471_ (_44052_, _44051_, _44050_);
  and _51472_ (_39206_, _44052_, _41806_);
  and _51473_ (_44053_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _51474_ (_44054_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _51475_ (_44055_, _44054_, _44053_);
  and _51476_ (_39207_, _44055_, _41806_);
  and _51477_ (_44056_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _51478_ (_44057_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _51479_ (_44058_, _44057_, _44056_);
  and _51480_ (_39208_, _44058_, _41806_);
  and _51481_ (_44059_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _51482_ (_44060_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _51483_ (_00008_, _44060_, _44059_);
  and _51484_ (_39209_, _00008_, _41806_);
  and _51485_ (_00009_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _51486_ (_00010_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _51487_ (_00011_, _00010_, _00009_);
  and _51488_ (_39210_, _00011_, _41806_);
  and _51489_ (_00012_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _51490_ (_00013_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _51491_ (_00014_, _00013_, _00012_);
  and _51492_ (_39211_, _00014_, _41806_);
  and _51493_ (_00015_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _51494_ (_00016_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _51495_ (_00017_, _00016_, _00015_);
  and _51496_ (_39212_, _00017_, _41806_);
  and _51497_ (_00018_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _51498_ (_00019_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _51499_ (_00020_, _00019_, _00018_);
  and _51500_ (_39213_, _00020_, _41806_);
  and _51501_ (_00021_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _51502_ (_00022_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _51503_ (_00023_, _00022_, _00021_);
  and _51504_ (_39215_, _00023_, _41806_);
  and _51505_ (_00024_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _51506_ (_00025_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _51507_ (_00026_, _00025_, _00024_);
  and _51508_ (_39216_, _00026_, _41806_);
  and _51509_ (_00027_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _51510_ (_00028_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _51511_ (_00029_, _00028_, _00027_);
  and _51512_ (_39217_, _00029_, _41806_);
  and _51513_ (_00030_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _51514_ (_00031_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _51515_ (_00032_, _00031_, _00030_);
  and _51516_ (_39218_, _00032_, _41806_);
  and _51517_ (_00033_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _51518_ (_00034_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _51519_ (_00035_, _00034_, _00033_);
  and _51520_ (_39219_, _00035_, _41806_);
  and _51521_ (_00036_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _51522_ (_00037_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _51523_ (_00038_, _00037_, _00036_);
  and _51524_ (_39220_, _00038_, _41806_);
  and _51525_ (_00039_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _51526_ (_00040_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _51527_ (_00041_, _00040_, _00039_);
  and _51528_ (_39221_, _00041_, _41806_);
  and _51529_ (_00042_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _51530_ (_00043_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _51531_ (_00044_, _00043_, _00042_);
  and _51532_ (_39222_, _00044_, _41806_);
  and _51533_ (_00045_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _51534_ (_00046_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _51535_ (_00047_, _00046_, _00045_);
  and _51536_ (_39223_, _00047_, _41806_);
  and _51537_ (_00048_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _51538_ (_00049_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _51539_ (_00050_, _00049_, _00048_);
  and _51540_ (_39224_, _00050_, _41806_);
  and _51541_ (_00051_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _51542_ (_00052_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _51543_ (_00053_, _00052_, _00051_);
  and _51544_ (_39226_, _00053_, _41806_);
  and _51545_ (_00054_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _51546_ (_00055_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _51547_ (_00056_, _00055_, _00054_);
  and _51548_ (_39227_, _00056_, _41806_);
  and _51549_ (_00057_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _51550_ (_00058_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _51551_ (_00059_, _00058_, _00057_);
  and _51552_ (_39228_, _00059_, _41806_);
  and _51553_ (_00060_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _51554_ (_00061_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _51555_ (_00062_, _00061_, _00060_);
  and _51556_ (_39229_, _00062_, _41806_);
  and _51557_ (_00063_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _51558_ (_00064_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _51559_ (_00065_, _00064_, _00063_);
  and _51560_ (_39230_, _00065_, _41806_);
  nor _51561_ (_39231_, _36409_, rst);
  nor _51562_ (_39232_, _35056_, rst);
  nor _51563_ (_39233_, _35286_, rst);
  nor _51564_ (_39234_, _40279_, rst);
  nor _51565_ (_39236_, _40408_, rst);
  nor _51566_ (_39237_, _40564_, rst);
  nor _51567_ (_39238_, _40492_, rst);
  nor _51568_ (_39239_, _40370_, rst);
  and _51569_ (_39240_, _40540_, _41806_);
  nor _51570_ (_39242_, _40442_, rst);
  nor _51571_ (_39243_, _40639_, rst);
  and _51572_ (_39259_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _41806_);
  and _51573_ (_39260_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _41806_);
  and _51574_ (_39261_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _41806_);
  and _51575_ (_39263_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _41806_);
  and _51576_ (_39264_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _41806_);
  and _51577_ (_39265_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _41806_);
  and _51578_ (_39266_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _41806_);
  or _51579_ (_00066_, _43132_, _43111_);
  and _51580_ (_00067_, _00066_, _29242_);
  and _51581_ (_00068_, _43266_, _40397_);
  and _51582_ (_00069_, _43114_, _43194_);
  or _51583_ (_00070_, _00069_, _00068_);
  and _51584_ (_00071_, _37624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _51585_ (_00072_, _00071_, _00070_);
  or _51586_ (_00073_, _00072_, _00067_);
  nor _51587_ (_00074_, _43198_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _51588_ (_00075_, _00074_, _43199_);
  nand _51589_ (_00076_, _00075_, _43261_);
  nand _51590_ (_00077_, _00076_, _43108_);
  or _51591_ (_00078_, _00077_, _00073_);
  or _51592_ (_00079_, _43108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _51593_ (_00080_, _00079_, _41806_);
  and _51594_ (_39267_, _00080_, _00078_);
  not _51595_ (_00081_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _51596_ (_00082_, _43109_, _00081_);
  and _51597_ (_00083_, _43114_, _43187_);
  and _51598_ (_00084_, _43266_, _40607_);
  or _51599_ (_00085_, _00084_, _00083_);
  or _51600_ (_00086_, _43202_, _43199_);
  not _51601_ (_00087_, _43261_);
  nor _51602_ (_00088_, _00087_, _43203_);
  and _51603_ (_00089_, _00088_, _00086_);
  or _51604_ (_00090_, _00089_, _00085_);
  and _51605_ (_00091_, _00066_, _29904_);
  or _51606_ (_00092_, _00091_, _00090_);
  and _51607_ (_00093_, _00092_, _43108_);
  or _51608_ (_00094_, _00093_, _00082_);
  and _51609_ (_39268_, _00094_, _41806_);
  and _51610_ (_00095_, _00066_, _30578_);
  and _51611_ (_00096_, _43266_, _40480_);
  and _51612_ (_00097_, _43114_, _43181_);
  or _51613_ (_00098_, _00097_, _00096_);
  or _51614_ (_00099_, _43209_, _43206_);
  nor _51615_ (_00100_, _00087_, _43210_);
  and _51616_ (_00101_, _00100_, _00099_);
  or _51617_ (_00102_, _00101_, _00098_);
  and _51618_ (_00103_, _37624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _51619_ (_00104_, _00103_, _00102_);
  nand _51620_ (_00105_, _00104_, _43108_);
  or _51621_ (_00106_, _00105_, _00095_);
  not _51622_ (_00107_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _51623_ (_00108_, _43309_, _00107_);
  and _51624_ (_00109_, _43309_, _00107_);
  nor _51625_ (_00110_, _00109_, _00108_);
  or _51626_ (_00111_, _00110_, _43108_);
  and _51627_ (_00112_, _00111_, _41806_);
  and _51628_ (_39269_, _00112_, _00106_);
  and _51629_ (_00113_, _00066_, _31349_);
  and _51630_ (_00114_, _43266_, _40357_);
  and _51631_ (_00115_, _43114_, _43174_);
  or _51632_ (_00116_, _00115_, _00114_);
  and _51633_ (_00117_, _37624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _51634_ (_00118_, _00117_, _00116_);
  or _51635_ (_00119_, _43179_, _43178_);
  or _51636_ (_00120_, _00119_, _43211_);
  nand _51637_ (_00121_, _00119_, _43211_);
  and _51638_ (_00122_, _00121_, _00120_);
  and _51639_ (_00123_, _00122_, _43261_);
  nor _51640_ (_00124_, _00123_, _00118_);
  nand _51641_ (_00125_, _00124_, _43108_);
  or _51642_ (_00126_, _00125_, _00113_);
  and _51643_ (_00127_, _00108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _51644_ (_00128_, _00108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _51645_ (_00129_, _00128_, _00127_);
  or _51646_ (_00130_, _00129_, _43108_);
  and _51647_ (_00131_, _00130_, _41806_);
  and _51648_ (_39270_, _00131_, _00126_);
  and _51649_ (_00132_, _00066_, _32055_);
  and _51650_ (_00133_, _43266_, _40528_);
  and _51651_ (_00134_, _43114_, _43167_);
  and _51652_ (_00135_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _51653_ (_00136_, _00135_, _00134_);
  or _51654_ (_00137_, _00136_, _00133_);
  or _51655_ (_00138_, _00137_, _00132_);
  or _51656_ (_00139_, _43216_, _43213_);
  and _51657_ (_00140_, _00139_, _43217_);
  nand _51658_ (_00141_, _00140_, _43261_);
  nand _51659_ (_00142_, _00141_, _43108_);
  or _51660_ (_00143_, _00142_, _00138_);
  and _51661_ (_00144_, _43294_, _43311_);
  nor _51662_ (_00145_, _00127_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _51663_ (_00146_, _00145_, _00144_);
  or _51664_ (_00147_, _00146_, _43108_);
  and _51665_ (_00148_, _00147_, _41806_);
  and _51666_ (_39271_, _00148_, _00143_);
  and _51667_ (_00149_, _00066_, _32864_);
  and _51668_ (_00150_, _43266_, _40459_);
  and _51669_ (_00151_, _43114_, _43160_);
  and _51670_ (_00152_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _51671_ (_00153_, _00152_, _00151_);
  or _51672_ (_00154_, _00153_, _00150_);
  or _51673_ (_00155_, _00154_, _00149_);
  or _51674_ (_00156_, _43165_, _43166_);
  or _51675_ (_00157_, _00156_, _43218_);
  nand _51676_ (_00158_, _00156_, _43218_);
  and _51677_ (_00159_, _00158_, _00157_);
  nand _51678_ (_00160_, _00159_, _43261_);
  nand _51679_ (_00161_, _00160_, _43108_);
  or _51680_ (_00162_, _00161_, _00155_);
  and _51681_ (_00163_, _43296_, _43311_);
  nor _51682_ (_00164_, _00144_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _51683_ (_00165_, _00164_, _00163_);
  or _51684_ (_00166_, _00165_, _43108_);
  and _51685_ (_00167_, _00166_, _41806_);
  and _51686_ (_39272_, _00167_, _00162_);
  not _51687_ (_00168_, _43108_);
  nor _51688_ (_00169_, _43221_, _43159_);
  nor _51689_ (_00170_, _00169_, _43222_);
  and _51690_ (_00171_, _00170_, _43261_);
  and _51691_ (_00172_, _00066_, _33609_);
  and _51692_ (_00173_, _43266_, _40683_);
  and _51693_ (_00174_, _43114_, _43152_);
  and _51694_ (_00175_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _51695_ (_00176_, _00175_, _00174_);
  or _51696_ (_00177_, _00176_, _00173_);
  or _51697_ (_00178_, _00177_, _00172_);
  or _51698_ (_00179_, _00178_, _00171_);
  or _51699_ (_00180_, _00179_, _00168_);
  and _51700_ (_00181_, _00163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _51701_ (_00182_, _00163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _51702_ (_00183_, _00182_, _00181_);
  or _51703_ (_00184_, _00183_, _43108_);
  and _51704_ (_00185_, _00184_, _41806_);
  and _51705_ (_39274_, _00185_, _00180_);
  and _51706_ (_00186_, _00066_, _28022_);
  and _51707_ (_00187_, _43266_, _40322_);
  and _51708_ (_00188_, _43114_, _43138_);
  and _51709_ (_00189_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _51710_ (_00190_, _00189_, _00188_);
  or _51711_ (_00191_, _00190_, _00187_);
  or _51712_ (_00192_, _43225_, _43150_);
  and _51713_ (_00193_, _00192_, _43226_);
  and _51714_ (_00194_, _00193_, _43261_);
  or _51715_ (_00195_, _00194_, _00191_);
  or _51716_ (_00196_, _00195_, _00186_);
  or _51717_ (_00197_, _00196_, _00168_);
  and _51718_ (_00198_, _00181_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _51719_ (_00199_, _00181_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _51720_ (_00200_, _00199_, _00198_);
  or _51721_ (_00201_, _00200_, _43108_);
  and _51722_ (_00202_, _00201_, _41806_);
  and _51723_ (_39275_, _00202_, _00197_);
  nor _51724_ (_00203_, _37635_, _29231_);
  nor _51725_ (_00204_, _43112_, _38617_);
  and _51726_ (_00205_, _43114_, _40397_);
  and _51727_ (_00206_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _51728_ (_00207_, _00206_, _00205_);
  and _51729_ (_00208_, _43266_, _42329_);
  nor _51730_ (_00209_, _43228_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _51731_ (_00210_, _43228_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _51732_ (_00211_, _00210_, _00209_);
  or _51733_ (_00212_, _00211_, _43238_);
  nand _51734_ (_00213_, _00211_, _43238_);
  and _51735_ (_00214_, _00213_, _43261_);
  and _51736_ (_00215_, _00214_, _00212_);
  or _51737_ (_00216_, _00215_, _00208_);
  or _51738_ (_00217_, _00216_, _00207_);
  or _51739_ (_00218_, _00217_, _00204_);
  or _51740_ (_00219_, _00218_, _00203_);
  or _51741_ (_00220_, _00219_, _00168_);
  and _51742_ (_00221_, _00198_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _51743_ (_00222_, _00198_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _51744_ (_00223_, _00222_, _00221_);
  or _51745_ (_00224_, _00223_, _43108_);
  and _51746_ (_00225_, _00224_, _41806_);
  and _51747_ (_39276_, _00225_, _00220_);
  nor _51748_ (_00226_, _43112_, _38645_);
  and _51749_ (_00227_, _43266_, _42353_);
  and _51750_ (_00228_, _43114_, _40607_);
  and _51751_ (_00229_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _51752_ (_00230_, _00229_, _00228_);
  or _51753_ (_00231_, _00230_, _00227_);
  or _51754_ (_00232_, _00231_, _00226_);
  nor _51755_ (_00233_, _37635_, _29893_);
  or _51756_ (_00234_, _00233_, _00232_);
  and _51757_ (_00235_, _43240_, _43146_);
  and _51758_ (_00236_, _43229_, _43238_);
  nor _51759_ (_00237_, _00236_, _00235_);
  nor _51760_ (_00238_, _00237_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _51761_ (_00239_, _00237_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _51762_ (_00240_, _00239_, _00238_);
  and _51763_ (_00241_, _00240_, _43261_);
  or _51764_ (_00242_, _00241_, _00168_);
  or _51765_ (_00243_, _00242_, _00234_);
  and _51766_ (_00244_, _43301_, _43311_);
  nor _51767_ (_00245_, _00221_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _51768_ (_00246_, _00245_, _00244_);
  or _51769_ (_00247_, _00246_, _43108_);
  and _51770_ (_00248_, _00247_, _41806_);
  and _51771_ (_39277_, _00248_, _00243_);
  or _51772_ (_00249_, _37635_, _30567_);
  or _51773_ (_00250_, _43112_, _38673_);
  nand _51774_ (_00251_, _43114_, _40480_);
  nand _51775_ (_00252_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _51776_ (_00253_, _00252_, _00251_);
  and _51777_ (_00254_, _00253_, _00250_);
  nand _51778_ (_00255_, _43266_, _42333_);
  and _51779_ (_00256_, _43241_, _43146_);
  and _51780_ (_00257_, _43230_, _43238_);
  nor _51781_ (_00258_, _00257_, _00256_);
  nor _51782_ (_00259_, _00258_, _38554_);
  and _51783_ (_00260_, _00258_, _38554_);
  or _51784_ (_00261_, _00260_, _00087_);
  or _51785_ (_00262_, _00261_, _00259_);
  and _51786_ (_00263_, _00262_, _00255_);
  and _51787_ (_00264_, _00263_, _00254_);
  and _51788_ (_00265_, _00264_, _00249_);
  nand _51789_ (_00266_, _00265_, _43108_);
  and _51790_ (_00267_, _00244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _51791_ (_00268_, _00244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _51792_ (_00269_, _00268_, _00267_);
  or _51793_ (_00270_, _00269_, _43108_);
  and _51794_ (_00271_, _00270_, _41806_);
  and _51795_ (_39278_, _00271_, _00266_);
  nor _51796_ (_00272_, _43278_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _51797_ (_00273_, _00272_, _43279_);
  and _51798_ (_00274_, _00273_, _43266_);
  and _51799_ (_00275_, _43232_, _43238_);
  and _51800_ (_00276_, _43243_, _43146_);
  nor _51801_ (_00277_, _00276_, _00275_);
  or _51802_ (_00278_, _00277_, _38539_);
  nand _51803_ (_00279_, _00277_, _38539_);
  and _51804_ (_00280_, _00279_, _43261_);
  and _51805_ (_00281_, _00280_, _00278_);
  nor _51806_ (_00282_, _37635_, _31338_);
  nor _51807_ (_00283_, _43112_, _38702_);
  and _51808_ (_00284_, _43114_, _40357_);
  and _51809_ (_00285_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _51810_ (_00286_, _00285_, _00284_);
  or _51811_ (_00287_, _00286_, _00283_);
  or _51812_ (_00288_, _00287_, _00282_);
  or _51813_ (_00289_, _00288_, _00281_);
  or _51814_ (_00290_, _00289_, _00274_);
  or _51815_ (_00291_, _00290_, _00168_);
  and _51816_ (_00292_, _00267_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _51817_ (_00293_, _00267_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _51818_ (_00294_, _00293_, _00292_);
  or _51819_ (_00295_, _00294_, _43108_);
  and _51820_ (_00296_, _00295_, _41806_);
  and _51821_ (_39279_, _00296_, _00291_);
  and _51822_ (_00297_, _43233_, _43238_);
  and _51823_ (_00298_, _43244_, _43146_);
  nor _51824_ (_00299_, _00298_, _00297_);
  or _51825_ (_00300_, _00299_, _38560_);
  nand _51826_ (_00301_, _00299_, _38560_);
  and _51827_ (_00302_, _00301_, _43261_);
  and _51828_ (_00303_, _00302_, _00300_);
  nor _51829_ (_00304_, _43279_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _51830_ (_00305_, _00304_, _43280_);
  and _51831_ (_00306_, _00305_, _43266_);
  nor _51832_ (_00307_, _37635_, _32044_);
  nor _51833_ (_00308_, _43112_, _38731_);
  and _51834_ (_00309_, _43114_, _40528_);
  and _51835_ (_00310_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _51836_ (_00311_, _00310_, _00309_);
  or _51837_ (_00312_, _00311_, _00308_);
  or _51838_ (_00313_, _00312_, _00307_);
  or _51839_ (_00314_, _00313_, _00306_);
  or _51840_ (_00315_, _00314_, _00303_);
  or _51841_ (_00316_, _00315_, _00168_);
  and _51842_ (_00317_, _00292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _51843_ (_00318_, _00292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _51844_ (_00319_, _00318_, _00317_);
  or _51845_ (_00320_, _00319_, _43108_);
  and _51846_ (_00321_, _00320_, _41806_);
  and _51847_ (_39280_, _00321_, _00316_);
  nor _51848_ (_00322_, _37635_, _32853_);
  nor _51849_ (_00323_, _43112_, _38760_);
  and _51850_ (_00324_, _43114_, _40459_);
  and _51851_ (_00325_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _51852_ (_00326_, _00325_, _00324_);
  or _51853_ (_00327_, _00326_, _00323_);
  or _51854_ (_00328_, _00327_, _00322_);
  and _51855_ (_00329_, _00297_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _51856_ (_00330_, _00298_, _38560_);
  nor _51857_ (_00331_, _00330_, _00329_);
  nand _51858_ (_00332_, _00331_, _38535_);
  or _51859_ (_00333_, _00331_, _38535_);
  and _51860_ (_00334_, _00333_, _00332_);
  and _51861_ (_00335_, _00334_, _43261_);
  or _51862_ (_00336_, _00335_, _00328_);
  nor _51863_ (_00337_, _43280_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _51864_ (_00338_, _00337_, _43281_);
  nand _51865_ (_00339_, _00338_, _43266_);
  nand _51866_ (_00340_, _00339_, _43108_);
  or _51867_ (_00341_, _00340_, _00336_);
  or _51868_ (_00342_, _00317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _51869_ (_00343_, _00317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _51870_ (_00344_, _00343_, _00342_);
  or _51871_ (_00345_, _00344_, _43108_);
  and _51872_ (_00346_, _00345_, _41806_);
  and _51873_ (_39281_, _00346_, _00341_);
  or _51874_ (_00347_, _43281_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _51875_ (_00348_, _00347_, _43282_);
  nand _51876_ (_00349_, _00348_, _43266_);
  or _51877_ (_00350_, _37635_, _33598_);
  or _51878_ (_00351_, _43112_, _38787_);
  nand _51879_ (_00352_, _43114_, _40683_);
  nand _51880_ (_00353_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _51881_ (_00354_, _00353_, _00352_);
  and _51882_ (_00355_, _00354_, _00351_);
  and _51883_ (_00356_, _00355_, _00350_);
  or _51884_ (_00357_, _43249_, _38566_);
  nand _51885_ (_00358_, _43249_, _38566_);
  and _51886_ (_00359_, _00358_, _00357_);
  or _51887_ (_00360_, _00359_, _00087_);
  and _51888_ (_00361_, _00360_, _00356_);
  and _51889_ (_00362_, _00361_, _00349_);
  nand _51890_ (_00363_, _00362_, _43108_);
  or _51891_ (_00364_, _43313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _51892_ (_00365_, _00364_, _43314_);
  or _51893_ (_00366_, _00365_, _43108_);
  and _51894_ (_00367_, _00366_, _41806_);
  and _51895_ (_39282_, _00367_, _00363_);
  and _51896_ (_00368_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _51897_ (_00369_, _43777_, _43774_);
  nor _51898_ (_00370_, _00369_, _43778_);
  or _51899_ (_00371_, _00370_, _43328_);
  or _51900_ (_00372_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _51901_ (_00373_, _00372_, _43821_);
  and _51902_ (_00374_, _00373_, _00371_);
  or _51903_ (_39283_, _00374_, _00368_);
  nor _51904_ (_00375_, _43781_, _43778_);
  nor _51905_ (_00376_, _00375_, _43782_);
  or _51906_ (_00377_, _00376_, _43328_);
  or _51907_ (_00378_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _51908_ (_00379_, _00378_, _43821_);
  and _51909_ (_00380_, _00379_, _00377_);
  and _51910_ (_00381_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _51911_ (_39285_, _00381_, _00380_);
  and _51912_ (_00382_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _51913_ (_00383_, _43787_, _43785_);
  nor _51914_ (_00384_, _00383_, _43789_);
  or _51915_ (_00385_, _00384_, _43328_);
  or _51916_ (_00386_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _51917_ (_00387_, _00386_, _43821_);
  and _51918_ (_00388_, _00387_, _00385_);
  or _51919_ (_39286_, _00388_, _00382_);
  and _51920_ (_00389_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _51921_ (_00390_, _43789_, _43441_);
  nor _51922_ (_00391_, _00390_, _43790_);
  or _51923_ (_00392_, _00391_, _43328_);
  or _51924_ (_00393_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _51925_ (_00394_, _00393_, _43821_);
  and _51926_ (_00395_, _00394_, _00392_);
  or _51927_ (_39287_, _00395_, _00389_);
  and _51928_ (_00396_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _51929_ (_00397_, _43794_, _43790_);
  nor _51930_ (_00398_, _00397_, _43795_);
  or _51931_ (_00399_, _00398_, _43328_);
  or _51932_ (_00400_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _51933_ (_00401_, _00400_, _43821_);
  and _51934_ (_00402_, _00401_, _00399_);
  or _51935_ (_39288_, _00402_, _00396_);
  and _51936_ (_00403_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _51937_ (_00404_, _43795_, _43434_);
  nor _51938_ (_00405_, _00404_, _43797_);
  or _51939_ (_00406_, _00405_, _43328_);
  or _51940_ (_00407_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _51941_ (_00408_, _00407_, _43821_);
  and _51942_ (_00409_, _00408_, _00406_);
  or _51943_ (_39289_, _00409_, _00403_);
  nor _51944_ (_00410_, _43797_, _43428_);
  nor _51945_ (_00411_, _00410_, _43798_);
  or _51946_ (_00412_, _00411_, _43328_);
  or _51947_ (_00413_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _51948_ (_00414_, _00413_, _43821_);
  and _51949_ (_00415_, _00414_, _00412_);
  and _51950_ (_00416_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _51951_ (_39290_, _00416_, _00415_);
  and _51952_ (_00417_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _51953_ (_00418_, _43798_, _43424_);
  nor _51954_ (_00419_, _00418_, _43799_);
  or _51955_ (_00420_, _00419_, _43328_);
  or _51956_ (_00421_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _51957_ (_00422_, _00421_, _43821_);
  and _51958_ (_00423_, _00422_, _00420_);
  or _51959_ (_39291_, _00423_, _00417_);
  nor _51960_ (_00424_, _43802_, _43799_);
  nor _51961_ (_00425_, _00424_, _43803_);
  or _51962_ (_00426_, _00425_, _43328_);
  or _51963_ (_00427_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _51964_ (_00428_, _00427_, _43821_);
  and _51965_ (_00429_, _00428_, _00426_);
  and _51966_ (_00430_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _51967_ (_39292_, _00430_, _00429_);
  nor _51968_ (_00431_, _43803_, _43418_);
  nor _51969_ (_00432_, _00431_, _43805_);
  or _51970_ (_00433_, _00432_, _43328_);
  or _51971_ (_00434_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _51972_ (_00435_, _00434_, _43821_);
  and _51973_ (_00436_, _00435_, _00433_);
  and _51974_ (_00437_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _51975_ (_39293_, _00437_, _00436_);
  nor _51976_ (_00438_, _43805_, _43409_);
  nor _51977_ (_00439_, _00438_, _43806_);
  or _51978_ (_00440_, _00439_, _43328_);
  or _51979_ (_00441_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _51980_ (_00442_, _00441_, _43821_);
  and _51981_ (_00443_, _00442_, _00440_);
  and _51982_ (_00444_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _51983_ (_39294_, _00444_, _00443_);
  nor _51984_ (_00445_, _43806_, _43406_);
  nor _51985_ (_00446_, _00445_, _43807_);
  or _51986_ (_00447_, _00446_, _43328_);
  or _51987_ (_00448_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _51988_ (_00449_, _00448_, _43821_);
  and _51989_ (_00450_, _00449_, _00447_);
  and _51990_ (_00451_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _51991_ (_39296_, _00451_, _00450_);
  nor _51992_ (_00452_, _43807_, _43399_);
  nor _51993_ (_00453_, _00452_, _43809_);
  or _51994_ (_00454_, _00453_, _43328_);
  or _51995_ (_00455_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _51996_ (_00456_, _00455_, _43821_);
  and _51997_ (_00457_, _00456_, _00454_);
  and _51998_ (_00458_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _51999_ (_39297_, _00458_, _00457_);
  nor _52000_ (_00459_, _43809_, _43393_);
  nor _52001_ (_00460_, _00459_, _43810_);
  or _52002_ (_00461_, _00460_, _43328_);
  or _52003_ (_00462_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _52004_ (_00463_, _00462_, _43821_);
  and _52005_ (_00464_, _00463_, _00461_);
  and _52006_ (_00465_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _52007_ (_39298_, _00465_, _00464_);
  nor _52008_ (_00466_, _43810_, _43387_);
  nor _52009_ (_00467_, _00466_, _43811_);
  or _52010_ (_00468_, _00467_, _43328_);
  or _52011_ (_00469_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _52012_ (_00470_, _00469_, _43821_);
  and _52013_ (_00471_, _00470_, _00468_);
  and _52014_ (_00472_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _52015_ (_39299_, _00472_, _00471_);
  and _52016_ (_00473_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _52017_ (_00474_, _00473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _52018_ (_39300_, _00474_, _41806_);
  and _52019_ (_00475_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _52020_ (_00476_, _00475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _52021_ (_39301_, _00476_, _41806_);
  and _52022_ (_00477_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _52023_ (_00478_, _00477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _52024_ (_39302_, _00478_, _41806_);
  and _52025_ (_00479_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _52026_ (_00480_, _00479_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _52027_ (_39303_, _00480_, _41806_);
  and _52028_ (_00481_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _52029_ (_00482_, _00481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _52030_ (_39304_, _00482_, _41806_);
  and _52031_ (_00483_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _52032_ (_00484_, _00483_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _52033_ (_39305_, _00484_, _41806_);
  and _52034_ (_00485_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _52035_ (_00486_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _52036_ (_39307_, _00486_, _41806_);
  nor _52037_ (_00487_, _43773_, _40305_);
  nand _52038_ (_00488_, _00487_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _52039_ (_00489_, _00487_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _52040_ (_00490_, _00489_, _43821_);
  and _52041_ (_39308_, _00490_, _00488_);
  nor _52042_ (_00491_, _43850_, _43848_);
  nor _52043_ (_00492_, _00491_, _43851_);
  or _52044_ (_00493_, _00492_, _40305_);
  or _52045_ (_00494_, _33860_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _52046_ (_00495_, _00494_, _43821_);
  and _52047_ (_39309_, _00495_, _00493_);
  and _52048_ (_00496_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _52049_ (_00497_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _52050_ (_00498_, _00497_, _38935_);
  or _52051_ (_39324_, _00498_, _00496_);
  and _52052_ (_00499_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _52053_ (_00500_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _52054_ (_00501_, _00500_, _38935_);
  or _52055_ (_39325_, _00501_, _00499_);
  and _52056_ (_00502_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _52057_ (_00503_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _52058_ (_00504_, _00503_, _38935_);
  or _52059_ (_39326_, _00504_, _00502_);
  and _52060_ (_00505_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _52061_ (_00506_, _44034_, _38935_);
  or _52062_ (_39328_, _00506_, _00505_);
  and _52063_ (_00507_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _52064_ (_00508_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _52065_ (_00509_, _00508_, _38935_);
  or _52066_ (_39329_, _00509_, _00507_);
  and _52067_ (_00510_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _52068_ (_00511_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _52069_ (_00512_, _00511_, _38935_);
  or _52070_ (_39330_, _00512_, _00510_);
  and _52071_ (_00513_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _52072_ (_00514_, _44044_, _38935_);
  or _52073_ (_39331_, _00514_, _00513_);
  and _52074_ (_39332_, _43882_, _41806_);
  nor _52075_ (_39333_, _43892_, rst);
  and _52076_ (_39334_, _43888_, _41806_);
  and _52077_ (_00515_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _52078_ (_00516_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or _52079_ (_00517_, _00516_, _00515_);
  and _52080_ (_39335_, _00517_, _41806_);
  and _52081_ (_00518_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _52082_ (_00519_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or _52083_ (_00520_, _00519_, _00518_);
  and _52084_ (_39336_, _00520_, _41806_);
  and _52085_ (_00521_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _52086_ (_00522_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or _52087_ (_00523_, _00522_, _00521_);
  and _52088_ (_39337_, _00523_, _41806_);
  and _52089_ (_00524_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _52090_ (_00525_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or _52091_ (_00526_, _00525_, _00524_);
  and _52092_ (_39339_, _00526_, _41806_);
  and _52093_ (_00527_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _52094_ (_00528_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or _52095_ (_00529_, _00528_, _00527_);
  and _52096_ (_39340_, _00529_, _41806_);
  and _52097_ (_00530_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _52098_ (_00531_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or _52099_ (_00532_, _00531_, _00530_);
  and _52100_ (_39341_, _00532_, _41806_);
  and _52101_ (_00533_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _52102_ (_00534_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or _52103_ (_00535_, _00534_, _00533_);
  and _52104_ (_39342_, _00535_, _41806_);
  and _52105_ (_00536_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _52106_ (_00537_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or _52107_ (_00538_, _00537_, _00536_);
  and _52108_ (_39343_, _00538_, _41806_);
  and _52109_ (_00539_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _52110_ (_00540_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _52111_ (_00541_, _00540_, _00539_);
  and _52112_ (_39344_, _00541_, _41806_);
  and _52113_ (_00542_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _52114_ (_00543_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _52115_ (_00544_, _00543_, _00542_);
  and _52116_ (_39345_, _00544_, _41806_);
  and _52117_ (_00545_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _52118_ (_00546_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _52119_ (_00547_, _00546_, _00545_);
  and _52120_ (_39346_, _00547_, _41806_);
  and _52121_ (_00548_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _52122_ (_00549_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _52123_ (_00550_, _00549_, _00548_);
  and _52124_ (_39347_, _00550_, _41806_);
  and _52125_ (_00551_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _52126_ (_00552_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _52127_ (_00553_, _00552_, _00551_);
  and _52128_ (_39348_, _00553_, _41806_);
  and _52129_ (_00554_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _52130_ (_00555_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _52131_ (_00556_, _00555_, _00554_);
  and _52132_ (_39350_, _00556_, _41806_);
  and _52133_ (_00557_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _52134_ (_00558_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _52135_ (_00559_, _00558_, _00557_);
  and _52136_ (_39351_, _00559_, _41806_);
  and _52137_ (_00560_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _52138_ (_00561_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _52139_ (_00562_, _00561_, _00560_);
  and _52140_ (_39352_, _00562_, _41806_);
  and _52141_ (_00563_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _52142_ (_00564_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _52143_ (_00565_, _00564_, _00563_);
  and _52144_ (_39353_, _00565_, _41806_);
  and _52145_ (_00566_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _52146_ (_00567_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _52147_ (_00568_, _00567_, _00566_);
  and _52148_ (_39354_, _00568_, _41806_);
  and _52149_ (_00569_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _52150_ (_00570_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _52151_ (_00571_, _00570_, _00569_);
  and _52152_ (_39355_, _00571_, _41806_);
  and _52153_ (_00572_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _52154_ (_00573_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _52155_ (_00574_, _00573_, _00572_);
  and _52156_ (_39356_, _00574_, _41806_);
  and _52157_ (_00575_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _52158_ (_00576_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _52159_ (_00577_, _00576_, _00575_);
  and _52160_ (_39357_, _00577_, _41806_);
  and _52161_ (_00578_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _52162_ (_00579_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _52163_ (_00580_, _00579_, _00578_);
  and _52164_ (_39358_, _00580_, _41806_);
  and _52165_ (_00581_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _52166_ (_00582_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _52167_ (_00583_, _00582_, _00581_);
  and _52168_ (_39359_, _00583_, _41806_);
  and _52169_ (_00584_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _52170_ (_00585_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _52171_ (_00586_, _00585_, _00584_);
  and _52172_ (_39361_, _00586_, _41806_);
  and _52173_ (_00587_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _52174_ (_00588_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _52175_ (_00589_, _00588_, _00587_);
  and _52176_ (_39362_, _00589_, _41806_);
  and _52177_ (_00590_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _52178_ (_00591_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _52179_ (_00592_, _00591_, _00590_);
  and _52180_ (_39363_, _00592_, _41806_);
  and _52181_ (_00593_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _52182_ (_00594_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _52183_ (_00595_, _00594_, _00593_);
  and _52184_ (_39364_, _00595_, _41806_);
  and _52185_ (_00596_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _52186_ (_00597_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _52187_ (_00598_, _00597_, _00596_);
  and _52188_ (_39365_, _00598_, _41806_);
  and _52189_ (_00599_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _52190_ (_00600_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _52191_ (_00601_, _00600_, _00599_);
  and _52192_ (_39366_, _00601_, _41806_);
  and _52193_ (_00602_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _52194_ (_00603_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _52195_ (_00604_, _00603_, _00602_);
  and _52196_ (_39367_, _00604_, _41806_);
  and _52197_ (_00605_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _52198_ (_00606_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _52199_ (_00607_, _00606_, _00605_);
  and _52200_ (_39368_, _00607_, _41806_);
  and _52201_ (_00608_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52202_ (_00609_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _52203_ (_00610_, _00609_, _00608_);
  and _52204_ (_39369_, _00610_, _41806_);
  and _52205_ (_00611_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52206_ (_00612_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _52207_ (_00613_, _00612_, _00611_);
  and _52208_ (_39370_, _00613_, _41806_);
  and _52209_ (_00614_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52210_ (_00615_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _52211_ (_00616_, _00615_, _00614_);
  and _52212_ (_39372_, _00616_, _41806_);
  and _52213_ (_00617_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52214_ (_00618_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _52215_ (_00619_, _00618_, _00617_);
  and _52216_ (_39373_, _00619_, _41806_);
  and _52217_ (_00620_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52218_ (_00621_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _52219_ (_00622_, _00621_, _00620_);
  and _52220_ (_39374_, _00622_, _41806_);
  and _52221_ (_00623_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52222_ (_00624_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _52223_ (_00625_, _00624_, _00623_);
  and _52224_ (_39375_, _00625_, _41806_);
  and _52225_ (_00626_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52226_ (_00627_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _52227_ (_00628_, _00627_, _00626_);
  and _52228_ (_39376_, _00628_, _41806_);
  and _52229_ (_00629_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52230_ (_00630_, _40408_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52231_ (_00631_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _52232_ (_00632_, _00631_, _43905_);
  and _52233_ (_00633_, _00632_, _00630_);
  or _52234_ (_00634_, _00633_, _00629_);
  and _52235_ (_39377_, _00634_, _41806_);
  and _52236_ (_00635_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52237_ (_00636_, _40564_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52238_ (_00637_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _52239_ (_00638_, _00637_, _43905_);
  and _52240_ (_00639_, _00638_, _00636_);
  or _52241_ (_00640_, _00639_, _00635_);
  and _52242_ (_39378_, _00640_, _41806_);
  and _52243_ (_00641_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52244_ (_00642_, _40492_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52245_ (_00643_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _52246_ (_00644_, _00643_, _43905_);
  and _52247_ (_00645_, _00644_, _00642_);
  or _52248_ (_00646_, _00645_, _00641_);
  and _52249_ (_39379_, _00646_, _41806_);
  and _52250_ (_00647_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52251_ (_00648_, _40370_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52252_ (_00649_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _52253_ (_00650_, _00649_, _43905_);
  and _52254_ (_00651_, _00650_, _00648_);
  or _52255_ (_00652_, _00651_, _00647_);
  and _52256_ (_39380_, _00652_, _41806_);
  and _52257_ (_00653_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52258_ (_00654_, _40540_, _43912_);
  or _52259_ (_00655_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _52260_ (_00656_, _00655_, _43905_);
  and _52261_ (_00657_, _00656_, _00654_);
  or _52262_ (_00658_, _00657_, _00653_);
  and _52263_ (_39381_, _00658_, _41806_);
  and _52264_ (_00659_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52265_ (_00660_, _40442_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52266_ (_00661_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _52267_ (_00662_, _00661_, _43905_);
  and _52268_ (_00663_, _00662_, _00660_);
  or _52269_ (_00664_, _00663_, _00659_);
  and _52270_ (_39383_, _00664_, _41806_);
  and _52271_ (_00665_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52272_ (_00666_, _40639_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52273_ (_00667_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _52274_ (_00668_, _00667_, _43905_);
  and _52275_ (_00669_, _00668_, _00666_);
  or _52276_ (_00670_, _00669_, _00665_);
  and _52277_ (_39384_, _00670_, _41806_);
  and _52278_ (_00671_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52279_ (_00672_, _40300_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52280_ (_00673_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _52281_ (_00674_, _00673_, _43905_);
  and _52282_ (_00675_, _00674_, _00672_);
  or _52283_ (_00676_, _00675_, _00671_);
  and _52284_ (_39385_, _00676_, _41806_);
  and _52285_ (_00677_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _52286_ (_00678_, _00677_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52287_ (_00679_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _43905_);
  and _52288_ (_00680_, _00679_, _41806_);
  and _52289_ (_39386_, _00680_, _00678_);
  and _52290_ (_00681_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _52291_ (_00682_, _00681_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52292_ (_00683_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _43905_);
  and _52293_ (_00684_, _00683_, _41806_);
  and _52294_ (_39387_, _00684_, _00682_);
  and _52295_ (_00685_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _52296_ (_00686_, _00685_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52297_ (_00687_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _43905_);
  and _52298_ (_00688_, _00687_, _41806_);
  and _52299_ (_39388_, _00688_, _00686_);
  and _52300_ (_00689_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _52301_ (_00690_, _00689_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52302_ (_00691_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _43905_);
  and _52303_ (_00692_, _00691_, _41806_);
  and _52304_ (_39389_, _00692_, _00690_);
  and _52305_ (_00693_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _52306_ (_00694_, _00693_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52307_ (_00695_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _43905_);
  and _52308_ (_00696_, _00695_, _41806_);
  and _52309_ (_39390_, _00696_, _00694_);
  and _52310_ (_00697_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _52311_ (_00698_, _00697_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52312_ (_00699_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _43905_);
  and _52313_ (_00700_, _00699_, _41806_);
  and _52314_ (_39391_, _00700_, _00698_);
  and _52315_ (_00701_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _52316_ (_00702_, _00701_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52317_ (_00703_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _43905_);
  and _52318_ (_00704_, _00703_, _41806_);
  and _52319_ (_39392_, _00704_, _00702_);
  nand _52320_ (_00705_, _43919_, _29231_);
  or _52321_ (_00706_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _52322_ (_00707_, _00706_, _41806_);
  and _52323_ (_39394_, _00707_, _00705_);
  nand _52324_ (_00708_, _43919_, _29893_);
  or _52325_ (_00709_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _52326_ (_00710_, _00709_, _41806_);
  and _52327_ (_39395_, _00710_, _00708_);
  nand _52328_ (_00711_, _43919_, _30567_);
  or _52329_ (_00712_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _52330_ (_00713_, _00712_, _41806_);
  and _52331_ (_39396_, _00713_, _00711_);
  nand _52332_ (_00714_, _43919_, _31338_);
  or _52333_ (_00715_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _52334_ (_00716_, _00715_, _41806_);
  and _52335_ (_39397_, _00716_, _00714_);
  nand _52336_ (_00717_, _43919_, _32044_);
  or _52337_ (_00718_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _52338_ (_00719_, _00718_, _41806_);
  and _52339_ (_39398_, _00719_, _00717_);
  nand _52340_ (_00720_, _43919_, _32853_);
  or _52341_ (_00721_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _52342_ (_00722_, _00721_, _41806_);
  and _52343_ (_39399_, _00722_, _00720_);
  nand _52344_ (_00723_, _43919_, _33598_);
  or _52345_ (_00724_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _52346_ (_00725_, _00724_, _41806_);
  and _52347_ (_39400_, _00725_, _00723_);
  nand _52348_ (_00726_, _43919_, _28011_);
  or _52349_ (_00727_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _52350_ (_00728_, _00727_, _41806_);
  and _52351_ (_39401_, _00728_, _00726_);
  nand _52352_ (_00729_, _43919_, _38617_);
  or _52353_ (_00730_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _52354_ (_00731_, _00730_, _41806_);
  and _52355_ (_39402_, _00731_, _00729_);
  nand _52356_ (_00732_, _43919_, _38645_);
  or _52357_ (_00733_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _52358_ (_00734_, _00733_, _41806_);
  and _52359_ (_39403_, _00734_, _00732_);
  nand _52360_ (_00735_, _43919_, _38673_);
  or _52361_ (_00736_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _52362_ (_00737_, _00736_, _41806_);
  and _52363_ (_39405_, _00737_, _00735_);
  nand _52364_ (_00738_, _43919_, _38702_);
  or _52365_ (_00739_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _52366_ (_00740_, _00739_, _41806_);
  and _52367_ (_39406_, _00740_, _00738_);
  nand _52368_ (_00741_, _43919_, _38731_);
  or _52369_ (_00742_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _52370_ (_00743_, _00742_, _41806_);
  and _52371_ (_39407_, _00743_, _00741_);
  nand _52372_ (_00744_, _43919_, _38760_);
  or _52373_ (_00745_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _52374_ (_00746_, _00745_, _41806_);
  and _52375_ (_39408_, _00746_, _00744_);
  nand _52376_ (_00747_, _43919_, _38787_);
  or _52377_ (_00748_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _52378_ (_00749_, _00748_, _41806_);
  and _52379_ (_39409_, _00749_, _00747_);
  nor _52380_ (_39617_, _40339_, rst);
  nor _52381_ (_00750_, _40703_, _40463_);
  nor _52382_ (_00751_, _40547_, _40327_);
  and _52383_ (_00752_, _00751_, _40380_);
  and _52384_ (_00753_, _00752_, _00750_);
  not _52385_ (_00754_, _00753_);
  nor _52386_ (_00755_, _00754_, _39024_);
  and _52387_ (_00756_, _40380_, _40547_);
  and _52388_ (_00757_, _00756_, _40463_);
  nor _52389_ (_00758_, _40703_, _40327_);
  and _52390_ (_00759_, _00758_, _00757_);
  not _52391_ (_00760_, _40500_);
  nor _52392_ (_00761_, _39128_, _39116_);
  and _52393_ (_00762_, _39128_, _39116_);
  nor _52394_ (_00763_, _00762_, _00761_);
  nor _52395_ (_00764_, _39140_, _39048_);
  and _52396_ (_00765_, _39140_, _39048_);
  nor _52397_ (_00766_, _00765_, _00764_);
  and _52398_ (_00767_, _00766_, _00763_);
  nor _52399_ (_00768_, _00766_, _00763_);
  or _52400_ (_00769_, _00768_, _00767_);
  and _52401_ (_00770_, _39073_, _39060_);
  nor _52402_ (_00771_, _39073_, _39060_);
  or _52403_ (_00772_, _00771_, _00770_);
  not _52404_ (_00773_, _00772_);
  nor _52405_ (_00774_, _39104_, _39093_);
  and _52406_ (_00775_, _39104_, _39093_);
  or _52407_ (_00776_, _00775_, _00774_);
  and _52408_ (_00777_, _00776_, _00773_);
  nor _52409_ (_00778_, _00776_, _00773_);
  nor _52410_ (_00779_, _00778_, _00777_);
  nor _52411_ (_00780_, _00779_, _00769_);
  and _52412_ (_00781_, _00779_, _00769_);
  nor _52413_ (_00782_, _00781_, _00780_);
  nor _52414_ (_00783_, _00782_, _00760_);
  and _52415_ (_00784_, _40415_, _40611_);
  nand _52416_ (_00785_, _00760_, _38964_);
  nand _52417_ (_00786_, _00785_, _00784_);
  or _52418_ (_00787_, _00786_, _00783_);
  not _52419_ (_00788_, _40415_);
  and _52420_ (_00789_, _00788_, _40611_);
  not _52421_ (_00790_, _00789_);
  and _52422_ (_00791_, _00760_, _38971_);
  and _52423_ (_00792_, _40500_, _38870_);
  nor _52424_ (_00793_, _00792_, _00791_);
  or _52425_ (_00794_, _00793_, _00790_);
  nor _52426_ (_00795_, _40415_, _40611_);
  not _52427_ (_00796_, _00795_);
  and _52428_ (_00797_, _00760_, _38862_);
  and _52429_ (_00798_, _40500_, _38933_);
  or _52430_ (_00799_, _00798_, _00797_);
  or _52431_ (_00800_, _00799_, _00796_);
  and _52432_ (_00801_, _00800_, _00794_);
  nor _52433_ (_00802_, _00760_, _38907_);
  nor _52434_ (_00803_, _00788_, _40611_);
  nand _52435_ (_00804_, _00760_, _39004_);
  nand _52436_ (_00805_, _00804_, _00803_);
  or _52437_ (_00806_, _00805_, _00802_);
  and _52438_ (_00807_, _00806_, _00801_);
  nand _52439_ (_00808_, _00807_, _00787_);
  and _52440_ (_00809_, _00808_, _00759_);
  and _52441_ (_00810_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _52442_ (_00811_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _52443_ (_00812_, _00811_, _00810_);
  and _52444_ (_00813_, _00812_, _00803_);
  or _52445_ (_00814_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _52446_ (_00815_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _52447_ (_00816_, _00815_, _00789_);
  and _52448_ (_00817_, _00816_, _00814_);
  and _52449_ (_00818_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _52450_ (_00819_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _52451_ (_00820_, _00819_, _00818_);
  and _52452_ (_00821_, _00820_, _00795_);
  nand _52453_ (_00822_, _40500_, _39870_);
  or _52454_ (_00823_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _52455_ (_00824_, _00823_, _00784_);
  and _52456_ (_00825_, _00824_, _00822_);
  or _52457_ (_00826_, _00825_, _00821_);
  or _52458_ (_00827_, _00826_, _00817_);
  or _52459_ (_00828_, _00827_, _00813_);
  and _52460_ (_00829_, _40703_, _40463_);
  and _52461_ (_00830_, _00751_, _40381_);
  and _52462_ (_00831_, _00830_, _00829_);
  and _52463_ (_00832_, _00831_, _00828_);
  and _52464_ (_00833_, _40703_, _40464_);
  and _52465_ (_00834_, _00830_, _00833_);
  and _52466_ (_00835_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _52467_ (_00836_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _52468_ (_00837_, _00836_, _00835_);
  and _52469_ (_00838_, _00837_, _00803_);
  or _52470_ (_00839_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _52471_ (_00840_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _52472_ (_00841_, _00840_, _00789_);
  and _52473_ (_00842_, _00841_, _00839_);
  nor _52474_ (_00843_, _40500_, _39908_);
  and _52475_ (_00844_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _52476_ (_00845_, _00844_, _00843_);
  and _52477_ (_00846_, _00845_, _00795_);
  or _52478_ (_00847_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _52479_ (_00848_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _52480_ (_00849_, _00848_, _00784_);
  and _52481_ (_00850_, _00849_, _00847_);
  or _52482_ (_00851_, _00850_, _00846_);
  or _52483_ (_00852_, _00851_, _00842_);
  or _52484_ (_00853_, _00852_, _00838_);
  and _52485_ (_00854_, _00853_, _00834_);
  nor _52486_ (_00855_, _00854_, _00832_);
  nor _52487_ (_00856_, _42622_, _37475_);
  and _52488_ (_00857_, _36069_, _37646_);
  or _52489_ (_00858_, _00857_, _37095_);
  nor _52490_ (_00859_, _00858_, _35839_);
  and _52491_ (_00860_, _42461_, _35915_);
  and _52492_ (_00861_, _34793_, _42458_);
  or _52493_ (_00863_, _00861_, _00860_);
  or _52494_ (_00864_, _00863_, _42524_);
  nor _52495_ (_00865_, _00864_, _37133_);
  and _52496_ (_00866_, _00865_, _00859_);
  nor _52497_ (_00867_, _42457_, _37056_);
  and _52498_ (_00868_, _00867_, _42526_);
  and _52499_ (_00869_, _00868_, _00866_);
  and _52500_ (_00870_, _00869_, _37373_);
  and _52501_ (_00871_, _00870_, _00856_);
  nor _52502_ (_00872_, _00871_, _33817_);
  and _52503_ (_00873_, _43004_, p2in_reg[2]);
  and _52504_ (_00874_, _43000_, p2_in[2]);
  nor _52505_ (_00875_, _00874_, _00873_);
  nor _52506_ (_00876_, _00875_, _00872_);
  and _52507_ (_00877_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _52508_ (_00878_, _00877_, _00876_);
  nor _52509_ (_00879_, _00878_, _00760_);
  and _52510_ (_00880_, _43004_, p2in_reg[6]);
  and _52511_ (_00881_, _43000_, p2_in[6]);
  nor _52512_ (_00882_, _00881_, _00880_);
  nor _52513_ (_00883_, _00882_, _00872_);
  and _52514_ (_00884_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _52515_ (_00885_, _00884_, _00883_);
  or _52516_ (_00886_, _00885_, _40500_);
  nand _52517_ (_00887_, _00886_, _00803_);
  or _52518_ (_00888_, _00887_, _00879_);
  not _52519_ (_00889_, _00784_);
  and _52520_ (_00890_, _43004_, p2in_reg[4]);
  and _52521_ (_00891_, _43000_, p2_in[4]);
  nor _52522_ (_00892_, _00891_, _00890_);
  nor _52523_ (_00894_, _00892_, _00872_);
  and _52524_ (_00895_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _52525_ (_00896_, _00895_, _00894_);
  nand _52526_ (_00897_, _00896_, _00760_);
  and _52527_ (_00898_, _43004_, p2in_reg[0]);
  and _52528_ (_00899_, _43000_, p2_in[0]);
  nor _52529_ (_00900_, _00899_, _00898_);
  nor _52530_ (_00901_, _00900_, _00872_);
  and _52531_ (_00902_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _52532_ (_00903_, _00902_, _00901_);
  nand _52533_ (_00904_, _00903_, _40500_);
  and _52534_ (_00905_, _00904_, _00897_);
  or _52535_ (_00906_, _00905_, _00889_);
  and _52536_ (_00907_, _43004_, p2in_reg[7]);
  and _52537_ (_00908_, _43000_, p2_in[7]);
  nor _52538_ (_00909_, _00908_, _00907_);
  nor _52539_ (_00910_, _00909_, _00872_);
  and _52540_ (_00911_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _52541_ (_00912_, _00911_, _00910_);
  nand _52542_ (_00913_, _00912_, _00760_);
  and _52543_ (_00915_, _43004_, p2in_reg[3]);
  and _52544_ (_00916_, _43000_, p2_in[3]);
  nor _52545_ (_00917_, _00916_, _00915_);
  nor _52546_ (_00918_, _00917_, _00872_);
  and _52547_ (_00919_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _52548_ (_00920_, _00919_, _00918_);
  nand _52549_ (_00921_, _00920_, _40500_);
  and _52550_ (_00922_, _00921_, _00913_);
  or _52551_ (_00923_, _00922_, _00796_);
  and _52552_ (_00924_, _00923_, _00906_);
  and _52553_ (_00925_, _43004_, p2in_reg[1]);
  and _52554_ (_00926_, _43000_, p2_in[1]);
  nor _52555_ (_00927_, _00926_, _00925_);
  nor _52556_ (_00928_, _00927_, _00872_);
  and _52557_ (_00929_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _52558_ (_00930_, _00929_, _00928_);
  nor _52559_ (_00931_, _00930_, _00760_);
  and _52560_ (_00932_, _43004_, p2in_reg[5]);
  and _52561_ (_00933_, _43000_, p2_in[5]);
  nor _52562_ (_00934_, _00933_, _00932_);
  nor _52563_ (_00935_, _00934_, _00872_);
  and _52564_ (_00936_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _52565_ (_00937_, _00936_, _00935_);
  or _52566_ (_00938_, _00937_, _40500_);
  nand _52567_ (_00939_, _00938_, _00789_);
  or _52568_ (_00940_, _00939_, _00931_);
  and _52569_ (_00941_, _00940_, _00924_);
  and _52570_ (_00942_, _00941_, _00888_);
  nand _52571_ (_00943_, _00833_, _00752_);
  or _52572_ (_00944_, _00943_, _00942_);
  and _52573_ (_00945_, _00944_, _00855_);
  not _52574_ (_00946_, _40327_);
  and _52575_ (_00947_, _00756_, _00946_);
  and _52576_ (_00948_, _00947_, _00750_);
  nand _52577_ (_00949_, _40500_, _29264_);
  or _52578_ (_00950_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _52579_ (_00951_, _00950_, _00784_);
  and _52580_ (_00952_, _00951_, _00949_);
  nor _52581_ (_00953_, _40500_, _28098_);
  and _52582_ (_00954_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _52583_ (_00955_, _00954_, _00953_);
  and _52584_ (_00956_, _00955_, _00795_);
  nor _52585_ (_00957_, _40500_, _33631_);
  and _52586_ (_00958_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _52587_ (_00959_, _00958_, _00957_);
  and _52588_ (_00960_, _00959_, _00803_);
  nand _52589_ (_00961_, _40500_, _29926_);
  or _52590_ (_00962_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _52591_ (_00963_, _00962_, _00789_);
  and _52592_ (_00964_, _00963_, _00961_);
  or _52593_ (_00965_, _00964_, _00960_);
  or _52594_ (_00966_, _00965_, _00956_);
  or _52595_ (_00967_, _00966_, _00952_);
  and _52596_ (_00968_, _00967_, _00948_);
  nor _52597_ (_00969_, _40380_, _40327_);
  and _52598_ (_00970_, _40703_, _40547_);
  and _52599_ (_00971_, _00970_, _00969_);
  and _52600_ (_00972_, _00971_, _40464_);
  nand _52601_ (_00973_, _40500_, _39920_);
  or _52602_ (_00974_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _52603_ (_00975_, _00974_, _00784_);
  and _52604_ (_00976_, _00975_, _00973_);
  and _52605_ (_00977_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _52606_ (_00978_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _52607_ (_00979_, _00978_, _00977_);
  and _52608_ (_00980_, _00979_, _00795_);
  and _52609_ (_00981_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _52610_ (_00982_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _52611_ (_00983_, _00982_, _00981_);
  and _52612_ (_00984_, _00983_, _00803_);
  nand _52613_ (_00985_, _40500_, _39922_);
  or _52614_ (_00986_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _52615_ (_00987_, _00986_, _00789_);
  and _52616_ (_00988_, _00987_, _00985_);
  or _52617_ (_00989_, _00988_, _00984_);
  or _52618_ (_00990_, _00989_, _00980_);
  or _52619_ (_00991_, _00990_, _00976_);
  and _52620_ (_00992_, _00991_, _00972_);
  nor _52621_ (_00993_, _00992_, _00968_);
  nand _52622_ (_00994_, _00947_, _00833_);
  and _52623_ (_00995_, _43004_, p3in_reg[2]);
  and _52624_ (_00996_, _43000_, p3_in[2]);
  nor _52625_ (_00997_, _00996_, _00995_);
  nor _52626_ (_00998_, _00997_, _00872_);
  and _52627_ (_00999_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _52628_ (_01000_, _00999_, _00998_);
  nor _52629_ (_01001_, _01000_, _00760_);
  and _52630_ (_01002_, _43004_, p3in_reg[6]);
  and _52631_ (_01003_, _43000_, p3_in[6]);
  nor _52632_ (_01004_, _01003_, _01002_);
  nor _52633_ (_01005_, _01004_, _00872_);
  and _52634_ (_01006_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _52635_ (_01007_, _01006_, _01005_);
  or _52636_ (_01008_, _01007_, _40500_);
  nand _52637_ (_01009_, _01008_, _00803_);
  or _52638_ (_01010_, _01009_, _01001_);
  and _52639_ (_01011_, _43004_, p3in_reg[4]);
  and _52640_ (_01012_, _43000_, p3_in[4]);
  nor _52641_ (_01013_, _01012_, _01011_);
  nor _52642_ (_01014_, _01013_, _00872_);
  and _52643_ (_01015_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _52644_ (_01016_, _01015_, _01014_);
  nand _52645_ (_01017_, _01016_, _00760_);
  and _52646_ (_01018_, _43004_, p3in_reg[0]);
  and _52647_ (_01019_, _43000_, p3_in[0]);
  nor _52648_ (_01020_, _01019_, _01018_);
  nor _52649_ (_01021_, _01020_, _00872_);
  and _52650_ (_01022_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _52651_ (_01023_, _01022_, _01021_);
  nand _52652_ (_01024_, _01023_, _40500_);
  and _52653_ (_01025_, _01024_, _01017_);
  or _52654_ (_01026_, _01025_, _00889_);
  and _52655_ (_01027_, _43004_, p3in_reg[7]);
  and _52656_ (_01028_, _43000_, p3_in[7]);
  nor _52657_ (_01029_, _01028_, _01027_);
  nor _52658_ (_01030_, _01029_, _00872_);
  and _52659_ (_01031_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _52660_ (_01032_, _01031_, _01030_);
  nand _52661_ (_01033_, _01032_, _00760_);
  and _52662_ (_01034_, _43004_, p3in_reg[3]);
  and _52663_ (_01035_, _43000_, p3_in[3]);
  nor _52664_ (_01036_, _01035_, _01034_);
  nor _52665_ (_01037_, _01036_, _00872_);
  and _52666_ (_01038_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _52667_ (_01039_, _01038_, _01037_);
  nand _52668_ (_01040_, _01039_, _40500_);
  and _52669_ (_01041_, _01040_, _01033_);
  or _52670_ (_01042_, _01041_, _00796_);
  and _52671_ (_01043_, _01042_, _01026_);
  and _52672_ (_01044_, _43004_, p3in_reg[1]);
  and _52673_ (_01045_, _43000_, p3_in[1]);
  nor _52674_ (_01046_, _01045_, _01044_);
  nor _52675_ (_01047_, _01046_, _00872_);
  and _52676_ (_01048_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _52677_ (_01049_, _01048_, _01047_);
  nor _52678_ (_01050_, _01049_, _00760_);
  and _52679_ (_01051_, _43004_, p3in_reg[5]);
  and _52680_ (_01052_, _43000_, p3_in[5]);
  nor _52681_ (_01053_, _01052_, _01051_);
  nor _52682_ (_01054_, _01053_, _00872_);
  and _52683_ (_01055_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _52684_ (_01056_, _01055_, _01054_);
  or _52685_ (_01057_, _01056_, _40500_);
  nand _52686_ (_01058_, _01057_, _00789_);
  or _52687_ (_01059_, _01058_, _01050_);
  and _52688_ (_01060_, _01059_, _01043_);
  and _52689_ (_01061_, _01060_, _01010_);
  or _52690_ (_01062_, _01061_, _00994_);
  and _52691_ (_01063_, _01062_, _00993_);
  and _52692_ (_01064_, _00830_, _40703_);
  or _52693_ (_01065_, _01064_, _00948_);
  nor _52694_ (_01066_, _01065_, _00759_);
  nor _52695_ (_01067_, _40381_, _40327_);
  and _52696_ (_01068_, _01067_, _40703_);
  nor _52697_ (_01069_, _01068_, _00971_);
  and _52698_ (_01070_, _01069_, _00754_);
  and _52699_ (_01071_, _01070_, _01066_);
  nand _52700_ (_01072_, _43104_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or _52701_ (_01073_, _01072_, _01071_);
  nand _52702_ (_01074_, _00947_, _00829_);
  and _52703_ (_01075_, _43004_, p1in_reg[5]);
  and _52704_ (_01076_, _43000_, p1_in[5]);
  nor _52705_ (_01077_, _01076_, _01075_);
  nor _52706_ (_01078_, _01077_, _00872_);
  and _52707_ (_01079_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _52708_ (_01080_, _01079_, _01078_);
  nand _52709_ (_01081_, _01080_, _00760_);
  and _52710_ (_01082_, _43004_, p1in_reg[1]);
  and _52711_ (_01083_, _43000_, p1_in[1]);
  nor _52712_ (_01084_, _01083_, _01082_);
  nor _52713_ (_01085_, _01084_, _00872_);
  and _52714_ (_01086_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _52715_ (_01087_, _01086_, _01085_);
  nand _52716_ (_01088_, _01087_, _40500_);
  and _52717_ (_01089_, _01088_, _01081_);
  or _52718_ (_01090_, _01089_, _00790_);
  and _52719_ (_01091_, _43004_, p1in_reg[7]);
  and _52720_ (_01092_, _43000_, p1_in[7]);
  nor _52721_ (_01093_, _01092_, _01091_);
  nor _52722_ (_01094_, _01093_, _00872_);
  and _52723_ (_01095_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _52724_ (_01096_, _01095_, _01094_);
  nand _52725_ (_01097_, _01096_, _00760_);
  and _52726_ (_01098_, _43004_, p1in_reg[3]);
  and _52727_ (_01099_, _43000_, p1_in[3]);
  nor _52728_ (_01100_, _01099_, _01098_);
  nor _52729_ (_01101_, _01100_, _00872_);
  and _52730_ (_01102_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _52731_ (_01103_, _01102_, _01101_);
  nand _52732_ (_01104_, _01103_, _40500_);
  and _52733_ (_01105_, _01104_, _01097_);
  or _52734_ (_01106_, _01105_, _00796_);
  and _52735_ (_01107_, _01106_, _01090_);
  not _52736_ (_01108_, _00803_);
  and _52737_ (_01109_, _43004_, p1in_reg[6]);
  and _52738_ (_01110_, _43000_, p1_in[6]);
  nor _52739_ (_01111_, _01110_, _01109_);
  nor _52740_ (_01112_, _01111_, _00872_);
  and _52741_ (_01113_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _52742_ (_01114_, _01113_, _01112_);
  nand _52743_ (_01115_, _01114_, _00760_);
  and _52744_ (_01116_, _43004_, p1in_reg[2]);
  and _52745_ (_01117_, _43000_, p1_in[2]);
  nor _52746_ (_01118_, _01117_, _01116_);
  nor _52747_ (_01119_, _01118_, _00872_);
  and _52748_ (_01120_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _52749_ (_01121_, _01120_, _01119_);
  nand _52750_ (_01122_, _01121_, _40500_);
  and _52751_ (_01123_, _01122_, _01115_);
  or _52752_ (_01124_, _01123_, _01108_);
  and _52753_ (_01125_, _43004_, p1in_reg[4]);
  and _52754_ (_01126_, _43000_, p1_in[4]);
  nor _52755_ (_01127_, _01126_, _01125_);
  nor _52756_ (_01128_, _01127_, _00872_);
  and _52757_ (_01129_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _52758_ (_01130_, _01129_, _01128_);
  nand _52759_ (_01131_, _01130_, _00760_);
  and _52760_ (_01132_, _43004_, p1in_reg[0]);
  and _52761_ (_01133_, _43000_, p1_in[0]);
  nor _52762_ (_01134_, _01133_, _01132_);
  nor _52763_ (_01135_, _01134_, _00872_);
  and _52764_ (_01136_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _52765_ (_01137_, _01136_, _01135_);
  nand _52766_ (_01138_, _01137_, _40500_);
  and _52767_ (_01139_, _01138_, _01131_);
  or _52768_ (_01140_, _01139_, _00889_);
  and _52769_ (_01141_, _01140_, _01124_);
  and _52770_ (_01142_, _01141_, _01107_);
  or _52771_ (_01143_, _01142_, _01074_);
  and _52772_ (_01144_, _00829_, _00752_);
  and _52773_ (_01145_, _43004_, p0in_reg[5]);
  and _52774_ (_01146_, _43000_, p0_in[5]);
  nor _52775_ (_01147_, _01146_, _01145_);
  nor _52776_ (_01148_, _01147_, _00872_);
  and _52777_ (_01149_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _52778_ (_01150_, _01149_, _01148_);
  nand _52779_ (_01151_, _01150_, _00760_);
  and _52780_ (_01152_, _43004_, p0in_reg[1]);
  and _52781_ (_01153_, _43000_, p0_in[1]);
  nor _52782_ (_01154_, _01153_, _01152_);
  nor _52783_ (_01155_, _01154_, _00872_);
  and _52784_ (_01156_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _52785_ (_01157_, _01156_, _01155_);
  nand _52786_ (_01158_, _01157_, _40500_);
  and _52787_ (_01159_, _01158_, _01151_);
  or _52788_ (_01160_, _01159_, _00790_);
  and _52789_ (_01161_, _43004_, p0in_reg[4]);
  and _52790_ (_01162_, _43000_, p0_in[4]);
  nor _52791_ (_01163_, _01162_, _01161_);
  nor _52792_ (_01164_, _01163_, _00872_);
  and _52793_ (_01165_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _52794_ (_01166_, _01165_, _01164_);
  nand _52795_ (_01167_, _01166_, _00760_);
  and _52796_ (_01168_, _43004_, p0in_reg[0]);
  and _52797_ (_01169_, _43000_, p0_in[0]);
  nor _52798_ (_01170_, _01169_, _01168_);
  nor _52799_ (_01171_, _01170_, _00872_);
  and _52800_ (_01172_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or _52801_ (_01173_, _01172_, _01171_);
  nand _52802_ (_01174_, _01173_, _40500_);
  and _52803_ (_01175_, _01174_, _01167_);
  or _52804_ (_01176_, _01175_, _00889_);
  and _52805_ (_01177_, _01176_, _01160_);
  and _52806_ (_01178_, _43004_, p0in_reg[6]);
  and _52807_ (_01179_, _43000_, p0_in[6]);
  nor _52808_ (_01180_, _01179_, _01178_);
  nor _52809_ (_01181_, _01180_, _00872_);
  and _52810_ (_01182_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _52811_ (_01183_, _01182_, _01181_);
  nand _52812_ (_01184_, _01183_, _00760_);
  and _52813_ (_01185_, _43004_, p0in_reg[2]);
  and _52814_ (_01186_, _43000_, p0_in[2]);
  nor _52815_ (_01187_, _01186_, _01185_);
  nor _52816_ (_01188_, _01187_, _00872_);
  and _52817_ (_01189_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _52818_ (_01190_, _01189_, _01188_);
  nand _52819_ (_01191_, _01190_, _40500_);
  and _52820_ (_01192_, _01191_, _01184_);
  or _52821_ (_01193_, _01192_, _01108_);
  and _52822_ (_01194_, _43004_, p0in_reg[7]);
  and _52823_ (_01195_, _43000_, p0_in[7]);
  nor _52824_ (_01196_, _01195_, _01194_);
  nor _52825_ (_01197_, _01196_, _00872_);
  and _52826_ (_01198_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _52827_ (_01199_, _01198_, _01197_);
  nand _52828_ (_01200_, _01199_, _00760_);
  and _52829_ (_01201_, _43004_, p0in_reg[3]);
  and _52830_ (_01202_, _43000_, p0_in[3]);
  nor _52831_ (_01203_, _01202_, _01201_);
  nor _52832_ (_01204_, _01203_, _00872_);
  and _52833_ (_01205_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _52834_ (_01206_, _01205_, _01204_);
  nand _52835_ (_01207_, _01206_, _40500_);
  and _52836_ (_01208_, _01207_, _01200_);
  or _52837_ (_01209_, _01208_, _00796_);
  and _52838_ (_01210_, _01209_, _01193_);
  nand _52839_ (_01211_, _01210_, _01177_);
  nand _52840_ (_01212_, _01211_, _01144_);
  and _52841_ (_01213_, _01212_, _01143_);
  and _52842_ (_01214_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _52843_ (_01215_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _52844_ (_01216_, _01215_, _01214_);
  and _52845_ (_01217_, _01216_, _00784_);
  or _52846_ (_01218_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _52847_ (_01219_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _52848_ (_01220_, _01219_, _00795_);
  and _52849_ (_01221_, _01220_, _01218_);
  and _52850_ (_01222_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _52851_ (_01223_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _52852_ (_01224_, _01223_, _01222_);
  and _52853_ (_01225_, _01224_, _00789_);
  nand _52854_ (_01226_, _40500_, _39082_);
  or _52855_ (_01227_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _52856_ (_01228_, _01227_, _00803_);
  and _52857_ (_01229_, _01228_, _01226_);
  or _52858_ (_01230_, _01229_, _01225_);
  or _52859_ (_01231_, _01230_, _01221_);
  or _52860_ (_01232_, _01231_, _01217_);
  nand _52861_ (_01233_, _01232_, _00753_);
  and _52862_ (_01234_, _01233_, _01213_);
  and _52863_ (_01235_, _01234_, _01073_);
  and _52864_ (_01236_, _01235_, _01063_);
  nand _52865_ (_01237_, _01236_, _00945_);
  or _52866_ (_01238_, _01237_, _00809_);
  or _52867_ (_01239_, _01073_, _29318_);
  and _52868_ (_01240_, _01239_, _01238_);
  or _52869_ (_01241_, _01240_, _00755_);
  and _52870_ (_01242_, _00789_, _39073_);
  and _52871_ (_01243_, _00784_, _39060_);
  or _52872_ (_01244_, _01243_, _01242_);
  nor _52873_ (_01245_, _00796_, _39104_);
  nor _52874_ (_01246_, _01108_, _39093_);
  or _52875_ (_01247_, _01246_, _01245_);
  or _52876_ (_01248_, _01247_, _01244_);
  and _52877_ (_01249_, _01248_, _40500_);
  and _52878_ (_01250_, _00789_, _39128_);
  and _52879_ (_01251_, _00795_, _39048_);
  or _52880_ (_01252_, _01251_, _01250_);
  and _52881_ (_01253_, _00784_, _39116_);
  and _52882_ (_01254_, _00803_, _39140_);
  or _52883_ (_01255_, _01254_, _01253_);
  or _52884_ (_01256_, _01255_, _01252_);
  nand _52885_ (_01257_, _01256_, _00760_);
  nand _52886_ (_01258_, _01257_, _00755_);
  or _52887_ (_01259_, _01258_, _01249_);
  and _52888_ (_01260_, _01259_, _01241_);
  not _52889_ (_01261_, _38817_);
  not _52890_ (_01262_, _00872_);
  and _52891_ (_01263_, _01068_, _01262_);
  nor _52892_ (_01264_, _01263_, _01261_);
  and _52893_ (_01265_, _01264_, _43027_);
  not _52894_ (_01266_, _01265_);
  nor _52895_ (_01267_, _01266_, _01071_);
  or _52896_ (_01268_, _01267_, _01260_);
  and _52897_ (_01269_, _00803_, _40633_);
  and _52898_ (_01270_, _00784_, _40538_);
  or _52899_ (_01271_, _01270_, _40500_);
  or _52900_ (_01272_, _01271_, _01269_);
  and _52901_ (_01273_, _00803_, _40482_);
  and _52902_ (_01274_, _00784_, _38426_);
  or _52903_ (_01275_, _01274_, _00760_);
  or _52904_ (_01276_, _01275_, _01273_);
  and _52905_ (_01277_, _01276_, _01272_);
  and _52906_ (_01278_, _40500_, _38418_);
  nor _52907_ (_01279_, _40500_, _38366_);
  or _52908_ (_01280_, _01279_, _01278_);
  and _52909_ (_01281_, _01280_, _00789_);
  and _52910_ (_01282_, _40500_, _40360_);
  nor _52911_ (_01283_, _40500_, _38162_);
  or _52912_ (_01284_, _01283_, _01282_);
  and _52913_ (_01285_, _01284_, _00795_);
  or _52914_ (_01286_, _01285_, _01281_);
  nor _52915_ (_01287_, _01286_, _01277_);
  nand _52916_ (_01288_, _01287_, _01267_);
  and _52917_ (_01289_, _01288_, _41806_);
  and _52918_ (_39648_, _01289_, _01268_);
  and _52919_ (_01290_, _40547_, _40463_);
  and _52920_ (_01291_, _40380_, _40500_);
  and _52921_ (_01292_, _01291_, _00784_);
  and _52922_ (_01293_, _01292_, _01290_);
  and _52923_ (_01294_, _01293_, _00758_);
  and _52924_ (_01295_, _01294_, _38823_);
  and _52925_ (_01296_, _00829_, _00751_);
  and _52926_ (_01297_, _01291_, _00795_);
  and _52927_ (_01298_, _01297_, _01296_);
  and _52928_ (_01299_, _01298_, _38493_);
  nor _52929_ (_01300_, _01299_, _01295_);
  nor _52930_ (_01301_, _01300_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _52931_ (_01302_, _01301_);
  nand _52932_ (_01303_, _39024_, _39022_);
  and _52933_ (_01304_, _00784_, _40500_);
  and _52934_ (_01305_, _01304_, _00753_);
  and _52935_ (_01306_, _01305_, _01303_);
  and _52936_ (_01307_, _00795_, _00760_);
  nor _52937_ (_01308_, _01307_, _38954_);
  and _52938_ (_01309_, _01308_, _43027_);
  nor _52939_ (_01310_, _01309_, _01306_);
  and _52940_ (_01311_, _01310_, _43107_);
  and _52941_ (_01312_, _01311_, _01302_);
  and _52942_ (_01313_, _01291_, _00803_);
  and _52943_ (_01314_, _01313_, _01296_);
  and _52944_ (_01315_, _01314_, _38493_);
  or _52945_ (_01316_, _01315_, rst);
  nor _52946_ (_39649_, _01316_, _01312_);
  not _52947_ (_01317_, _01315_);
  and _52948_ (_01318_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _52949_ (_01319_, _40703_, _00946_);
  and _52950_ (_01320_, _40547_, _40464_);
  and _52951_ (_01321_, _01320_, _01319_);
  and _52952_ (_01322_, _01304_, _40381_);
  and _52953_ (_01323_, _01322_, _01321_);
  and _52954_ (_01324_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _52955_ (_01325_, _01324_, _01318_);
  and _52956_ (_01326_, _01322_, _01296_);
  and _52957_ (_01327_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _52958_ (_01328_, _00833_, _00751_);
  and _52959_ (_01329_, _01328_, _01322_);
  and _52960_ (_01330_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _52961_ (_01331_, _01330_, _01327_);
  or _52962_ (_01332_, _01331_, _01325_);
  and _52963_ (_01333_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _52964_ (_01334_, _01320_, _00758_);
  and _52965_ (_01335_, _01334_, _01292_);
  and _52966_ (_01336_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _52967_ (_01337_, _01336_, _01333_);
  and _52968_ (_01338_, _01291_, _00789_);
  and _52969_ (_01339_, _01338_, _01296_);
  and _52970_ (_01340_, _01339_, _40266_);
  and _52971_ (_01341_, _01292_, _01321_);
  and _52972_ (_01342_, _01341_, _01032_);
  or _52973_ (_01343_, _01342_, _01340_);
  or _52974_ (_01344_, _01343_, _01337_);
  or _52975_ (_01345_, _01344_, _01332_);
  and _52976_ (_01346_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _52977_ (_01347_, _01328_, _01292_);
  and _52978_ (_01348_, _01347_, _00912_);
  and _52979_ (_01349_, _01319_, _01290_);
  and _52980_ (_01350_, _01349_, _01292_);
  and _52981_ (_01351_, _01350_, _01096_);
  or _52982_ (_01352_, _01351_, _01348_);
  and _52983_ (_01353_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _52984_ (_01354_, _01296_, _01292_);
  and _52985_ (_01355_, _01354_, _01199_);
  or _52986_ (_01356_, _01355_, _01353_);
  or _52987_ (_01357_, _01356_, _01352_);
  or _52988_ (_01358_, _01357_, _01346_);
  or _52989_ (_01359_, _01358_, _01345_);
  and _52990_ (_01360_, _01359_, _01312_);
  nor _52991_ (_01361_, _01312_, _17497_);
  or _52992_ (_01362_, _01361_, _01360_);
  and _52993_ (_01363_, _01362_, _01317_);
  nor _52994_ (_01364_, _01317_, _28011_);
  or _52995_ (_01365_, _01364_, _01363_);
  and _52996_ (_39650_, _01365_, _41806_);
  and _52997_ (_01366_, _01294_, _00782_);
  and _52998_ (_01367_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _52999_ (_01368_, _01304_, _01144_);
  and _53000_ (_01369_, _01368_, _01173_);
  and _53001_ (_01370_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _53002_ (_01371_, _01293_, _01319_);
  and _53003_ (_01372_, _01371_, _01137_);
  or _53004_ (_01373_, _01372_, _01370_);
  or _53005_ (_01374_, _01373_, _01369_);
  or _53006_ (_01375_, _01374_, _01367_);
  and _53007_ (_01376_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _53008_ (_01377_, _01341_, _01023_);
  or _53009_ (_01378_, _01377_, _01376_);
  and _53010_ (_01379_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _53011_ (_01380_, _01339_, _40411_);
  or _53012_ (_01381_, _01380_, _01379_);
  or _53013_ (_01382_, _01381_, _01378_);
  and _53014_ (_01383_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _53015_ (_01384_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _53016_ (_01385_, _01384_, _01383_);
  and _53017_ (_01386_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _53018_ (_01387_, _01347_, _00903_);
  or _53019_ (_01388_, _01387_, _01386_);
  or _53020_ (_01389_, _01388_, _01385_);
  or _53021_ (_01390_, _01389_, _01382_);
  nor _53022_ (_01391_, _01390_, _01375_);
  nand _53023_ (_01392_, _01391_, _01312_);
  or _53024_ (_01393_, _01392_, _01366_);
  or _53025_ (_01394_, _01312_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _53026_ (_01395_, _01394_, _01393_);
  or _53027_ (_01396_, _01395_, _01315_);
  nand _53028_ (_01397_, _01315_, _29231_);
  and _53029_ (_01398_, _01397_, _41806_);
  and _53030_ (_39713_, _01398_, _01396_);
  and _53031_ (_01399_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _53032_ (_01400_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or _53033_ (_01401_, _01400_, _01399_);
  and _53034_ (_01402_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _53035_ (_01403_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _53036_ (_01404_, _01403_, _01402_);
  or _53037_ (_01405_, _01404_, _01401_);
  and _53038_ (_01407_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _53039_ (_01409_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _53040_ (_01411_, _01409_, _01407_);
  and _53041_ (_01413_, _01341_, _01049_);
  and _53042_ (_01415_, _01339_, _40550_);
  or _53043_ (_01417_, _01415_, _01413_);
  or _53044_ (_01419_, _01417_, _01411_);
  or _53045_ (_01420_, _01419_, _01405_);
  and _53046_ (_01421_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _53047_ (_01422_, _01347_, _00930_);
  and _53048_ (_01423_, _01350_, _01087_);
  or _53049_ (_01424_, _01423_, _01422_);
  and _53050_ (_01425_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _53051_ (_01427_, _01354_, _01157_);
  or _53052_ (_01428_, _01427_, _01425_);
  or _53053_ (_01430_, _01428_, _01424_);
  or _53054_ (_01431_, _01430_, _01421_);
  or _53055_ (_01432_, _01431_, _01420_);
  and _53056_ (_01434_, _01432_, _01312_);
  nor _53057_ (_01435_, _01312_, _17323_);
  or _53058_ (_01436_, _01435_, _01434_);
  and _53059_ (_01438_, _01436_, _01317_);
  nor _53060_ (_01439_, _01317_, _29893_);
  or _53061_ (_01440_, _01439_, _01438_);
  and _53062_ (_39714_, _01440_, _41806_);
  and _53063_ (_01442_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _53064_ (_01443_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _53065_ (_01445_, _01443_, _01442_);
  and _53066_ (_01446_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _53067_ (_01447_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _53068_ (_01449_, _01447_, _01446_);
  or _53069_ (_01450_, _01449_, _01445_);
  and _53070_ (_01451_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _53071_ (_01453_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _53072_ (_01454_, _01453_, _01451_);
  and _53073_ (_01455_, _01339_, _40496_);
  and _53074_ (_01457_, _01341_, _01000_);
  or _53075_ (_01458_, _01457_, _01455_);
  or _53076_ (_01459_, _01458_, _01454_);
  or _53077_ (_01460_, _01459_, _01450_);
  and _53078_ (_01461_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _53079_ (_01462_, _01347_, _00878_);
  and _53080_ (_01463_, _01350_, _01121_);
  or _53081_ (_01464_, _01463_, _01462_);
  and _53082_ (_01465_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _53083_ (_01466_, _01354_, _01190_);
  or _53084_ (_01467_, _01466_, _01465_);
  or _53085_ (_01468_, _01467_, _01464_);
  or _53086_ (_01469_, _01468_, _01461_);
  or _53087_ (_01470_, _01469_, _01460_);
  and _53088_ (_01471_, _01470_, _01312_);
  nor _53089_ (_01472_, _01312_, _15975_);
  or _53090_ (_01473_, _01472_, _01471_);
  and _53091_ (_01474_, _01473_, _01317_);
  nor _53092_ (_01475_, _01317_, _30567_);
  or _53093_ (_01476_, _01475_, _01474_);
  and _53094_ (_39715_, _01476_, _41806_);
  and _53095_ (_01478_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _53096_ (_01479_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _53097_ (_01481_, _01479_, _01478_);
  and _53098_ (_01482_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _53099_ (_01483_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _53100_ (_01485_, _01483_, _01482_);
  or _53101_ (_01486_, _01485_, _01481_);
  and _53102_ (_01487_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _53103_ (_01489_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _53104_ (_01490_, _01489_, _01487_);
  and _53105_ (_01491_, _01341_, _01039_);
  and _53106_ (_01493_, _01339_, _40373_);
  or _53107_ (_01494_, _01493_, _01491_);
  or _53108_ (_01495_, _01494_, _01490_);
  or _53109_ (_01497_, _01495_, _01486_);
  and _53110_ (_01498_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _53111_ (_01499_, _01347_, _00920_);
  and _53112_ (_01501_, _01350_, _01103_);
  or _53113_ (_01502_, _01501_, _01499_);
  and _53114_ (_01503_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _53115_ (_01505_, _01354_, _01206_);
  or _53116_ (_01506_, _01505_, _01503_);
  or _53117_ (_01507_, _01506_, _01502_);
  or _53118_ (_01509_, _01507_, _01498_);
  or _53119_ (_01510_, _01509_, _01497_);
  and _53120_ (_01511_, _01510_, _01312_);
  nor _53121_ (_01512_, _01312_, _17007_);
  or _53122_ (_01513_, _01512_, _01511_);
  and _53123_ (_01514_, _01513_, _01317_);
  nor _53124_ (_01515_, _01317_, _31338_);
  or _53125_ (_01516_, _01515_, _01514_);
  and _53126_ (_39716_, _01516_, _41806_);
  and _53127_ (_01517_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _53128_ (_01518_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or _53129_ (_01519_, _01518_, _01517_);
  and _53130_ (_01520_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _53131_ (_01521_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _53132_ (_01522_, _01521_, _01520_);
  or _53133_ (_01523_, _01522_, _01519_);
  and _53134_ (_01524_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _53135_ (_01525_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _53136_ (_01526_, _01525_, _01524_);
  and _53137_ (_01527_, _01339_, _40511_);
  and _53138_ (_01528_, _01341_, _01016_);
  or _53139_ (_01530_, _01528_, _01527_);
  or _53140_ (_01531_, _01530_, _01526_);
  or _53141_ (_01533_, _01531_, _01523_);
  and _53142_ (_01534_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _53143_ (_01535_, _01347_, _00896_);
  and _53144_ (_01537_, _01350_, _01130_);
  or _53145_ (_01538_, _01537_, _01535_);
  and _53146_ (_01539_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _53147_ (_01541_, _01354_, _01166_);
  or _53148_ (_01542_, _01541_, _01539_);
  or _53149_ (_01543_, _01542_, _01538_);
  or _53150_ (_01545_, _01543_, _01534_);
  or _53151_ (_01546_, _01545_, _01533_);
  and _53152_ (_01547_, _01546_, _01312_);
  nor _53153_ (_01549_, _01312_, _16172_);
  or _53154_ (_01550_, _01549_, _01547_);
  and _53155_ (_01551_, _01550_, _01317_);
  nor _53156_ (_01553_, _01317_, _32044_);
  or _53157_ (_01554_, _01553_, _01551_);
  and _53158_ (_39717_, _01554_, _41806_);
  and _53159_ (_01556_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _53160_ (_01557_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or _53161_ (_01558_, _01557_, _01556_);
  and _53162_ (_01560_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _53163_ (_01561_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _53164_ (_01562_, _01561_, _01560_);
  or _53165_ (_01563_, _01562_, _01558_);
  and _53166_ (_01564_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _53167_ (_01565_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _53168_ (_01566_, _01565_, _01564_);
  and _53169_ (_01567_, _01339_, _40427_);
  and _53170_ (_01568_, _01341_, _01056_);
  or _53171_ (_01569_, _01568_, _01567_);
  or _53172_ (_01570_, _01569_, _01566_);
  or _53173_ (_01571_, _01570_, _01563_);
  and _53174_ (_01572_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _53175_ (_01573_, _01347_, _00937_);
  and _53176_ (_01574_, _01350_, _01080_);
  or _53177_ (_01575_, _01574_, _01573_);
  and _53178_ (_01576_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _53179_ (_01577_, _01354_, _01150_);
  or _53180_ (_01578_, _01577_, _01576_);
  or _53181_ (_01579_, _01578_, _01575_);
  or _53182_ (_01580_, _01579_, _01572_);
  or _53183_ (_01582_, _01580_, _01571_);
  and _53184_ (_01583_, _01582_, _01312_);
  nor _53185_ (_01585_, _01312_, _17160_);
  or _53186_ (_01586_, _01585_, _01583_);
  and _53187_ (_01587_, _01586_, _01317_);
  nor _53188_ (_01589_, _01317_, _32853_);
  or _53189_ (_01590_, _01589_, _01587_);
  and _53190_ (_39718_, _01590_, _41806_);
  and _53191_ (_01592_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _53192_ (_01593_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _53193_ (_01594_, _01593_, _01592_);
  and _53194_ (_01596_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _53195_ (_01597_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _53196_ (_01598_, _01597_, _01596_);
  or _53197_ (_01600_, _01598_, _01594_);
  and _53198_ (_01601_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _53199_ (_01602_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _53200_ (_01604_, _01602_, _01601_);
  and _53201_ (_01605_, _01339_, _40695_);
  and _53202_ (_01606_, _01341_, _01007_);
  or _53203_ (_01608_, _01606_, _01605_);
  or _53204_ (_01609_, _01608_, _01604_);
  or _53205_ (_01610_, _01609_, _01600_);
  and _53206_ (_01612_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _53207_ (_01613_, _01347_, _00885_);
  and _53208_ (_01614_, _01350_, _01114_);
  or _53209_ (_01615_, _01614_, _01613_);
  and _53210_ (_01616_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _53211_ (_01617_, _01354_, _01183_);
  or _53212_ (_01618_, _01617_, _01616_);
  or _53213_ (_01619_, _01618_, _01615_);
  or _53214_ (_01620_, _01619_, _01612_);
  or _53215_ (_01621_, _01620_, _01610_);
  and _53216_ (_01622_, _01621_, _01312_);
  nor _53217_ (_01623_, _01312_, _16512_);
  or _53218_ (_01624_, _01623_, _01622_);
  and _53219_ (_01625_, _01624_, _01317_);
  nor _53220_ (_01626_, _01317_, _33598_);
  or _53221_ (_01627_, _01626_, _01625_);
  and _53222_ (_39719_, _01627_, _41806_);
  and _53223_ (_39764_, _40734_, _41806_);
  and _53224_ (_39765_, _40870_, _41806_);
  nor _53225_ (_39767_, _40500_, rst);
  and _53226_ (_39783_, _40888_, _41806_);
  and _53227_ (_39784_, _40901_, _41806_);
  and _53228_ (_39785_, _40914_, _41806_);
  and _53229_ (_39786_, _40922_, _41806_);
  and _53230_ (_39787_, _40932_, _41806_);
  and _53231_ (_39788_, _40942_, _41806_);
  and _53232_ (_39789_, _40952_, _41806_);
  nor _53233_ (_39790_, _40415_, rst);
  nor _53234_ (_39791_, _40611_, rst);
  not _53235_ (_01632_, _41697_);
  nor _53236_ (_01633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _53237_ (_01635_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53238_ (_01636_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01635_);
  nor _53239_ (_01637_, _01636_, _01633_);
  nor _53240_ (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53241_ (_01640_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01635_);
  nor _53242_ (_01641_, _01640_, _01639_);
  not _53243_ (_01643_, _01641_);
  nor _53244_ (_01644_, _01643_, _01637_);
  nor _53245_ (_01645_, _00129_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53246_ (_01647_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01635_);
  nor _53247_ (_01648_, _01647_, _01645_);
  not _53248_ (_01649_, _01648_);
  nor _53249_ (_01651_, _01641_, _01637_);
  not _53250_ (_01652_, _01651_);
  nor _53251_ (_01653_, _00110_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53252_ (_01654_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01635_);
  nor _53253_ (_01655_, _01654_, _01653_);
  and _53254_ (_01656_, _01655_, _01652_);
  or _53255_ (_01657_, _01656_, _01649_);
  nor _53256_ (_01658_, _01655_, _01652_);
  or _53257_ (_01659_, _01658_, _01648_);
  and _53258_ (_01660_, _01659_, _01657_);
  and _53259_ (_01661_, _01660_, _01644_);
  and _53260_ (_01662_, _01661_, _01632_);
  not _53261_ (_01663_, _41738_);
  and _53262_ (_01664_, _01641_, _01637_);
  and _53263_ (_01665_, _01660_, _01664_);
  and _53264_ (_01666_, _01665_, _01663_);
  or _53265_ (_01667_, _01666_, _01662_);
  not _53266_ (_01668_, _41656_);
  and _53267_ (_01669_, _01643_, _01637_);
  and _53268_ (_01670_, _01669_, _01660_);
  and _53269_ (_01671_, _01670_, _01668_);
  not _53270_ (_01673_, _42040_);
  and _53271_ (_01674_, _01649_, _01655_);
  and _53272_ (_01676_, _01674_, _01644_);
  and _53273_ (_01677_, _01676_, _01673_);
  not _53274_ (_01678_, _42081_);
  and _53275_ (_01680_, _01674_, _01664_);
  and _53276_ (_01681_, _01680_, _01678_);
  or _53277_ (_01682_, _01681_, _01677_);
  not _53278_ (_01684_, _41999_);
  and _53279_ (_01685_, _01669_, _01674_);
  and _53280_ (_01686_, _01685_, _01684_);
  not _53281_ (_01688_, _41786_);
  and _53282_ (_01689_, _01658_, _01649_);
  and _53283_ (_01690_, _01689_, _01688_);
  or _53284_ (_01692_, _01690_, _01686_);
  or _53285_ (_01693_, _01692_, _01682_);
  or _53286_ (_01694_, _01693_, _01671_);
  or _53287_ (_01696_, _01694_, _01667_);
  not _53288_ (_01697_, _41917_);
  nor _53289_ (_01698_, _01658_, _01656_);
  and _53290_ (_01700_, _01698_, _01649_);
  and _53291_ (_01701_, _01700_, _01664_);
  and _53292_ (_01702_, _01701_, _01697_);
  not _53293_ (_01704_, _42204_);
  and _53294_ (_01705_, _01698_, _01648_);
  and _53295_ (_01706_, _01705_, _01644_);
  and _53296_ (_01707_, _01706_, _01704_);
  not _53297_ (_01708_, _42163_);
  and _53298_ (_01709_, _01705_, _01669_);
  and _53299_ (_01710_, _01709_, _01708_);
  or _53300_ (_01711_, _01710_, _01707_);
  or _53301_ (_01712_, _01711_, _01702_);
  not _53302_ (_01713_, _41876_);
  and _53303_ (_01714_, _01700_, _01644_);
  and _53304_ (_01715_, _01714_, _01713_);
  not _53305_ (_01716_, _41958_);
  and _53306_ (_01717_, _01674_, _01651_);
  and _53307_ (_01718_, _01717_, _01716_);
  not _53308_ (_01719_, _42286_);
  and _53309_ (_01720_, _01655_, _01651_);
  and _53310_ (_01721_, _01720_, _01648_);
  and _53311_ (_01722_, _01721_, _01719_);
  not _53312_ (_01723_, _42122_);
  and _53313_ (_01724_, _01658_, _01648_);
  and _53314_ (_01726_, _01724_, _01723_);
  or _53315_ (_01727_, _01726_, _01722_);
  or _53316_ (_01729_, _01727_, _01718_);
  or _53317_ (_01730_, _01729_, _01715_);
  not _53318_ (_01731_, _42245_);
  and _53319_ (_01733_, _01705_, _01664_);
  and _53320_ (_01734_, _01733_, _01731_);
  not _53321_ (_01735_, _41835_);
  and _53322_ (_01737_, _01700_, _01669_);
  and _53323_ (_01738_, _01737_, _01735_);
  or _53324_ (_01739_, _01738_, _01734_);
  or _53325_ (_01741_, _01739_, _01730_);
  or _53326_ (_01742_, _01741_, _01712_);
  or _53327_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01742_, _01696_);
  and _53328_ (_01744_, _01661_, _01719_);
  and _53329_ (_01745_, _01680_, _01684_);
  and _53330_ (_01746_, _01676_, _01716_);
  or _53331_ (_01748_, _01746_, _01745_);
  and _53332_ (_01749_, _01689_, _01632_);
  and _53333_ (_01750_, _01685_, _01697_);
  or _53334_ (_01752_, _01750_, _01749_);
  or _53335_ (_01753_, _01752_, _01748_);
  or _53336_ (_01754_, _01753_, _01744_);
  and _53337_ (_01756_, _01665_, _01668_);
  and _53338_ (_01757_, _01670_, _01731_);
  or _53339_ (_01758_, _01757_, _01756_);
  or _53340_ (_01759_, _01758_, _01754_);
  and _53341_ (_01760_, _01737_, _01663_);
  and _53342_ (_01761_, _01714_, _01688_);
  and _53343_ (_01762_, _01706_, _01723_);
  or _53344_ (_01763_, _01762_, _01761_);
  or _53345_ (_01764_, _01763_, _01760_);
  and _53346_ (_01765_, _01709_, _01678_);
  and _53347_ (_01766_, _01717_, _01713_);
  and _53348_ (_01767_, _01724_, _01673_);
  and _53349_ (_01768_, _01721_, _01704_);
  or _53350_ (_01769_, _01768_, _01767_);
  or _53351_ (_01770_, _01769_, _01766_);
  or _53352_ (_01771_, _01770_, _01765_);
  and _53353_ (_01772_, _01701_, _01735_);
  and _53354_ (_01773_, _01733_, _01708_);
  or _53355_ (_01774_, _01773_, _01772_);
  or _53356_ (_01775_, _01774_, _01771_);
  or _53357_ (_01776_, _01775_, _01764_);
  or _53358_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01776_, _01759_);
  and _53359_ (_01778_, _01665_, _01632_);
  and _53360_ (_01780_, _01717_, _01697_);
  and _53361_ (_01781_, _01676_, _01684_);
  or _53362_ (_01782_, _01781_, _01780_);
  and _53363_ (_01784_, _01689_, _01663_);
  and _53364_ (_01785_, _01680_, _01673_);
  or _53365_ (_01786_, _01785_, _01784_);
  or _53366_ (_01788_, _01786_, _01782_);
  or _53367_ (_01789_, _01788_, _01778_);
  and _53368_ (_01790_, _01670_, _01719_);
  and _53369_ (_01792_, _01661_, _01668_);
  or _53370_ (_01793_, _01792_, _01790_);
  or _53371_ (_01794_, _01793_, _01789_);
  and _53372_ (_01796_, _01714_, _01735_);
  and _53373_ (_01797_, _01701_, _01713_);
  and _53374_ (_01798_, _01709_, _01723_);
  or _53375_ (_01800_, _01798_, _01797_);
  or _53376_ (_01801_, _01800_, _01796_);
  and _53377_ (_01802_, _01737_, _01688_);
  and _53378_ (_01804_, _01685_, _01716_);
  and _53379_ (_01805_, _01724_, _01678_);
  and _53380_ (_01806_, _01721_, _01731_);
  or _53381_ (_01808_, _01806_, _01805_);
  or _53382_ (_01809_, _01808_, _01804_);
  or _53383_ (_01810_, _01809_, _01802_);
  and _53384_ (_01811_, _01733_, _01704_);
  and _53385_ (_01812_, _01706_, _01708_);
  or _53386_ (_01813_, _01812_, _01811_);
  or _53387_ (_01814_, _01813_, _01810_);
  or _53388_ (_01815_, _01814_, _01801_);
  or _53389_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01815_, _01794_);
  and _53390_ (_01816_, _01665_, _01719_);
  and _53391_ (_01817_, _01661_, _01731_);
  or _53392_ (_01818_, _01817_, _01816_);
  and _53393_ (_01819_, _01670_, _01704_);
  and _53394_ (_01820_, _01676_, _01697_);
  and _53395_ (_01821_, _01685_, _01713_);
  or _53396_ (_01822_, _01821_, _01820_);
  and _53397_ (_01823_, _01689_, _01668_);
  and _53398_ (_01824_, _01717_, _01735_);
  or _53399_ (_01825_, _01824_, _01823_);
  or _53400_ (_01826_, _01825_, _01822_);
  or _53401_ (_01827_, _01826_, _01819_);
  or _53402_ (_01829_, _01827_, _01818_);
  and _53403_ (_01830_, _01714_, _01663_);
  and _53404_ (_01832_, _01733_, _01723_);
  and _53405_ (_01833_, _01737_, _01632_);
  or _53406_ (_01834_, _01833_, _01832_);
  or _53407_ (_01836_, _01834_, _01830_);
  and _53408_ (_01837_, _01709_, _01673_);
  and _53409_ (_01838_, _01680_, _01716_);
  and _53410_ (_01840_, _01721_, _01708_);
  and _53411_ (_01841_, _01724_, _01684_);
  or _53412_ (_01842_, _01841_, _01840_);
  or _53413_ (_01844_, _01842_, _01838_);
  or _53414_ (_01845_, _01844_, _01837_);
  and _53415_ (_01846_, _01706_, _01678_);
  and _53416_ (_01848_, _01701_, _01688_);
  or _53417_ (_01849_, _01848_, _01846_);
  or _53418_ (_01850_, _01849_, _01845_);
  or _53419_ (_01852_, _01850_, _01836_);
  or _53420_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01852_, _01829_);
  not _53421_ (_01853_, _41743_);
  and _53422_ (_01855_, _01665_, _01853_);
  not _53423_ (_01856_, _41791_);
  and _53424_ (_01857_, _01689_, _01856_);
  not _53425_ (_01859_, _42086_);
  and _53426_ (_01860_, _01680_, _01859_);
  or _53427_ (_01861_, _01860_, _01857_);
  not _53428_ (_01862_, _42045_);
  and _53429_ (_01863_, _01676_, _01862_);
  not _53430_ (_01864_, _42004_);
  and _53431_ (_01865_, _01685_, _01864_);
  or _53432_ (_01866_, _01865_, _01863_);
  or _53433_ (_01867_, _01866_, _01861_);
  or _53434_ (_01868_, _01867_, _01855_);
  not _53435_ (_01869_, _41661_);
  and _53436_ (_01870_, _01670_, _01869_);
  not _53437_ (_01871_, _41702_);
  and _53438_ (_01872_, _01661_, _01871_);
  or _53439_ (_01873_, _01872_, _01870_);
  or _53440_ (_01874_, _01873_, _01868_);
  not _53441_ (_01875_, _42168_);
  and _53442_ (_01876_, _01709_, _01875_);
  not _53443_ (_01877_, _41922_);
  and _53444_ (_01878_, _01701_, _01877_);
  not _53445_ (_01879_, _42209_);
  and _53446_ (_01881_, _01706_, _01879_);
  or _53447_ (_01882_, _01881_, _01878_);
  or _53448_ (_01884_, _01882_, _01876_);
  not _53449_ (_01885_, _41881_);
  and _53450_ (_01886_, _01714_, _01885_);
  not _53451_ (_01888_, _41963_);
  and _53452_ (_01889_, _01717_, _01888_);
  not _53453_ (_01890_, _42291_);
  and _53454_ (_01892_, _01721_, _01890_);
  not _53455_ (_01893_, _42127_);
  and _53456_ (_01894_, _01724_, _01893_);
  or _53457_ (_01896_, _01894_, _01892_);
  or _53458_ (_01897_, _01896_, _01889_);
  or _53459_ (_01898_, _01897_, _01886_);
  not _53460_ (_01900_, _41840_);
  and _53461_ (_01901_, _01737_, _01900_);
  not _53462_ (_01902_, _42250_);
  and _53463_ (_01904_, _01733_, _01902_);
  or _53464_ (_01905_, _01904_, _01901_);
  or _53465_ (_01906_, _01905_, _01898_);
  or _53466_ (_01908_, _01906_, _01884_);
  or _53467_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01908_, _01874_);
  not _53468_ (_01909_, _41749_);
  and _53469_ (_01911_, _01665_, _01909_);
  not _53470_ (_01912_, _42050_);
  and _53471_ (_01913_, _01676_, _01912_);
  not _53472_ (_01914_, _42091_);
  and _53473_ (_01915_, _01680_, _01914_);
  or _53474_ (_01916_, _01915_, _01913_);
  not _53475_ (_01917_, _41968_);
  and _53476_ (_01918_, _01717_, _01917_);
  not _53477_ (_01919_, _42009_);
  and _53478_ (_01920_, _01685_, _01919_);
  or _53479_ (_01921_, _01920_, _01918_);
  or _53480_ (_01922_, _01921_, _01916_);
  or _53481_ (_01923_, _01922_, _01911_);
  not _53482_ (_01924_, _41666_);
  and _53483_ (_01925_, _01670_, _01924_);
  not _53484_ (_01926_, _41707_);
  and _53485_ (_01927_, _01661_, _01926_);
  or _53486_ (_01928_, _01927_, _01925_);
  or _53487_ (_01929_, _01928_, _01923_);
  not _53488_ (_01930_, _41886_);
  and _53489_ (_01931_, _01714_, _01930_);
  not _53490_ (_01933_, _41927_);
  and _53491_ (_01934_, _01701_, _01933_);
  or _53492_ (_01936_, _01934_, _01931_);
  not _53493_ (_01937_, _42214_);
  and _53494_ (_01938_, _01706_, _01937_);
  or _53495_ (_01940_, _01938_, _01936_);
  not _53496_ (_01941_, _42173_);
  and _53497_ (_01942_, _01709_, _01941_);
  not _53498_ (_01944_, _41801_);
  and _53499_ (_01945_, _01689_, _01944_);
  not _53500_ (_01946_, _42296_);
  and _53501_ (_01948_, _01721_, _01946_);
  not _53502_ (_01949_, _42132_);
  and _53503_ (_01950_, _01724_, _01949_);
  or _53504_ (_01952_, _01950_, _01948_);
  or _53505_ (_01953_, _01952_, _01945_);
  or _53506_ (_01954_, _01953_, _01942_);
  not _53507_ (_01956_, _41845_);
  and _53508_ (_01957_, _01737_, _01956_);
  not _53509_ (_01958_, _42255_);
  and _53510_ (_01960_, _01733_, _01958_);
  or _53511_ (_01961_, _01960_, _01957_);
  or _53512_ (_01962_, _01961_, _01954_);
  or _53513_ (_01964_, _01962_, _01940_);
  or _53514_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01964_, _01929_);
  not _53515_ (_01965_, _41671_);
  and _53516_ (_01966_, _01670_, _01965_);
  not _53517_ (_01967_, _41758_);
  and _53518_ (_01968_, _01665_, _01967_);
  or _53519_ (_01969_, _01968_, _01966_);
  not _53520_ (_01970_, _41712_);
  and _53521_ (_01971_, _01661_, _01970_);
  not _53522_ (_01972_, _42096_);
  and _53523_ (_01973_, _01680_, _01972_);
  not _53524_ (_01974_, _42055_);
  and _53525_ (_01975_, _01676_, _01974_);
  or _53526_ (_01976_, _01975_, _01973_);
  not _53527_ (_01977_, _41973_);
  and _53528_ (_01978_, _01717_, _01977_);
  not _53529_ (_01979_, _41809_);
  and _53530_ (_01980_, _01689_, _01979_);
  or _53531_ (_01981_, _01980_, _01978_);
  or _53532_ (_01982_, _01981_, _01976_);
  or _53533_ (_01983_, _01982_, _01971_);
  or _53534_ (_01985_, _01983_, _01969_);
  not _53535_ (_01986_, _41891_);
  and _53536_ (_01988_, _01714_, _01986_);
  not _53537_ (_01989_, _42260_);
  and _53538_ (_01990_, _01733_, _01989_);
  not _53539_ (_01992_, _41932_);
  and _53540_ (_01993_, _01701_, _01992_);
  or _53541_ (_01994_, _01993_, _01990_);
  or _53542_ (_01996_, _01994_, _01988_);
  not _53543_ (_01997_, _42219_);
  and _53544_ (_01998_, _01706_, _01997_);
  not _53545_ (_02000_, _42014_);
  and _53546_ (_02001_, _01685_, _02000_);
  not _53547_ (_02002_, _42301_);
  and _53548_ (_02004_, _01721_, _02002_);
  not _53549_ (_02005_, _42137_);
  and _53550_ (_02006_, _01724_, _02005_);
  or _53551_ (_02008_, _02006_, _02004_);
  or _53552_ (_02009_, _02008_, _02001_);
  or _53553_ (_02010_, _02009_, _01998_);
  not _53554_ (_02012_, _42178_);
  and _53555_ (_02013_, _01709_, _02012_);
  not _53556_ (_02014_, _41850_);
  and _53557_ (_02016_, _01737_, _02014_);
  or _53558_ (_02017_, _02016_, _02013_);
  or _53559_ (_02018_, _02017_, _02010_);
  or _53560_ (_02019_, _02018_, _01996_);
  or _53561_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _02019_, _01985_);
  not _53562_ (_02020_, _41676_);
  and _53563_ (_02021_, _01670_, _02020_);
  not _53564_ (_02022_, _41765_);
  and _53565_ (_02023_, _01665_, _02022_);
  or _53566_ (_02024_, _02023_, _02021_);
  not _53567_ (_02025_, _41978_);
  and _53568_ (_02026_, _01717_, _02025_);
  not _53569_ (_02027_, _42019_);
  and _53570_ (_02028_, _01685_, _02027_);
  or _53571_ (_02029_, _02028_, _02026_);
  not _53572_ (_02030_, _42101_);
  and _53573_ (_02031_, _01680_, _02030_);
  not _53574_ (_02032_, _42060_);
  and _53575_ (_02033_, _01676_, _02032_);
  or _53576_ (_02034_, _02033_, _02031_);
  or _53577_ (_02035_, _02034_, _02029_);
  not _53578_ (_02037_, _41717_);
  and _53579_ (_02038_, _01661_, _02037_);
  or _53580_ (_02040_, _02038_, _02035_);
  or _53581_ (_02041_, _02040_, _02024_);
  not _53582_ (_02042_, _41937_);
  and _53583_ (_02044_, _01701_, _02042_);
  not _53584_ (_02045_, _42224_);
  and _53585_ (_02046_, _01706_, _02045_);
  not _53586_ (_02048_, _41896_);
  and _53587_ (_02049_, _01714_, _02048_);
  or _53588_ (_02050_, _02049_, _02046_);
  or _53589_ (_02052_, _02050_, _02044_);
  not _53590_ (_02053_, _41855_);
  and _53591_ (_02054_, _01737_, _02053_);
  not _53592_ (_02056_, _41814_);
  and _53593_ (_02057_, _01689_, _02056_);
  not _53594_ (_02058_, _42306_);
  and _53595_ (_02060_, _01721_, _02058_);
  not _53596_ (_02061_, _42142_);
  and _53597_ (_02062_, _01724_, _02061_);
  or _53598_ (_02064_, _02062_, _02060_);
  or _53599_ (_02065_, _02064_, _02057_);
  or _53600_ (_02066_, _02065_, _02054_);
  not _53601_ (_02068_, _42265_);
  and _53602_ (_02069_, _01733_, _02068_);
  not _53603_ (_02070_, _42183_);
  and _53604_ (_02071_, _01709_, _02070_);
  or _53605_ (_02072_, _02071_, _02069_);
  or _53606_ (_02073_, _02072_, _02066_);
  or _53607_ (_02074_, _02073_, _02052_);
  or _53608_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _02074_, _02041_);
  not _53609_ (_02075_, _41681_);
  and _53610_ (_02076_, _01670_, _02075_);
  not _53611_ (_02077_, _41770_);
  and _53612_ (_02078_, _01665_, _02077_);
  or _53613_ (_02079_, _02078_, _02076_);
  not _53614_ (_02080_, _41722_);
  and _53615_ (_02081_, _01661_, _02080_);
  not _53616_ (_02082_, _42065_);
  and _53617_ (_02083_, _01676_, _02082_);
  not _53618_ (_02084_, _42106_);
  and _53619_ (_02085_, _01680_, _02084_);
  or _53620_ (_02086_, _02085_, _02083_);
  not _53621_ (_02087_, _41983_);
  and _53622_ (_02089_, _01717_, _02087_);
  not _53623_ (_02090_, _42024_);
  and _53624_ (_02092_, _01685_, _02090_);
  or _53625_ (_02093_, _02092_, _02089_);
  or _53626_ (_02094_, _02093_, _02086_);
  or _53627_ (_02096_, _02094_, _02081_);
  or _53628_ (_02097_, _02096_, _02079_);
  not _53629_ (_02098_, _42270_);
  and _53630_ (_02100_, _01733_, _02098_);
  not _53631_ (_02101_, _41901_);
  and _53632_ (_02102_, _01714_, _02101_);
  not _53633_ (_02104_, _42229_);
  and _53634_ (_02105_, _01706_, _02104_);
  or _53635_ (_02106_, _02105_, _02102_);
  or _53636_ (_02108_, _02106_, _02100_);
  not _53637_ (_02109_, _42188_);
  and _53638_ (_02110_, _01709_, _02109_);
  not _53639_ (_02112_, _41819_);
  and _53640_ (_02113_, _01689_, _02112_);
  not _53641_ (_02114_, _42311_);
  and _53642_ (_02116_, _01721_, _02114_);
  not _53643_ (_02117_, _42147_);
  and _53644_ (_02118_, _01724_, _02117_);
  or _53645_ (_02120_, _02118_, _02116_);
  or _53646_ (_02121_, _02120_, _02113_);
  or _53647_ (_02122_, _02121_, _02110_);
  not _53648_ (_02123_, _41942_);
  and _53649_ (_02124_, _01701_, _02123_);
  not _53650_ (_02125_, _41860_);
  and _53651_ (_02126_, _01737_, _02125_);
  or _53652_ (_02127_, _02126_, _02124_);
  or _53653_ (_02128_, _02127_, _02122_);
  or _53654_ (_02129_, _02128_, _02108_);
  or _53655_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _02129_, _02097_);
  not _53656_ (_02130_, _41727_);
  and _53657_ (_02131_, _01661_, _02130_);
  not _53658_ (_02132_, _41775_);
  and _53659_ (_02133_, _01665_, _02132_);
  or _53660_ (_02134_, _02133_, _02131_);
  not _53661_ (_02135_, _41686_);
  and _53662_ (_02136_, _01670_, _02135_);
  not _53663_ (_02137_, _42111_);
  and _53664_ (_02138_, _01680_, _02137_);
  not _53665_ (_02139_, _41824_);
  and _53666_ (_02141_, _01689_, _02139_);
  or _53667_ (_02142_, _02141_, _02138_);
  not _53668_ (_02144_, _42070_);
  and _53669_ (_02145_, _01676_, _02144_);
  not _53670_ (_02146_, _41988_);
  and _53671_ (_02148_, _01717_, _02146_);
  or _53672_ (_02149_, _02148_, _02145_);
  or _53673_ (_02150_, _02149_, _02142_);
  or _53674_ (_02152_, _02150_, _02136_);
  or _53675_ (_02153_, _02152_, _02134_);
  not _53676_ (_02154_, _42275_);
  and _53677_ (_02156_, _01733_, _02154_);
  not _53678_ (_02157_, _42193_);
  and _53679_ (_02158_, _01709_, _02157_);
  not _53680_ (_02160_, _41947_);
  and _53681_ (_02161_, _01701_, _02160_);
  or _53682_ (_02162_, _02161_, _02158_);
  or _53683_ (_02164_, _02162_, _02156_);
  not _53684_ (_02165_, _42234_);
  and _53685_ (_02166_, _01706_, _02165_);
  not _53686_ (_02168_, _42029_);
  and _53687_ (_02169_, _01685_, _02168_);
  not _53688_ (_02170_, _42316_);
  and _53689_ (_02172_, _01721_, _02170_);
  not _53690_ (_02173_, _42152_);
  and _53691_ (_02174_, _01724_, _02173_);
  or _53692_ (_02175_, _02174_, _02172_);
  or _53693_ (_02176_, _02175_, _02169_);
  or _53694_ (_02177_, _02176_, _02166_);
  not _53695_ (_02178_, _41906_);
  and _53696_ (_02179_, _01714_, _02178_);
  not _53697_ (_02180_, _41865_);
  and _53698_ (_02181_, _01737_, _02180_);
  or _53699_ (_02182_, _02181_, _02179_);
  or _53700_ (_02183_, _02182_, _02177_);
  or _53701_ (_02184_, _02183_, _02164_);
  or _53702_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _02184_, _02153_);
  not _53703_ (_02185_, _41691_);
  and _53704_ (_02186_, _01670_, _02185_);
  not _53705_ (_02187_, _41780_);
  and _53706_ (_02188_, _01665_, _02187_);
  or _53707_ (_02189_, _02188_, _02186_);
  not _53708_ (_02190_, _41732_);
  and _53709_ (_02191_, _01661_, _02190_);
  not _53710_ (_02193_, _42116_);
  and _53711_ (_02194_, _01680_, _02193_);
  not _53712_ (_02196_, _42075_);
  and _53713_ (_02197_, _01676_, _02196_);
  or _53714_ (_02198_, _02197_, _02194_);
  not _53715_ (_02200_, _42034_);
  and _53716_ (_02201_, _01685_, _02200_);
  not _53717_ (_02202_, _41829_);
  and _53718_ (_02204_, _01689_, _02202_);
  or _53719_ (_02205_, _02204_, _02201_);
  or _53720_ (_02206_, _02205_, _02198_);
  or _53721_ (_02208_, _02206_, _02191_);
  or _53722_ (_02209_, _02208_, _02189_);
  not _53723_ (_02210_, _41952_);
  and _53724_ (_02212_, _01701_, _02210_);
  not _53725_ (_02213_, _41911_);
  and _53726_ (_02214_, _01714_, _02213_);
  or _53727_ (_02216_, _02214_, _02212_);
  not _53728_ (_02217_, _41870_);
  and _53729_ (_02218_, _01737_, _02217_);
  or _53730_ (_02220_, _02218_, _02216_);
  not _53731_ (_02221_, _42280_);
  and _53732_ (_02222_, _01733_, _02221_);
  not _53733_ (_02224_, _41993_);
  and _53734_ (_02225_, _01717_, _02224_);
  not _53735_ (_02226_, _42321_);
  and _53736_ (_02227_, _01721_, _02226_);
  not _53737_ (_02228_, _42157_);
  and _53738_ (_02229_, _01724_, _02228_);
  or _53739_ (_02230_, _02229_, _02227_);
  or _53740_ (_02231_, _02230_, _02225_);
  or _53741_ (_02232_, _02231_, _02222_);
  not _53742_ (_02233_, _42239_);
  and _53743_ (_02234_, _01706_, _02233_);
  not _53744_ (_02235_, _42198_);
  and _53745_ (_02236_, _01709_, _02235_);
  or _53746_ (_02237_, _02236_, _02234_);
  or _53747_ (_02238_, _02237_, _02232_);
  or _53748_ (_02239_, _02238_, _02220_);
  or _53749_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _02239_, _02209_);
  and _53750_ (_02240_, _01665_, _01871_);
  and _53751_ (_02241_, _01680_, _01862_);
  and _53752_ (_02242_, _01685_, _01888_);
  or _53753_ (_02243_, _02242_, _02241_);
  and _53754_ (_02244_, _01689_, _01853_);
  and _53755_ (_02245_, _01676_, _01864_);
  or _53756_ (_02246_, _02245_, _02244_);
  or _53757_ (_02247_, _02246_, _02243_);
  or _53758_ (_02248_, _02247_, _02240_);
  and _53759_ (_02249_, _01670_, _01890_);
  and _53760_ (_02250_, _01661_, _01869_);
  or _53761_ (_02251_, _02250_, _02249_);
  or _53762_ (_02252_, _02251_, _02248_);
  and _53763_ (_02253_, _01709_, _01893_);
  and _53764_ (_02254_, _01714_, _01900_);
  and _53765_ (_02255_, _01706_, _01875_);
  or _53766_ (_02256_, _02255_, _02254_);
  or _53767_ (_02257_, _02256_, _02253_);
  and _53768_ (_02258_, _01737_, _01856_);
  and _53769_ (_02259_, _01717_, _01877_);
  and _53770_ (_02260_, _01724_, _01859_);
  and _53771_ (_02261_, _01721_, _01902_);
  or _53772_ (_02262_, _02261_, _02260_);
  or _53773_ (_02263_, _02262_, _02259_);
  or _53774_ (_02264_, _02263_, _02258_);
  and _53775_ (_02265_, _01701_, _01885_);
  and _53776_ (_02266_, _01733_, _01879_);
  or _53777_ (_02267_, _02266_, _02265_);
  or _53778_ (_02268_, _02267_, _02264_);
  or _53779_ (_02269_, _02268_, _02257_);
  or _53780_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _02269_, _02252_);
  and _53781_ (_02270_, _01665_, _01926_);
  and _53782_ (_02271_, _01689_, _01909_);
  and _53783_ (_02272_, _01680_, _01912_);
  or _53784_ (_02273_, _02272_, _02271_);
  and _53785_ (_02274_, _01717_, _01933_);
  and _53786_ (_02275_, _01676_, _01919_);
  or _53787_ (_02276_, _02275_, _02274_);
  or _53788_ (_02277_, _02276_, _02273_);
  or _53789_ (_02278_, _02277_, _02270_);
  and _53790_ (_02279_, _01670_, _01946_);
  and _53791_ (_02280_, _01661_, _01924_);
  or _53792_ (_02281_, _02280_, _02279_);
  or _53793_ (_02282_, _02281_, _02278_);
  and _53794_ (_02283_, _01706_, _01941_);
  and _53795_ (_02284_, _01714_, _01956_);
  and _53796_ (_02285_, _01733_, _01937_);
  or _53797_ (_02286_, _02285_, _02284_);
  or _53798_ (_02287_, _02286_, _02283_);
  and _53799_ (_02288_, _01737_, _01944_);
  and _53800_ (_02289_, _01685_, _01917_);
  and _53801_ (_02290_, _01724_, _01914_);
  and _53802_ (_02291_, _01721_, _01958_);
  or _53803_ (_02292_, _02291_, _02290_);
  or _53804_ (_02293_, _02292_, _02289_);
  or _53805_ (_02294_, _02293_, _02288_);
  and _53806_ (_02295_, _01701_, _01930_);
  and _53807_ (_02296_, _01709_, _01949_);
  or _53808_ (_02297_, _02296_, _02295_);
  or _53809_ (_02298_, _02297_, _02294_);
  or _53810_ (_02299_, _02298_, _02287_);
  or _53811_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02299_, _02282_);
  and _53812_ (_02300_, _01661_, _01965_);
  and _53813_ (_02301_, _01689_, _01967_);
  and _53814_ (_02302_, _01685_, _01977_);
  or _53815_ (_02303_, _02302_, _02301_);
  and _53816_ (_02304_, _01680_, _01974_);
  and _53817_ (_02305_, _01676_, _02000_);
  or _53818_ (_02306_, _02305_, _02304_);
  or _53819_ (_02307_, _02306_, _02303_);
  or _53820_ (_02308_, _02307_, _02300_);
  and _53821_ (_02309_, _01670_, _02002_);
  and _53822_ (_02310_, _01665_, _01970_);
  or _53823_ (_02311_, _02310_, _02309_);
  or _53824_ (_02312_, _02311_, _02308_);
  and _53825_ (_02313_, _01714_, _02014_);
  and _53826_ (_02314_, _01737_, _01979_);
  or _53827_ (_02315_, _02314_, _02313_);
  and _53828_ (_02316_, _01701_, _01986_);
  or _53829_ (_02317_, _02316_, _02315_);
  and _53830_ (_02318_, _01709_, _02005_);
  and _53831_ (_02319_, _01717_, _01992_);
  and _53832_ (_02320_, _01724_, _01972_);
  and _53833_ (_02321_, _01721_, _01989_);
  or _53834_ (_02322_, _02321_, _02320_);
  or _53835_ (_02323_, _02322_, _02319_);
  or _53836_ (_02324_, _02323_, _02318_);
  and _53837_ (_02325_, _01733_, _01997_);
  and _53838_ (_02326_, _01706_, _02012_);
  or _53839_ (_02327_, _02326_, _02325_);
  or _53840_ (_02328_, _02327_, _02324_);
  or _53841_ (_02329_, _02328_, _02317_);
  or _53842_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02329_, _02312_);
  and _53843_ (_02330_, _01665_, _02037_);
  and _53844_ (_02331_, _01685_, _02025_);
  and _53845_ (_02332_, _01717_, _02042_);
  or _53846_ (_02333_, _02332_, _02331_);
  and _53847_ (_02334_, _01680_, _02032_);
  and _53848_ (_02335_, _01676_, _02027_);
  or _53849_ (_02336_, _02335_, _02334_);
  or _53850_ (_02337_, _02336_, _02333_);
  or _53851_ (_02338_, _02337_, _02330_);
  and _53852_ (_02339_, _01670_, _02058_);
  and _53853_ (_02340_, _01661_, _02020_);
  or _53854_ (_02341_, _02340_, _02339_);
  or _53855_ (_02342_, _02341_, _02338_);
  and _53856_ (_02343_, _01733_, _02045_);
  and _53857_ (_02344_, _01706_, _02070_);
  and _53858_ (_02345_, _01701_, _02048_);
  or _53859_ (_02346_, _02345_, _02344_);
  or _53860_ (_02347_, _02346_, _02343_);
  and _53861_ (_02348_, _01737_, _02056_);
  and _53862_ (_02349_, _01714_, _02053_);
  or _53863_ (_02350_, _02349_, _02348_);
  and _53864_ (_02351_, _01709_, _02061_);
  and _53865_ (_02352_, _01689_, _02022_);
  and _53866_ (_02353_, _01721_, _02068_);
  and _53867_ (_02354_, _01724_, _02030_);
  or _53868_ (_02355_, _02354_, _02353_);
  or _53869_ (_02356_, _02355_, _02352_);
  or _53870_ (_02357_, _02356_, _02351_);
  or _53871_ (_02358_, _02357_, _02350_);
  or _53872_ (_02359_, _02358_, _02347_);
  or _53873_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02359_, _02342_);
  and _53874_ (_02360_, _01661_, _02075_);
  and _53875_ (_02361_, _01680_, _02082_);
  and _53876_ (_02362_, _01689_, _02077_);
  or _53877_ (_02363_, _02362_, _02361_);
  and _53878_ (_02364_, _01676_, _02090_);
  and _53879_ (_02365_, _01717_, _02123_);
  or _53880_ (_02366_, _02365_, _02364_);
  or _53881_ (_02367_, _02366_, _02363_);
  or _53882_ (_02368_, _02367_, _02360_);
  and _53883_ (_02369_, _01670_, _02114_);
  and _53884_ (_02370_, _01665_, _02080_);
  or _53885_ (_02371_, _02370_, _02369_);
  or _53886_ (_02372_, _02371_, _02368_);
  and _53887_ (_02373_, _01733_, _02104_);
  and _53888_ (_02374_, _01701_, _02101_);
  and _53889_ (_02375_, _01737_, _02112_);
  or _53890_ (_02376_, _02375_, _02374_);
  or _53891_ (_02377_, _02376_, _02373_);
  and _53892_ (_02378_, _01709_, _02117_);
  and _53893_ (_02379_, _01706_, _02109_);
  or _53894_ (_02380_, _02379_, _02378_);
  and _53895_ (_02381_, _01714_, _02125_);
  and _53896_ (_02382_, _01685_, _02087_);
  and _53897_ (_02383_, _01721_, _02098_);
  and _53898_ (_02384_, _01724_, _02084_);
  or _53899_ (_02385_, _02384_, _02383_);
  or _53900_ (_02386_, _02385_, _02382_);
  or _53901_ (_02387_, _02386_, _02381_);
  or _53902_ (_02388_, _02387_, _02380_);
  or _53903_ (_02389_, _02388_, _02377_);
  or _53904_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _02389_, _02372_);
  and _53905_ (_02390_, _01665_, _02130_);
  and _53906_ (_02391_, _01676_, _02168_);
  and _53907_ (_02392_, _01689_, _02132_);
  or _53908_ (_02393_, _02392_, _02391_);
  and _53909_ (_02394_, _01685_, _02146_);
  and _53910_ (_02395_, _01717_, _02160_);
  or _53911_ (_02396_, _02395_, _02394_);
  or _53912_ (_02397_, _02396_, _02393_);
  or _53913_ (_02398_, _02397_, _02390_);
  and _53914_ (_02399_, _01670_, _02170_);
  and _53915_ (_02400_, _01661_, _02135_);
  or _53916_ (_02401_, _02400_, _02399_);
  or _53917_ (_02402_, _02401_, _02398_);
  and _53918_ (_02403_, _01733_, _02165_);
  and _53919_ (_02404_, _01701_, _02178_);
  and _53920_ (_02405_, _01714_, _02180_);
  or _53921_ (_02406_, _02405_, _02404_);
  or _53922_ (_02407_, _02406_, _02403_);
  and _53923_ (_02408_, _01709_, _02173_);
  and _53924_ (_02409_, _01706_, _02157_);
  or _53925_ (_02410_, _02409_, _02408_);
  and _53926_ (_02411_, _01737_, _02139_);
  and _53927_ (_02412_, _01680_, _02144_);
  and _53928_ (_02413_, _01721_, _02154_);
  and _53929_ (_02414_, _01724_, _02137_);
  or _53930_ (_02415_, _02414_, _02413_);
  or _53931_ (_02416_, _02415_, _02412_);
  or _53932_ (_02417_, _02416_, _02411_);
  or _53933_ (_02418_, _02417_, _02410_);
  or _53934_ (_02419_, _02418_, _02407_);
  or _53935_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _02419_, _02402_);
  and _53936_ (_02420_, _01670_, _02226_);
  and _53937_ (_02421_, _01680_, _02196_);
  and _53938_ (_02422_, _01685_, _02224_);
  or _53939_ (_02423_, _02422_, _02421_);
  and _53940_ (_02424_, _01676_, _02200_);
  and _53941_ (_02425_, _01689_, _02187_);
  or _53942_ (_02426_, _02425_, _02424_);
  or _53943_ (_02427_, _02426_, _02423_);
  or _53944_ (_02428_, _02427_, _02420_);
  and _53945_ (_02429_, _01661_, _02185_);
  and _53946_ (_02430_, _01665_, _02190_);
  or _53947_ (_02431_, _02430_, _02429_);
  or _53948_ (_02432_, _02431_, _02428_);
  and _53949_ (_02433_, _01706_, _02235_);
  and _53950_ (_02434_, _01733_, _02233_);
  and _53951_ (_02435_, _01701_, _02213_);
  or _53952_ (_02436_, _02435_, _02434_);
  or _53953_ (_02437_, _02436_, _02433_);
  and _53954_ (_02438_, _01714_, _02217_);
  and _53955_ (_02439_, _01717_, _02210_);
  and _53956_ (_02440_, _01721_, _02221_);
  and _53957_ (_02441_, _01724_, _02193_);
  or _53958_ (_02442_, _02441_, _02440_);
  or _53959_ (_02443_, _02442_, _02439_);
  or _53960_ (_02444_, _02443_, _02438_);
  and _53961_ (_02445_, _01709_, _02228_);
  and _53962_ (_02446_, _01737_, _02202_);
  or _53963_ (_02447_, _02446_, _02445_);
  or _53964_ (_02448_, _02447_, _02444_);
  or _53965_ (_02449_, _02448_, _02437_);
  or _53966_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02449_, _02432_);
  and _53967_ (_02450_, _01661_, _01890_);
  and _53968_ (_02451_, _01670_, _01902_);
  or _53969_ (_02452_, _02451_, _02450_);
  and _53970_ (_02453_, _01665_, _01869_);
  and _53971_ (_02454_, _01685_, _01877_);
  and _53972_ (_02455_, _01676_, _01888_);
  or _53973_ (_02456_, _02455_, _02454_);
  and _53974_ (_02457_, _01717_, _01885_);
  and _53975_ (_02458_, _01680_, _01864_);
  or _53976_ (_02459_, _02458_, _02457_);
  or _53977_ (_02460_, _02459_, _02456_);
  or _53978_ (_02461_, _02460_, _02453_);
  or _53979_ (_02462_, _02461_, _02452_);
  and _53980_ (_02463_, _01706_, _01893_);
  and _53981_ (_02464_, _01701_, _01900_);
  and _53982_ (_02466_, _01733_, _01875_);
  or _53983_ (_02467_, _02466_, _02464_);
  or _53984_ (_02468_, _02467_, _02463_);
  and _53985_ (_02469_, _01737_, _01853_);
  and _53986_ (_02470_, _01689_, _01871_);
  and _53987_ (_02471_, _01724_, _01862_);
  and _53988_ (_02472_, _01721_, _01879_);
  or _53989_ (_02473_, _02472_, _02471_);
  or _53990_ (_02474_, _02473_, _02470_);
  or _53991_ (_02475_, _02474_, _02469_);
  and _53992_ (_02476_, _01714_, _01856_);
  and _53993_ (_02477_, _01709_, _01859_);
  or _53994_ (_02478_, _02477_, _02476_);
  or _53995_ (_02479_, _02478_, _02475_);
  or _53996_ (_02480_, _02479_, _02468_);
  or _53997_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _02480_, _02462_);
  and _53998_ (_02481_, _01661_, _01946_);
  and _53999_ (_02482_, _01676_, _01917_);
  and _54000_ (_02483_, _01685_, _01933_);
  or _54001_ (_02484_, _02483_, _02482_);
  and _54002_ (_02485_, _01717_, _01930_);
  and _54003_ (_02486_, _01689_, _01926_);
  or _54004_ (_02487_, _02486_, _02485_);
  or _54005_ (_02488_, _02487_, _02484_);
  or _54006_ (_02489_, _02488_, _02481_);
  and _54007_ (_02490_, _01670_, _01958_);
  and _54008_ (_02491_, _01665_, _01924_);
  or _54009_ (_02492_, _02491_, _02490_);
  or _54010_ (_02493_, _02492_, _02489_);
  and _54011_ (_02494_, _01706_, _01949_);
  and _54012_ (_02495_, _01709_, _01914_);
  and _54013_ (_02496_, _01737_, _01909_);
  or _54014_ (_02497_, _02496_, _02495_);
  or _54015_ (_02498_, _02497_, _02494_);
  and _54016_ (_02499_, _01701_, _01956_);
  and _54017_ (_02500_, _01714_, _01944_);
  or _54018_ (_02501_, _02500_, _02499_);
  and _54019_ (_02502_, _01733_, _01941_);
  and _54020_ (_02503_, _01680_, _01919_);
  and _54021_ (_02504_, _01721_, _01937_);
  and _54022_ (_02505_, _01724_, _01912_);
  or _54023_ (_02506_, _02505_, _02504_);
  or _54024_ (_02507_, _02506_, _02503_);
  or _54025_ (_02508_, _02507_, _02502_);
  or _54026_ (_02509_, _02508_, _02501_);
  or _54027_ (_02510_, _02509_, _02498_);
  or _54028_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _02510_, _02493_);
  and _54029_ (_02511_, _01661_, _02002_);
  and _54030_ (_02512_, _01670_, _01989_);
  or _54031_ (_02513_, _02512_, _02511_);
  and _54032_ (_02514_, _01665_, _01965_);
  and _54033_ (_02515_, _01676_, _01977_);
  and _54034_ (_02516_, _01685_, _01992_);
  or _54035_ (_02517_, _02516_, _02515_);
  and _54036_ (_02518_, _01717_, _01986_);
  and _54037_ (_02519_, _01689_, _01970_);
  or _54038_ (_02520_, _02519_, _02518_);
  or _54039_ (_02521_, _02520_, _02517_);
  or _54040_ (_02522_, _02521_, _02514_);
  or _54041_ (_02523_, _02522_, _02513_);
  and _54042_ (_02524_, _01737_, _01967_);
  and _54043_ (_02525_, _01709_, _01972_);
  and _54044_ (_02526_, _01706_, _02005_);
  or _54045_ (_02527_, _02526_, _02525_);
  or _54046_ (_02528_, _02527_, _02524_);
  and _54047_ (_02529_, _01701_, _02014_);
  and _54048_ (_02530_, _01714_, _01979_);
  or _54049_ (_02531_, _02530_, _02529_);
  and _54050_ (_02532_, _01733_, _02012_);
  and _54051_ (_02533_, _01680_, _02000_);
  and _54052_ (_02534_, _01724_, _01974_);
  and _54053_ (_02535_, _01721_, _01997_);
  or _54054_ (_02536_, _02535_, _02534_);
  or _54055_ (_02537_, _02536_, _02533_);
  or _54056_ (_02538_, _02537_, _02532_);
  or _54057_ (_02539_, _02538_, _02531_);
  or _54058_ (_02540_, _02539_, _02528_);
  or _54059_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _02540_, _02523_);
  and _54060_ (_02541_, _01661_, _02058_);
  and _54061_ (_02542_, _01676_, _02025_);
  and _54062_ (_02543_, _01685_, _02042_);
  or _54063_ (_02544_, _02543_, _02542_);
  and _54064_ (_02545_, _01689_, _02037_);
  and _54065_ (_02546_, _01717_, _02048_);
  or _54066_ (_02547_, _02546_, _02545_);
  or _54067_ (_02548_, _02547_, _02544_);
  or _54068_ (_02549_, _02548_, _02541_);
  and _54069_ (_02550_, _01670_, _02068_);
  and _54070_ (_02551_, _01665_, _02020_);
  or _54071_ (_02552_, _02551_, _02550_);
  or _54072_ (_02553_, _02552_, _02549_);
  and _54073_ (_02554_, _01706_, _02061_);
  and _54074_ (_02555_, _01709_, _02030_);
  and _54075_ (_02556_, _01737_, _02022_);
  or _54076_ (_02557_, _02556_, _02555_);
  or _54077_ (_02558_, _02557_, _02554_);
  and _54078_ (_02559_, _01701_, _02053_);
  and _54079_ (_02560_, _01714_, _02056_);
  or _54080_ (_02561_, _02560_, _02559_);
  and _54081_ (_02562_, _01733_, _02070_);
  and _54082_ (_02563_, _01680_, _02027_);
  and _54083_ (_02564_, _01721_, _02045_);
  and _54084_ (_02565_, _01724_, _02032_);
  or _54085_ (_02566_, _02565_, _02564_);
  or _54086_ (_02567_, _02566_, _02563_);
  or _54087_ (_02568_, _02567_, _02562_);
  or _54088_ (_02569_, _02568_, _02561_);
  or _54089_ (_02570_, _02569_, _02558_);
  or _54090_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _02570_, _02553_);
  and _54091_ (_02571_, _01661_, _02114_);
  and _54092_ (_02572_, _01680_, _02090_);
  and _54093_ (_02573_, _01676_, _02087_);
  or _54094_ (_02574_, _02573_, _02572_);
  and _54095_ (_02575_, _01717_, _02101_);
  and _54096_ (_02576_, _01689_, _02080_);
  or _54097_ (_02577_, _02576_, _02575_);
  or _54098_ (_02578_, _02577_, _02574_);
  or _54099_ (_02579_, _02578_, _02571_);
  and _54100_ (_02580_, _01665_, _02075_);
  and _54101_ (_02581_, _01670_, _02098_);
  or _54102_ (_02582_, _02581_, _02580_);
  or _54103_ (_02583_, _02582_, _02579_);
  and _54104_ (_02584_, _01737_, _02077_);
  and _54105_ (_02585_, _01701_, _02125_);
  and _54106_ (_02586_, _01706_, _02117_);
  or _54107_ (_02587_, _02586_, _02585_);
  or _54108_ (_02588_, _02587_, _02584_);
  and _54109_ (_02589_, _01709_, _02084_);
  and _54110_ (_02590_, _01685_, _02123_);
  and _54111_ (_02591_, _01724_, _02082_);
  and _54112_ (_02592_, _01721_, _02104_);
  or _54113_ (_02593_, _02592_, _02591_);
  or _54114_ (_02594_, _02593_, _02590_);
  or _54115_ (_02595_, _02594_, _02589_);
  and _54116_ (_02596_, _01714_, _02112_);
  and _54117_ (_02597_, _01733_, _02109_);
  or _54118_ (_02598_, _02597_, _02596_);
  or _54119_ (_02599_, _02598_, _02595_);
  or _54120_ (_02600_, _02599_, _02588_);
  or _54121_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _02600_, _02583_);
  and _54122_ (_02601_, _01661_, _02170_);
  and _54123_ (_02602_, _01670_, _02154_);
  or _54124_ (_02603_, _02602_, _02601_);
  and _54125_ (_02604_, _01665_, _02135_);
  and _54126_ (_02605_, _01685_, _02160_);
  and _54127_ (_02606_, _01676_, _02146_);
  or _54128_ (_02607_, _02606_, _02605_);
  and _54129_ (_02608_, _01717_, _02178_);
  and _54130_ (_02609_, _01680_, _02168_);
  or _54131_ (_02610_, _02609_, _02608_);
  or _54132_ (_02611_, _02610_, _02607_);
  or _54133_ (_02612_, _02611_, _02604_);
  or _54134_ (_02613_, _02612_, _02603_);
  and _54135_ (_02614_, _01709_, _02137_);
  and _54136_ (_02615_, _01714_, _02139_);
  and _54137_ (_02616_, _01706_, _02173_);
  or _54138_ (_02617_, _02616_, _02615_);
  or _54139_ (_02618_, _02617_, _02614_);
  and _54140_ (_02619_, _01733_, _02157_);
  and _54141_ (_02620_, _01689_, _02130_);
  and _54142_ (_02621_, _01724_, _02144_);
  and _54143_ (_02622_, _01721_, _02165_);
  or _54144_ (_02623_, _02622_, _02621_);
  or _54145_ (_02624_, _02623_, _02620_);
  or _54146_ (_02625_, _02624_, _02619_);
  and _54147_ (_02626_, _01701_, _02180_);
  and _54148_ (_02627_, _01737_, _02132_);
  or _54149_ (_02628_, _02627_, _02626_);
  or _54150_ (_02629_, _02628_, _02625_);
  or _54151_ (_02630_, _02629_, _02618_);
  or _54152_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _02630_, _02613_);
  and _54153_ (_02631_, _01670_, _02221_);
  and _54154_ (_02632_, _01676_, _02224_);
  and _54155_ (_02633_, _01717_, _02213_);
  or _54156_ (_02634_, _02633_, _02632_);
  and _54157_ (_02635_, _01680_, _02200_);
  and _54158_ (_02636_, _01689_, _02190_);
  or _54159_ (_02637_, _02636_, _02635_);
  or _54160_ (_02638_, _02637_, _02634_);
  or _54161_ (_02639_, _02638_, _02631_);
  and _54162_ (_02640_, _01661_, _02226_);
  and _54163_ (_02641_, _01665_, _02185_);
  or _54164_ (_02642_, _02641_, _02640_);
  or _54165_ (_02643_, _02642_, _02639_);
  and _54166_ (_02644_, _01709_, _02193_);
  and _54167_ (_02645_, _01733_, _02235_);
  and _54168_ (_02646_, _01714_, _02202_);
  or _54169_ (_02647_, _02646_, _02645_);
  or _54170_ (_02648_, _02647_, _02644_);
  and _54171_ (_02649_, _01737_, _02187_);
  and _54172_ (_02650_, _01685_, _02210_);
  and _54173_ (_02651_, _01721_, _02233_);
  and _54174_ (_02652_, _01724_, _02196_);
  or _54175_ (_02653_, _02652_, _02651_);
  or _54176_ (_02654_, _02653_, _02650_);
  or _54177_ (_02655_, _02654_, _02649_);
  and _54178_ (_02656_, _01706_, _02228_);
  and _54179_ (_02657_, _01701_, _02217_);
  or _54180_ (_02658_, _02657_, _02656_);
  or _54181_ (_02659_, _02658_, _02655_);
  or _54182_ (_02661_, _02659_, _02648_);
  or _54183_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _02661_, _02643_);
  and _54184_ (_02662_, _01661_, _01902_);
  and _54185_ (_02663_, _01670_, _01879_);
  or _54186_ (_02664_, _02663_, _02662_);
  and _54187_ (_02665_, _01665_, _01890_);
  and _54188_ (_02666_, _01685_, _01885_);
  and _54189_ (_02667_, _01717_, _01900_);
  or _54190_ (_02668_, _02667_, _02666_);
  and _54191_ (_02669_, _01680_, _01888_);
  and _54192_ (_02670_, _01676_, _01877_);
  or _54193_ (_02671_, _02670_, _02669_);
  or _54194_ (_02672_, _02671_, _02668_);
  or _54195_ (_02673_, _02672_, _02665_);
  or _54196_ (_02674_, _02673_, _02664_);
  and _54197_ (_02675_, _01706_, _01859_);
  and _54198_ (_02676_, _01733_, _01893_);
  and _54199_ (_02677_, _01701_, _01856_);
  or _54200_ (_02678_, _02677_, _02676_);
  or _54201_ (_02679_, _02678_, _02675_);
  and _54202_ (_02680_, _01714_, _01853_);
  and _54203_ (_02681_, _01689_, _01869_);
  and _54204_ (_02682_, _01724_, _01864_);
  and _54205_ (_02683_, _01721_, _01875_);
  or _54206_ (_02684_, _02683_, _02682_);
  or _54207_ (_02685_, _02684_, _02681_);
  or _54208_ (_02686_, _02685_, _02680_);
  and _54209_ (_02687_, _01709_, _01862_);
  and _54210_ (_02688_, _01737_, _01871_);
  or _54211_ (_02689_, _02688_, _02687_);
  or _54212_ (_02690_, _02689_, _02686_);
  or _54213_ (_02691_, _02690_, _02679_);
  or _54214_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02691_, _02674_);
  and _54215_ (_02692_, _01670_, _01937_);
  and _54216_ (_02693_, _01661_, _01958_);
  or _54217_ (_02694_, _02693_, _02692_);
  and _54218_ (_02695_, _01665_, _01946_);
  and _54219_ (_02696_, _01717_, _01956_);
  and _54220_ (_02697_, _01689_, _01924_);
  or _54221_ (_02698_, _02697_, _02696_);
  and _54222_ (_02699_, _01680_, _01917_);
  and _54223_ (_02700_, _01676_, _01933_);
  or _54224_ (_02701_, _02700_, _02699_);
  or _54225_ (_02702_, _02701_, _02698_);
  or _54226_ (_02703_, _02702_, _02695_);
  or _54227_ (_02704_, _02703_, _02694_);
  and _54228_ (_02705_, _01709_, _01912_);
  and _54229_ (_02706_, _01706_, _01914_);
  and _54230_ (_02707_, _01737_, _01926_);
  or _54231_ (_02708_, _02707_, _02706_);
  or _54232_ (_02709_, _02708_, _02705_);
  and _54233_ (_02710_, _01714_, _01909_);
  and _54234_ (_02711_, _01685_, _01930_);
  and _54235_ (_02712_, _01721_, _01941_);
  and _54236_ (_02713_, _01724_, _01919_);
  or _54237_ (_02714_, _02713_, _02712_);
  or _54238_ (_02715_, _02714_, _02711_);
  or _54239_ (_02716_, _02715_, _02710_);
  and _54240_ (_02717_, _01733_, _01949_);
  and _54241_ (_02718_, _01701_, _01944_);
  or _54242_ (_02719_, _02718_, _02717_);
  or _54243_ (_02720_, _02719_, _02716_);
  or _54244_ (_02721_, _02720_, _02709_);
  or _54245_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02721_, _02704_);
  and _54246_ (_02722_, _01661_, _01989_);
  and _54247_ (_02723_, _01680_, _01977_);
  and _54248_ (_02724_, _01685_, _01986_);
  or _54249_ (_02725_, _02724_, _02723_);
  and _54250_ (_02726_, _01676_, _01992_);
  and _54251_ (_02727_, _01717_, _02014_);
  or _54252_ (_02728_, _02727_, _02726_);
  or _54253_ (_02729_, _02728_, _02725_);
  or _54254_ (_02730_, _02729_, _02722_);
  and _54255_ (_02731_, _01665_, _02002_);
  and _54256_ (_02732_, _01670_, _01997_);
  or _54257_ (_02733_, _02732_, _02731_);
  or _54258_ (_02734_, _02733_, _02730_);
  and _54259_ (_02735_, _01709_, _01974_);
  and _54260_ (_02736_, _01701_, _01979_);
  and _54261_ (_02737_, _01714_, _01967_);
  or _54262_ (_02738_, _02737_, _02736_);
  or _54263_ (_02739_, _02738_, _02735_);
  and _54264_ (_02740_, _01733_, _02005_);
  and _54265_ (_02741_, _01689_, _01965_);
  and _54266_ (_02742_, _01721_, _02012_);
  and _54267_ (_02743_, _01724_, _02000_);
  or _54268_ (_02744_, _02743_, _02742_);
  or _54269_ (_02745_, _02744_, _02741_);
  or _54270_ (_02746_, _02745_, _02740_);
  and _54271_ (_02747_, _01706_, _01972_);
  and _54272_ (_02748_, _01737_, _01970_);
  or _54273_ (_02749_, _02748_, _02747_);
  or _54274_ (_02750_, _02749_, _02746_);
  or _54275_ (_02751_, _02750_, _02739_);
  or _54276_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02751_, _02734_);
  and _54277_ (_02752_, _01661_, _02068_);
  and _54278_ (_02753_, _01717_, _02053_);
  and _54279_ (_02754_, _01680_, _02025_);
  or _54280_ (_02755_, _02754_, _02753_);
  and _54281_ (_02756_, _01676_, _02042_);
  and _54282_ (_02757_, _01689_, _02020_);
  or _54283_ (_02758_, _02757_, _02756_);
  or _54284_ (_02759_, _02758_, _02755_);
  or _54285_ (_02760_, _02759_, _02752_);
  and _54286_ (_02761_, _01665_, _02058_);
  and _54287_ (_02762_, _01670_, _02045_);
  or _54288_ (_02763_, _02762_, _02761_);
  or _54289_ (_02764_, _02763_, _02760_);
  and _54290_ (_02765_, _01709_, _02032_);
  and _54291_ (_02766_, _01737_, _02037_);
  and _54292_ (_02767_, _01706_, _02030_);
  or _54293_ (_02768_, _02767_, _02766_);
  or _54294_ (_02769_, _02768_, _02765_);
  and _54295_ (_02770_, _01701_, _02056_);
  and _54296_ (_02771_, _01685_, _02048_);
  and _54297_ (_02772_, _01724_, _02027_);
  and _54298_ (_02773_, _01721_, _02070_);
  or _54299_ (_02774_, _02773_, _02772_);
  or _54300_ (_02775_, _02774_, _02771_);
  or _54301_ (_02776_, _02775_, _02770_);
  and _54302_ (_02777_, _01714_, _02022_);
  and _54303_ (_02778_, _01733_, _02061_);
  or _54304_ (_02779_, _02778_, _02777_);
  or _54305_ (_02780_, _02779_, _02776_);
  or _54306_ (_02781_, _02780_, _02769_);
  or _54307_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02781_, _02764_);
  and _54308_ (_02782_, _01661_, _02098_);
  and _54309_ (_02783_, _01689_, _02075_);
  and _54310_ (_02784_, _01676_, _02123_);
  or _54311_ (_02785_, _02784_, _02783_);
  and _54312_ (_02786_, _01680_, _02087_);
  and _54313_ (_02787_, _01685_, _02101_);
  or _54314_ (_02788_, _02787_, _02786_);
  or _54315_ (_02789_, _02788_, _02785_);
  or _54316_ (_02790_, _02789_, _02782_);
  and _54317_ (_02791_, _01665_, _02114_);
  and _54318_ (_02792_, _01670_, _02104_);
  or _54319_ (_02793_, _02792_, _02791_);
  or _54320_ (_02794_, _02793_, _02790_);
  and _54321_ (_02795_, _01714_, _02077_);
  and _54322_ (_02796_, _01733_, _02117_);
  and _54323_ (_02797_, _01709_, _02082_);
  or _54324_ (_02798_, _02797_, _02796_);
  or _54325_ (_02799_, _02798_, _02795_);
  and _54326_ (_02800_, _01737_, _02080_);
  and _54327_ (_02801_, _01717_, _02125_);
  and _54328_ (_02802_, _01721_, _02109_);
  and _54329_ (_02803_, _01724_, _02090_);
  or _54330_ (_02804_, _02803_, _02802_);
  or _54331_ (_02805_, _02804_, _02801_);
  or _54332_ (_02806_, _02805_, _02800_);
  and _54333_ (_02807_, _01706_, _02084_);
  and _54334_ (_02808_, _01701_, _02112_);
  or _54335_ (_02809_, _02808_, _02807_);
  or _54336_ (_02810_, _02809_, _02806_);
  or _54337_ (_02811_, _02810_, _02799_);
  or _54338_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02811_, _02794_);
  and _54339_ (_02812_, _01661_, _02154_);
  and _54340_ (_02813_, _01689_, _02135_);
  and _54341_ (_02814_, _01676_, _02160_);
  or _54342_ (_02815_, _02814_, _02813_);
  and _54343_ (_02816_, _01685_, _02178_);
  and _54344_ (_02817_, _01717_, _02180_);
  or _54345_ (_02818_, _02817_, _02816_);
  or _54346_ (_02819_, _02818_, _02815_);
  or _54347_ (_02820_, _02819_, _02812_);
  and _54348_ (_02821_, _01665_, _02170_);
  and _54349_ (_02822_, _01670_, _02165_);
  or _54350_ (_02823_, _02822_, _02821_);
  or _54351_ (_02824_, _02823_, _02820_);
  and _54352_ (_02825_, _01714_, _02132_);
  and _54353_ (_02826_, _01733_, _02173_);
  and _54354_ (_02827_, _01706_, _02137_);
  or _54355_ (_02828_, _02827_, _02826_);
  or _54356_ (_02829_, _02828_, _02825_);
  and _54357_ (_02830_, _01701_, _02139_);
  and _54358_ (_02831_, _01680_, _02146_);
  and _54359_ (_02832_, _01721_, _02157_);
  and _54360_ (_02833_, _01724_, _02168_);
  or _54361_ (_02834_, _02833_, _02832_);
  or _54362_ (_02835_, _02834_, _02831_);
  or _54363_ (_02836_, _02835_, _02830_);
  and _54364_ (_02837_, _01709_, _02144_);
  and _54365_ (_02838_, _01737_, _02130_);
  or _54366_ (_02839_, _02838_, _02837_);
  or _54367_ (_02840_, _02839_, _02836_);
  or _54368_ (_02841_, _02840_, _02829_);
  or _54369_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02841_, _02824_);
  and _54370_ (_02842_, _01661_, _02221_);
  and _54371_ (_02843_, _01676_, _02210_);
  and _54372_ (_02844_, _01685_, _02213_);
  or _54373_ (_02845_, _02844_, _02843_);
  and _54374_ (_02846_, _01680_, _02224_);
  and _54375_ (_02847_, _01689_, _02185_);
  or _54376_ (_02848_, _02847_, _02846_);
  or _54377_ (_02849_, _02848_, _02845_);
  or _54378_ (_02850_, _02849_, _02842_);
  and _54379_ (_02851_, _01665_, _02226_);
  and _54380_ (_02852_, _01670_, _02233_);
  or _54381_ (_02853_, _02852_, _02851_);
  or _54382_ (_02855_, _02853_, _02850_);
  and _54383_ (_02856_, _01733_, _02228_);
  and _54384_ (_02857_, _01709_, _02196_);
  and _54385_ (_02858_, _01737_, _02190_);
  or _54386_ (_02859_, _02858_, _02857_);
  or _54387_ (_02860_, _02859_, _02856_);
  and _54388_ (_02861_, _01706_, _02193_);
  and _54389_ (_02862_, _01717_, _02217_);
  and _54390_ (_02863_, _01721_, _02235_);
  and _54391_ (_02864_, _01724_, _02200_);
  or _54392_ (_02865_, _02864_, _02863_);
  or _54393_ (_02866_, _02865_, _02862_);
  or _54394_ (_02867_, _02866_, _02861_);
  and _54395_ (_02868_, _01701_, _02202_);
  and _54396_ (_02869_, _01714_, _02187_);
  or _54397_ (_02870_, _02869_, _02868_);
  or _54398_ (_02871_, _02870_, _02867_);
  or _54399_ (_02872_, _02871_, _02860_);
  or _54400_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02872_, _02855_);
  nand _54401_ (_02873_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not _54402_ (_02874_, \oc8051_golden_model_1.PC [3]);
  or _54403_ (_02875_, \oc8051_golden_model_1.PC [2], _02874_);
  or _54404_ (_02876_, _02875_, _02873_);
  or _54405_ (_02877_, _02876_, _42137_);
  not _54406_ (_02878_, \oc8051_golden_model_1.PC [1]);
  or _54407_ (_02879_, _02878_, \oc8051_golden_model_1.PC [0]);
  or _54408_ (_02880_, _02879_, _02875_);
  or _54409_ (_02881_, _02880_, _42096_);
  and _54410_ (_02882_, _02881_, _02877_);
  not _54411_ (_02883_, \oc8051_golden_model_1.PC [2]);
  or _54412_ (_02884_, _02883_, \oc8051_golden_model_1.PC [3]);
  or _54413_ (_02885_, _02884_, _02873_);
  or _54414_ (_02886_, _02885_, _41973_);
  or _54415_ (_02887_, _02884_, _02879_);
  or _54416_ (_02888_, _02887_, _41932_);
  and _54417_ (_02889_, _02888_, _02886_);
  and _54418_ (_02890_, _02889_, _02882_);
  nand _54419_ (_02891_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _54420_ (_02892_, _02891_, _02873_);
  or _54421_ (_02893_, _02892_, _42301_);
  or _54422_ (_02894_, _02891_, _02879_);
  or _54423_ (_02895_, _02894_, _42260_);
  and _54424_ (_02896_, _02895_, _02893_);
  or _54425_ (_02897_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _54426_ (_02898_, _02897_, _02873_);
  or _54427_ (_02899_, _02898_, _41809_);
  or _54428_ (_02900_, _02897_, _02879_);
  or _54429_ (_02901_, _02900_, _41758_);
  and _54430_ (_02902_, _02901_, _02899_);
  and _54431_ (_02903_, _02902_, _02896_);
  and _54432_ (_02904_, _02903_, _02890_);
  not _54433_ (_02905_, \oc8051_golden_model_1.PC [0]);
  or _54434_ (_02906_, \oc8051_golden_model_1.PC [1], _02905_);
  or _54435_ (_02907_, _02906_, _02891_);
  or _54436_ (_02908_, _02907_, _42219_);
  or _54437_ (_02909_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or _54438_ (_02910_, _02909_, _02891_);
  or _54439_ (_02911_, _02910_, _42178_);
  and _54440_ (_02912_, _02911_, _02908_);
  or _54441_ (_02913_, _02897_, _02909_);
  or _54442_ (_02914_, _02913_, _41671_);
  or _54443_ (_02915_, _02897_, _02906_);
  or _54444_ (_02916_, _02915_, _41712_);
  and _54445_ (_02917_, _02916_, _02914_);
  and _54446_ (_02918_, _02917_, _02912_);
  or _54447_ (_02919_, _02906_, _02875_);
  or _54448_ (_02920_, _02919_, _42055_);
  or _54449_ (_02921_, _02909_, _02875_);
  or _54450_ (_02922_, _02921_, _42014_);
  and _54451_ (_02923_, _02922_, _02920_);
  or _54452_ (_02924_, _02906_, _02884_);
  or _54453_ (_02925_, _02924_, _41891_);
  or _54454_ (_02926_, _02909_, _02884_);
  or _54455_ (_02927_, _02926_, _41850_);
  and _54456_ (_02928_, _02927_, _02925_);
  and _54457_ (_02929_, _02928_, _02923_);
  and _54458_ (_02930_, _02929_, _02918_);
  nand _54459_ (_02931_, _02930_, _02904_);
  or _54460_ (_02932_, _02876_, _42142_);
  or _54461_ (_02933_, _02880_, _42101_);
  and _54462_ (_02934_, _02933_, _02932_);
  or _54463_ (_02935_, _02885_, _41978_);
  or _54464_ (_02936_, _02887_, _41937_);
  and _54465_ (_02937_, _02936_, _02935_);
  and _54466_ (_02938_, _02937_, _02934_);
  or _54467_ (_02939_, _02892_, _42306_);
  or _54468_ (_02940_, _02894_, _42265_);
  and _54469_ (_02941_, _02940_, _02939_);
  or _54470_ (_02942_, _02898_, _41814_);
  or _54471_ (_02943_, _02900_, _41765_);
  and _54472_ (_02944_, _02943_, _02942_);
  and _54473_ (_02945_, _02944_, _02941_);
  and _54474_ (_02946_, _02945_, _02938_);
  or _54475_ (_02947_, _02907_, _42224_);
  or _54476_ (_02948_, _02910_, _42183_);
  and _54477_ (_02949_, _02948_, _02947_);
  or _54478_ (_02950_, _02913_, _41676_);
  or _54479_ (_02951_, _02915_, _41717_);
  and _54480_ (_02952_, _02951_, _02950_);
  and _54481_ (_02953_, _02952_, _02949_);
  or _54482_ (_02954_, _02919_, _42060_);
  or _54483_ (_02955_, _02921_, _42019_);
  and _54484_ (_02956_, _02955_, _02954_);
  or _54485_ (_02957_, _02924_, _41896_);
  or _54486_ (_02958_, _02926_, _41855_);
  and _54487_ (_02959_, _02958_, _02957_);
  and _54488_ (_02960_, _02959_, _02956_);
  and _54489_ (_02961_, _02960_, _02953_);
  nand _54490_ (_02962_, _02961_, _02946_);
  or _54491_ (_02963_, _02962_, _02931_);
  or _54492_ (_02964_, _02876_, _42127_);
  or _54493_ (_02965_, _02880_, _42086_);
  and _54494_ (_02966_, _02965_, _02964_);
  or _54495_ (_02967_, _02885_, _41963_);
  or _54496_ (_02968_, _02887_, _41922_);
  and _54497_ (_02969_, _02968_, _02967_);
  and _54498_ (_02970_, _02969_, _02966_);
  or _54499_ (_02971_, _02892_, _42291_);
  or _54500_ (_02972_, _02894_, _42250_);
  and _54501_ (_02973_, _02972_, _02971_);
  or _54502_ (_02974_, _02898_, _41791_);
  or _54503_ (_02975_, _02900_, _41743_);
  and _54504_ (_02976_, _02975_, _02974_);
  and _54505_ (_02977_, _02976_, _02973_);
  and _54506_ (_02978_, _02977_, _02970_);
  or _54507_ (_02979_, _02907_, _42209_);
  or _54508_ (_02980_, _02910_, _42168_);
  and _54509_ (_02981_, _02980_, _02979_);
  or _54510_ (_02982_, _02913_, _41661_);
  or _54511_ (_02983_, _02915_, _41702_);
  and _54512_ (_02984_, _02983_, _02982_);
  and _54513_ (_02985_, _02984_, _02981_);
  or _54514_ (_02986_, _02919_, _42045_);
  or _54515_ (_02987_, _02921_, _42004_);
  and _54516_ (_02988_, _02987_, _02986_);
  or _54517_ (_02989_, _02924_, _41881_);
  or _54518_ (_02990_, _02926_, _41840_);
  and _54519_ (_02991_, _02990_, _02989_);
  and _54520_ (_02992_, _02991_, _02988_);
  and _54521_ (_02993_, _02992_, _02985_);
  and _54522_ (_02994_, _02993_, _02978_);
  or _54523_ (_02995_, _02876_, _42132_);
  or _54524_ (_02996_, _02880_, _42091_);
  and _54525_ (_02997_, _02996_, _02995_);
  or _54526_ (_02998_, _02885_, _41968_);
  or _54527_ (_02999_, _02887_, _41927_);
  and _54528_ (_03000_, _02999_, _02998_);
  and _54529_ (_03001_, _03000_, _02997_);
  or _54530_ (_03002_, _02892_, _42296_);
  or _54531_ (_03003_, _02894_, _42255_);
  and _54532_ (_03004_, _03003_, _03002_);
  or _54533_ (_03005_, _02898_, _41801_);
  or _54534_ (_03006_, _02900_, _41749_);
  and _54535_ (_03007_, _03006_, _03005_);
  and _54536_ (_03008_, _03007_, _03004_);
  and _54537_ (_03009_, _03008_, _03001_);
  or _54538_ (_03010_, _02907_, _42214_);
  or _54539_ (_03011_, _02910_, _42173_);
  and _54540_ (_03012_, _03011_, _03010_);
  or _54541_ (_03013_, _02913_, _41666_);
  or _54542_ (_03015_, _02915_, _41707_);
  and _54543_ (_03016_, _03015_, _03013_);
  and _54544_ (_03017_, _03016_, _03012_);
  or _54545_ (_03018_, _02919_, _42050_);
  or _54546_ (_03019_, _02921_, _42009_);
  and _54547_ (_03020_, _03019_, _03018_);
  or _54548_ (_03021_, _02924_, _41886_);
  or _54549_ (_03022_, _02926_, _41845_);
  and _54550_ (_03023_, _03022_, _03021_);
  and _54551_ (_03024_, _03023_, _03020_);
  and _54552_ (_03026_, _03024_, _03017_);
  nand _54553_ (_03027_, _03026_, _03009_);
  or _54554_ (_03028_, _03027_, _02994_);
  or _54555_ (_03029_, _03028_, _02963_);
  not _54556_ (_03030_, _03029_);
  or _54557_ (_03031_, _02876_, _42147_);
  or _54558_ (_03032_, _02880_, _42106_);
  and _54559_ (_03033_, _03032_, _03031_);
  or _54560_ (_03034_, _02885_, _41983_);
  or _54561_ (_03035_, _02887_, _41942_);
  and _54562_ (_03036_, _03035_, _03034_);
  and _54563_ (_03037_, _03036_, _03033_);
  or _54564_ (_03038_, _02892_, _42311_);
  or _54565_ (_03039_, _02894_, _42270_);
  and _54566_ (_03040_, _03039_, _03038_);
  or _54567_ (_03041_, _02898_, _41819_);
  or _54568_ (_03042_, _02900_, _41770_);
  and _54569_ (_03043_, _03042_, _03041_);
  and _54570_ (_03044_, _03043_, _03040_);
  and _54571_ (_03045_, _03044_, _03037_);
  or _54572_ (_03047_, _02907_, _42229_);
  or _54573_ (_03048_, _02910_, _42188_);
  and _54574_ (_03049_, _03048_, _03047_);
  or _54575_ (_03050_, _02913_, _41681_);
  or _54576_ (_03051_, _02915_, _41722_);
  and _54577_ (_03052_, _03051_, _03050_);
  and _54578_ (_03053_, _03052_, _03049_);
  or _54579_ (_03054_, _02919_, _42065_);
  or _54580_ (_03055_, _02921_, _42024_);
  and _54581_ (_03056_, _03055_, _03054_);
  or _54582_ (_03058_, _02924_, _41901_);
  or _54583_ (_03059_, _02926_, _41860_);
  and _54584_ (_03060_, _03059_, _03058_);
  and _54585_ (_03061_, _03060_, _03056_);
  and _54586_ (_03062_, _03061_, _03053_);
  nand _54587_ (_03063_, _03062_, _03045_);
  or _54588_ (_03064_, _02876_, _42152_);
  or _54589_ (_03065_, _02880_, _42111_);
  and _54590_ (_03066_, _03065_, _03064_);
  or _54591_ (_03067_, _02885_, _41988_);
  or _54592_ (_03069_, _02887_, _41947_);
  and _54593_ (_03070_, _03069_, _03067_);
  and _54594_ (_03071_, _03070_, _03066_);
  or _54595_ (_03072_, _02892_, _42316_);
  or _54596_ (_03073_, _02894_, _42275_);
  and _54597_ (_03074_, _03073_, _03072_);
  or _54598_ (_03075_, _02898_, _41824_);
  or _54599_ (_03076_, _02900_, _41775_);
  and _54600_ (_03077_, _03076_, _03075_);
  and _54601_ (_03078_, _03077_, _03074_);
  and _54602_ (_03079_, _03078_, _03071_);
  or _54603_ (_03080_, _02907_, _42234_);
  or _54604_ (_03081_, _02910_, _42193_);
  and _54605_ (_03082_, _03081_, _03080_);
  or _54606_ (_03083_, _02913_, _41686_);
  or _54607_ (_03084_, _02915_, _41727_);
  and _54608_ (_03085_, _03084_, _03083_);
  and _54609_ (_03086_, _03085_, _03082_);
  or _54610_ (_03087_, _02919_, _42070_);
  or _54611_ (_03088_, _02921_, _42029_);
  and _54612_ (_03090_, _03088_, _03087_);
  or _54613_ (_03091_, _02924_, _41906_);
  or _54614_ (_03092_, _02926_, _41865_);
  and _54615_ (_03093_, _03092_, _03091_);
  and _54616_ (_03094_, _03093_, _03090_);
  and _54617_ (_03095_, _03094_, _03086_);
  nand _54618_ (_03096_, _03095_, _03079_);
  or _54619_ (_03097_, _03096_, _03063_);
  or _54620_ (_03098_, _02876_, _42157_);
  or _54621_ (_03099_, _02880_, _42116_);
  and _54622_ (_03101_, _03099_, _03098_);
  or _54623_ (_03102_, _02885_, _41993_);
  or _54624_ (_03103_, _02887_, _41952_);
  and _54625_ (_03104_, _03103_, _03102_);
  and _54626_ (_03105_, _03104_, _03101_);
  or _54627_ (_03106_, _02892_, _42321_);
  or _54628_ (_03107_, _02894_, _42280_);
  and _54629_ (_03108_, _03107_, _03106_);
  or _54630_ (_03109_, _02898_, _41829_);
  or _54631_ (_03110_, _02900_, _41780_);
  and _54632_ (_03112_, _03110_, _03109_);
  and _54633_ (_03113_, _03112_, _03108_);
  and _54634_ (_03114_, _03113_, _03105_);
  or _54635_ (_03115_, _02907_, _42239_);
  or _54636_ (_03116_, _02910_, _42198_);
  and _54637_ (_03117_, _03116_, _03115_);
  or _54638_ (_03118_, _02913_, _41691_);
  or _54639_ (_03119_, _02915_, _41732_);
  and _54640_ (_03120_, _03119_, _03118_);
  and _54641_ (_03121_, _03120_, _03117_);
  or _54642_ (_03123_, _02919_, _42075_);
  or _54643_ (_03124_, _02921_, _42034_);
  and _54644_ (_03125_, _03124_, _03123_);
  or _54645_ (_03126_, _02924_, _41911_);
  or _54646_ (_03127_, _02926_, _41870_);
  and _54647_ (_03128_, _03127_, _03126_);
  and _54648_ (_03129_, _03128_, _03125_);
  and _54649_ (_03130_, _03129_, _03121_);
  nand _54650_ (_03131_, _03130_, _03114_);
  or _54651_ (_03132_, _02876_, _42122_);
  or _54652_ (_03134_, _02880_, _42081_);
  and _54653_ (_03135_, _03134_, _03132_);
  or _54654_ (_03136_, _02885_, _41958_);
  or _54655_ (_03137_, _02887_, _41917_);
  and _54656_ (_03138_, _03137_, _03136_);
  and _54657_ (_03139_, _03138_, _03135_);
  or _54658_ (_03140_, _02892_, _42286_);
  or _54659_ (_03141_, _02894_, _42245_);
  and _54660_ (_03142_, _03141_, _03140_);
  or _54661_ (_03143_, _02898_, _41786_);
  or _54662_ (_03145_, _02900_, _41738_);
  and _54663_ (_03146_, _03145_, _03143_);
  and _54664_ (_03147_, _03146_, _03142_);
  and _54665_ (_03148_, _03147_, _03139_);
  or _54666_ (_03149_, _02907_, _42204_);
  or _54667_ (_03150_, _02910_, _42163_);
  and _54668_ (_03151_, _03150_, _03149_);
  or _54669_ (_03152_, _02913_, _41656_);
  or _54670_ (_03153_, _02915_, _41697_);
  and _54671_ (_03154_, _03153_, _03152_);
  and _54672_ (_03156_, _03154_, _03151_);
  or _54673_ (_03157_, _02919_, _42040_);
  or _54674_ (_03158_, _02921_, _41999_);
  and _54675_ (_03159_, _03158_, _03157_);
  or _54676_ (_03160_, _02924_, _41876_);
  or _54677_ (_03161_, _02926_, _41835_);
  and _54678_ (_03162_, _03161_, _03160_);
  and _54679_ (_03163_, _03162_, _03159_);
  and _54680_ (_03164_, _03163_, _03156_);
  and _54681_ (_03165_, _03164_, _03148_);
  or _54682_ (_03167_, _03165_, _03131_);
  nor _54683_ (_03168_, _03167_, _03097_);
  and _54684_ (_03169_, _03168_, _03030_);
  not _54685_ (_03170_, _03169_);
  and _54686_ (_03171_, _03165_, _03131_);
  and _54687_ (_03172_, _03062_, _03045_);
  and _54688_ (_03173_, _03095_, _03079_);
  or _54689_ (_03174_, _03173_, _03172_);
  not _54690_ (_03175_, _03174_);
  and _54691_ (_03176_, _03175_, _03171_);
  and _54692_ (_03178_, _03176_, _03030_);
  or _54693_ (_03179_, _03173_, _03063_);
  not _54694_ (_03180_, _03179_);
  and _54695_ (_03181_, _03180_, _03171_);
  and _54696_ (_03182_, _03181_, _03030_);
  nor _54697_ (_03183_, _03182_, _03178_);
  and _54698_ (_03184_, _03183_, _03170_);
  and _54699_ (_03185_, _03130_, _03114_);
  and _54700_ (_03186_, _03165_, _03185_);
  and _54701_ (_03187_, _03175_, _03186_);
  and _54702_ (_03188_, _03187_, _03030_);
  or _54703_ (_03189_, _03096_, _03172_);
  not _54704_ (_03190_, _03189_);
  and _54705_ (_03191_, _03171_, _03190_);
  and _54706_ (_03192_, _03191_, _03030_);
  nor _54707_ (_03193_, _03192_, _03188_);
  not _54708_ (_03194_, _03097_);
  and _54709_ (_03195_, _03194_, _03186_);
  and _54710_ (_03196_, _03195_, _03030_);
  and _54711_ (_03197_, _03190_, _03186_);
  and _54712_ (_03198_, _03030_, _03197_);
  nor _54713_ (_03199_, _03198_, _03196_);
  and _54714_ (_03200_, _03171_, _03194_);
  and _54715_ (_03201_, _03200_, _03030_);
  and _54716_ (_03202_, _03180_, _03186_);
  and _54717_ (_03203_, _03202_, _03030_);
  nor _54718_ (_03204_, _03203_, _03201_);
  and _54719_ (_03205_, _03204_, _03199_);
  and _54720_ (_03206_, _03205_, _03193_);
  and _54721_ (_03207_, _03206_, _03184_);
  and _54722_ (_03208_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _54723_ (_03209_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _54724_ (_03210_, _03209_, _03208_);
  or _54725_ (_03211_, _03210_, _03207_);
  not _54726_ (_03212_, _03168_);
  not _54727_ (_03213_, _03027_);
  or _54728_ (_03214_, _03213_, _02994_);
  or _54729_ (_03215_, _03214_, _02963_);
  nor _54730_ (_03216_, _03215_, _03212_);
  not _54731_ (_03217_, _03216_);
  not _54732_ (_03218_, _03028_);
  not _54733_ (_03219_, _02962_);
  and _54734_ (_03220_, _03219_, _02931_);
  and _54735_ (_03221_, _03220_, _03218_);
  and _54736_ (_03222_, _03221_, _03168_);
  nor _54737_ (_03223_, _03167_, _03189_);
  and _54738_ (_03224_, _03223_, _03030_);
  nor _54739_ (_03225_, _03224_, _03222_);
  or _54740_ (_03226_, _03167_, _03174_);
  or _54741_ (_03227_, _03226_, _03029_);
  or _54742_ (_03228_, _03165_, _03185_);
  or _54743_ (_03229_, _03228_, _03189_);
  or _54744_ (_03230_, _03229_, _03029_);
  and _54745_ (_03231_, _03230_, _03227_);
  or _54746_ (_03232_, _03228_, _03097_);
  or _54747_ (_03233_, _03232_, _03029_);
  or _54748_ (_03234_, _03228_, _03179_);
  or _54749_ (_03235_, _03234_, _03029_);
  and _54750_ (_03236_, _03235_, _03233_);
  or _54751_ (_03237_, _03167_, _03179_);
  or _54752_ (_03238_, _03237_, _03029_);
  or _54753_ (_03239_, _03228_, _03174_);
  or _54754_ (_03240_, _03239_, _03029_);
  and _54755_ (_03241_, _03240_, _03238_);
  and _54756_ (_03242_, _03241_, _03236_);
  and _54757_ (_03243_, _03242_, _03231_);
  and _54758_ (_03244_, _03243_, _03225_);
  not _54759_ (_03245_, _03210_);
  or _54760_ (_03246_, _03245_, _03244_);
  not _54761_ (_03247_, _03223_);
  or _54762_ (_03248_, _03247_, _03215_);
  and _54763_ (_03249_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and _54764_ (_03250_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _54765_ (_03251_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _54766_ (_03252_, _03251_, _03249_);
  and _54767_ (_03253_, _03252_, _03250_);
  nor _54768_ (_03254_, _03253_, _03249_);
  and _54769_ (_03255_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _54770_ (_03256_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _54771_ (_03257_, _03256_, _03255_);
  not _54772_ (_03258_, _03257_);
  nor _54773_ (_03259_, _03258_, _03254_);
  and _54774_ (_03260_, _03258_, _03254_);
  nor _54775_ (_03261_, _03260_, _03259_);
  not _54776_ (_03262_, _03261_);
  or _54777_ (_03263_, _03262_, _03248_);
  nor _54778_ (_03264_, _02873_, _02883_);
  and _54779_ (_03265_, _02873_, _02883_);
  nor _54780_ (_03266_, _03265_, _03264_);
  and _54781_ (_03267_, _03266_, _03248_);
  nand _54782_ (_03269_, _03267_, _03243_);
  nand _54783_ (_03270_, _03269_, _03263_);
  nand _54784_ (_03271_, _03270_, _03225_);
  nand _54785_ (_03272_, _03271_, _03246_);
  nand _54786_ (_03273_, _03272_, _03217_);
  not _54787_ (_03274_, \oc8051_golden_model_1.ACC [1]);
  and _54788_ (_03275_, _02906_, _02879_);
  nor _54789_ (_03276_, _03275_, _03274_);
  and _54790_ (_03277_, \oc8051_golden_model_1.ACC [0], _02905_);
  and _54791_ (_03278_, _03275_, _03274_);
  nor _54792_ (_03279_, _03278_, _03276_);
  and _54793_ (_03280_, _03279_, _03277_);
  nor _54794_ (_03281_, _03280_, _03276_);
  and _54795_ (_03282_, _03266_, \oc8051_golden_model_1.ACC [2]);
  nor _54796_ (_03283_, _03266_, \oc8051_golden_model_1.ACC [2]);
  nor _54797_ (_03284_, _03283_, _03282_);
  not _54798_ (_03285_, _03284_);
  nor _54799_ (_03286_, _03285_, _03281_);
  and _54800_ (_03287_, _03285_, _03281_);
  nor _54801_ (_03288_, _03287_, _03286_);
  and _54802_ (_03289_, _03288_, _03216_);
  not _54803_ (_03290_, _03289_);
  and _54804_ (_03291_, _03290_, _03207_);
  nand _54805_ (_03292_, _03291_, _03273_);
  nand _54806_ (_03293_, _03292_, _03211_);
  and _54807_ (_03294_, _03244_, _03207_);
  nor _54808_ (_03295_, _02891_, _02878_);
  nor _54809_ (_03296_, _03208_, \oc8051_golden_model_1.PC [3]);
  nor _54810_ (_03297_, _03296_, _03295_);
  or _54811_ (_03298_, _03297_, _03294_);
  and _54812_ (_03299_, _03225_, _03217_);
  nor _54813_ (_03300_, _03259_, _03255_);
  and _54814_ (_03301_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _54815_ (_03302_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _54816_ (_03303_, _03302_, _03301_);
  not _54817_ (_03304_, _03303_);
  nor _54818_ (_03305_, _03304_, _03300_);
  and _54819_ (_03306_, _03304_, _03300_);
  nor _54820_ (_03307_, _03306_, _03305_);
  or _54821_ (_03308_, _03307_, _03248_);
  not _54822_ (_03309_, _02885_);
  nor _54823_ (_03310_, _03264_, _02874_);
  nor _54824_ (_03311_, _03310_, _03309_);
  and _54825_ (_03312_, _03248_, _03311_);
  nand _54826_ (_03313_, _03312_, _03243_);
  nand _54827_ (_03314_, _03313_, _03308_);
  and _54828_ (_03315_, _03314_, _03299_);
  nor _54829_ (_03316_, _03286_, _03282_);
  nor _54830_ (_03317_, _03311_, \oc8051_golden_model_1.ACC [3]);
  and _54831_ (_03318_, _03311_, \oc8051_golden_model_1.ACC [3]);
  nor _54832_ (_03319_, _03318_, _03317_);
  and _54833_ (_03320_, _03319_, _03316_);
  nor _54834_ (_03321_, _03319_, _03316_);
  nor _54835_ (_03322_, _03321_, _03320_);
  nor _54836_ (_03323_, _03322_, _03217_);
  or _54837_ (_03324_, _03323_, _03315_);
  nand _54838_ (_03325_, _03324_, _03207_);
  and _54839_ (_03326_, _03325_, _03298_);
  or _54840_ (_03327_, _03326_, _03293_);
  nor _54841_ (_03328_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _54842_ (_03329_, _03328_, _03250_);
  or _54843_ (_03330_, _03329_, _03248_);
  and _54844_ (_03331_, _03248_, \oc8051_golden_model_1.PC [0]);
  nand _54845_ (_03332_, _03331_, _03243_);
  nand _54846_ (_03333_, _03332_, _03330_);
  and _54847_ (_03334_, _03333_, _03299_);
  not _54848_ (_03335_, \oc8051_golden_model_1.ACC [0]);
  and _54849_ (_03336_, _03335_, \oc8051_golden_model_1.PC [0]);
  nor _54850_ (_03337_, _03336_, _03277_);
  nor _54851_ (_03338_, _03337_, _03217_);
  or _54852_ (_03339_, _03338_, _03334_);
  nand _54853_ (_03340_, _03339_, _03207_);
  or _54854_ (_03341_, _03294_, \oc8051_golden_model_1.PC [0]);
  and _54855_ (_03342_, _03341_, _03340_);
  or _54856_ (_03343_, _03294_, _02878_);
  nor _54857_ (_03344_, _03252_, _03250_);
  nor _54858_ (_03345_, _03344_, _03253_);
  or _54859_ (_03346_, _03345_, _03248_);
  and _54860_ (_03347_, _03275_, _03248_);
  nand _54861_ (_03348_, _03347_, _03243_);
  nand _54862_ (_03349_, _03348_, _03346_);
  and _54863_ (_03350_, _03349_, _03299_);
  nor _54864_ (_03351_, _03279_, _03277_);
  nor _54865_ (_03352_, _03351_, _03280_);
  nor _54866_ (_03353_, _03352_, _03217_);
  or _54867_ (_03354_, _03353_, _03350_);
  nand _54868_ (_03355_, _03354_, _03207_);
  nand _54869_ (_03356_, _03355_, _03343_);
  or _54870_ (_03357_, _03356_, _03342_);
  or _54871_ (_03358_, _03357_, _03327_);
  nor _54872_ (_03359_, _03358_, _41927_);
  nand _54873_ (_03360_, _03341_, _03340_);
  and _54874_ (_03361_, _03355_, _03343_);
  or _54875_ (_03362_, _03361_, _03360_);
  or _54876_ (_03363_, _03362_, _03327_);
  nor _54877_ (_03364_, _03363_, _41886_);
  nor _54878_ (_03365_, _03364_, _03359_);
  or _54879_ (_03366_, _03356_, _03360_);
  and _54880_ (_03367_, _03292_, _03211_);
  nand _54881_ (_03368_, _03325_, _03298_);
  or _54882_ (_03369_, _03368_, _03367_);
  or _54883_ (_03370_, _03369_, _03366_);
  nor _54884_ (_03371_, _03370_, _42132_);
  or _54885_ (_03372_, _03326_, _03367_);
  or _54886_ (_03373_, _03361_, _03342_);
  or _54887_ (_03374_, _03373_, _03372_);
  nor _54888_ (_03375_, _03374_, _41666_);
  nor _54889_ (_03376_, _03375_, _03371_);
  and _54890_ (_03377_, _03376_, _03365_);
  or _54891_ (_03378_, _03369_, _03357_);
  nor _54892_ (_03379_, _03378_, _42091_);
  or _54893_ (_03380_, _03369_, _03362_);
  nor _54894_ (_03381_, _03380_, _42050_);
  nor _54895_ (_03382_, _03381_, _03379_);
  or _54896_ (_03383_, _03368_, _03293_);
  or _54897_ (_03384_, _03383_, _03357_);
  nor _54898_ (_03385_, _03384_, _42255_);
  or _54899_ (_03386_, _03372_, _03366_);
  nor _54900_ (_03387_, _03386_, _41801_);
  nor _54901_ (_03388_, _03387_, _03385_);
  and _54902_ (_03389_, _03388_, _03382_);
  and _54903_ (_03390_, _03389_, _03377_);
  or _54904_ (_03391_, _03383_, _03366_);
  nor _54905_ (_03392_, _03391_, _42296_);
  or _54906_ (_03393_, _03373_, _03383_);
  nor _54907_ (_03394_, _03393_, _42173_);
  nor _54908_ (_03395_, _03394_, _03392_);
  or _54909_ (_03396_, _03327_, _03366_);
  nor _54910_ (_03397_, _03396_, _41968_);
  or _54911_ (_03398_, _03373_, _03327_);
  nor _54912_ (_03399_, _03398_, _41845_);
  nor _54913_ (_03400_, _03399_, _03397_);
  and _54914_ (_03401_, _03400_, _03395_);
  or _54915_ (_03402_, _03369_, _03373_);
  nor _54916_ (_03403_, _03402_, _42009_);
  or _54917_ (_03404_, _03357_, _03372_);
  nor _54918_ (_03405_, _03404_, _41749_);
  nor _54919_ (_03406_, _03405_, _03403_);
  or _54920_ (_03407_, _03362_, _03383_);
  nor _54921_ (_03408_, _03407_, _42214_);
  or _54922_ (_03409_, _03362_, _03372_);
  nor _54923_ (_03410_, _03409_, _41707_);
  nor _54924_ (_03411_, _03410_, _03408_);
  and _54925_ (_03412_, _03411_, _03406_);
  and _54926_ (_03413_, _03412_, _03401_);
  and _54927_ (_03414_, _03413_, _03390_);
  not _54928_ (_03415_, _03414_);
  or _54929_ (_03416_, _03396_, _41958_);
  or _54930_ (_03417_, _03386_, _41786_);
  and _54931_ (_03418_, _03417_, _03416_);
  or _54932_ (_03419_, _03384_, _42245_);
  or _54933_ (_03420_, _03393_, _42163_);
  and _54934_ (_03421_, _03420_, _03419_);
  and _54935_ (_03422_, _03421_, _03418_);
  or _54936_ (_03423_, _03358_, _41917_);
  or _54937_ (_03424_, _03363_, _41876_);
  and _54938_ (_03425_, _03424_, _03423_);
  or _54939_ (_03426_, _03374_, _41656_);
  or _54940_ (_03427_, _03404_, _41738_);
  and _54941_ (_03428_, _03427_, _03426_);
  and _54942_ (_03429_, _03428_, _03425_);
  and _54943_ (_03430_, _03429_, _03422_);
  or _54944_ (_03431_, _03378_, _42081_);
  or _54945_ (_03432_, _03402_, _41999_);
  and _54946_ (_03433_, _03432_, _03431_);
  or _54947_ (_03434_, _03391_, _42286_);
  or _54948_ (_03435_, _03407_, _42204_);
  and _54949_ (_03436_, _03435_, _03434_);
  and _54950_ (_03437_, _03436_, _03433_);
  or _54951_ (_03438_, _03398_, _41835_);
  or _54952_ (_03439_, _03409_, _41697_);
  and _54953_ (_03440_, _03439_, _03438_);
  or _54954_ (_03441_, _03370_, _42122_);
  or _54955_ (_03442_, _03380_, _42040_);
  and _54956_ (_03443_, _03442_, _03441_);
  and _54957_ (_03444_, _03443_, _03440_);
  and _54958_ (_03445_, _03444_, _03437_);
  and _54959_ (_03446_, _03445_, _03430_);
  and _54960_ (_03447_, _03221_, _03195_);
  and _54961_ (_03448_, _03447_, _03446_);
  and _54962_ (_03449_, _03448_, _03415_);
  not _54963_ (_03450_, _02963_);
  and _54964_ (_03451_, _03213_, _02994_);
  and _54965_ (_03452_, _03451_, _03450_);
  and _54966_ (_03453_, _03452_, _03197_);
  not _54967_ (_03454_, _03446_);
  nor _54968_ (_03455_, _03358_, _41942_);
  nor _54969_ (_03456_, _03363_, _41901_);
  nor _54970_ (_03457_, _03456_, _03455_);
  nor _54971_ (_03458_, _03391_, _42311_);
  nor _54972_ (_03459_, _03370_, _42147_);
  nor _54973_ (_03460_, _03459_, _03458_);
  and _54974_ (_03461_, _03460_, _03457_);
  nor _54975_ (_03462_, _03384_, _42270_);
  nor _54976_ (_03463_, _03407_, _42229_);
  nor _54977_ (_03464_, _03463_, _03462_);
  nor _54978_ (_03465_, _03378_, _42106_);
  nor _54979_ (_03466_, _03402_, _42024_);
  nor _54980_ (_03467_, _03466_, _03465_);
  and _54981_ (_03468_, _03467_, _03464_);
  and _54982_ (_03470_, _03468_, _03461_);
  nor _54983_ (_03471_, _03374_, _41681_);
  nor _54984_ (_03472_, _03404_, _41770_);
  nor _54985_ (_03473_, _03472_, _03471_);
  nor _54986_ (_03474_, _03396_, _41983_);
  nor _54987_ (_03475_, _03398_, _41860_);
  nor _54988_ (_03476_, _03475_, _03474_);
  and _54989_ (_03477_, _03476_, _03473_);
  nor _54990_ (_03478_, _03393_, _42188_);
  nor _54991_ (_03479_, _03380_, _42065_);
  nor _54992_ (_03480_, _03479_, _03478_);
  nor _54993_ (_03481_, _03386_, _41819_);
  nor _54994_ (_03482_, _03409_, _41722_);
  nor _54995_ (_03483_, _03482_, _03481_);
  and _54996_ (_03484_, _03483_, _03480_);
  and _54997_ (_03485_, _03484_, _03477_);
  and _54998_ (_03486_, _03485_, _03470_);
  nor _54999_ (_03487_, _03486_, _03454_);
  and _55000_ (_03488_, _03487_, _03453_);
  and _55001_ (_03489_, _02962_, _02931_);
  and _55002_ (_03490_, _03489_, _03213_);
  and _55003_ (_03491_, _03490_, _03197_);
  not _55004_ (_03492_, _03491_);
  nor _55005_ (_03493_, _03219_, _02931_);
  and _55006_ (_03494_, _03493_, _03213_);
  and _55007_ (_03495_, _03494_, _03197_);
  not _55008_ (_03496_, \oc8051_golden_model_1.SP [1]);
  and _55009_ (_03497_, _03496_, \oc8051_golden_model_1.SP [0]);
  not _55010_ (_03498_, \oc8051_golden_model_1.SP [0]);
  and _55011_ (_03499_, \oc8051_golden_model_1.SP [1], _03498_);
  nor _55012_ (_03500_, _03499_, _03497_);
  not _55013_ (_03501_, _03500_);
  and _55014_ (_03502_, _03501_, _03188_);
  and _55015_ (_03503_, _03027_, _02994_);
  and _55016_ (_03504_, _03503_, _03450_);
  and _55017_ (_03505_, _03504_, _03223_);
  and _55018_ (_03506_, _03487_, _03505_);
  not _55019_ (_03507_, _03232_);
  and _55020_ (_03508_, _03507_, _03452_);
  and _55021_ (_03509_, _03501_, _03508_);
  not _55022_ (_03510_, _03508_);
  nand _55023_ (_03511_, _03220_, _03027_);
  nor _55024_ (_03512_, _03511_, _03239_);
  not _55025_ (_03513_, _03240_);
  not _55026_ (_03514_, _03447_);
  and _55027_ (_03515_, _03504_, _03202_);
  not _55028_ (_03516_, _03515_);
  and _55029_ (_03517_, _03221_, _03202_);
  not _55030_ (_03518_, _03517_);
  nor _55031_ (_03519_, _03396_, _41993_);
  nor _55032_ (_03520_, _03409_, _41732_);
  nor _55033_ (_03521_, _03520_, _03519_);
  nor _55034_ (_03522_, _03402_, _42034_);
  nor _55035_ (_03523_, _03386_, _41829_);
  nor _55036_ (_03524_, _03523_, _03522_);
  and _55037_ (_03525_, _03524_, _03521_);
  nor _55038_ (_03526_, _03370_, _42157_);
  nor _55039_ (_03527_, _03374_, _41691_);
  nor _55040_ (_03528_, _03527_, _03526_);
  nor _55041_ (_03529_, _03407_, _42239_);
  nor _55042_ (_03530_, _03393_, _42198_);
  nor _55043_ (_03531_, _03530_, _03529_);
  and _55044_ (_03532_, _03531_, _03528_);
  and _55045_ (_03533_, _03532_, _03525_);
  nor _55046_ (_03534_, _03384_, _42280_);
  nor _55047_ (_03535_, _03404_, _41780_);
  nor _55048_ (_03536_, _03535_, _03534_);
  nor _55049_ (_03537_, _03380_, _42075_);
  nor _55050_ (_03538_, _03358_, _41952_);
  nor _55051_ (_03539_, _03538_, _03537_);
  and _55052_ (_03540_, _03539_, _03536_);
  nor _55053_ (_03541_, _03378_, _42116_);
  nor _55054_ (_03542_, _03398_, _41870_);
  nor _55055_ (_03543_, _03542_, _03541_);
  nor _55056_ (_03544_, _03391_, _42321_);
  nor _55057_ (_03545_, _03363_, _41911_);
  nor _55058_ (_03546_, _03545_, _03544_);
  and _55059_ (_03547_, _03546_, _03543_);
  and _55060_ (_03548_, _03547_, _03540_);
  and _55061_ (_03549_, _03548_, _03533_);
  nor _55062_ (_03550_, _03549_, _03454_);
  or _55063_ (_03551_, _03391_, _42306_);
  or _55064_ (_03552_, _03402_, _42019_);
  and _55065_ (_03553_, _03552_, _03551_);
  or _55066_ (_03554_, _03378_, _42101_);
  or _55067_ (_03555_, _03386_, _41814_);
  and _55068_ (_03556_, _03555_, _03554_);
  and _55069_ (_03557_, _03556_, _03553_);
  or _55070_ (_03558_, _03384_, _42265_);
  or _55071_ (_03559_, _03407_, _42224_);
  and _55072_ (_03560_, _03559_, _03558_);
  or _55073_ (_03561_, _03396_, _41978_);
  or _55074_ (_03562_, _03398_, _41855_);
  and _55075_ (_03563_, _03562_, _03561_);
  and _55076_ (_03564_, _03563_, _03560_);
  and _55077_ (_03565_, _03564_, _03557_);
  or _55078_ (_03566_, _03363_, _41896_);
  or _55079_ (_03567_, _03404_, _41765_);
  and _55080_ (_03568_, _03567_, _03566_);
  or _55081_ (_03569_, _03374_, _41676_);
  or _55082_ (_03570_, _03409_, _41717_);
  and _55083_ (_03571_, _03570_, _03569_);
  and _55084_ (_03572_, _03571_, _03568_);
  or _55085_ (_03573_, _03393_, _42183_);
  or _55086_ (_03574_, _03358_, _41937_);
  and _55087_ (_03575_, _03574_, _03573_);
  or _55088_ (_03576_, _03370_, _42142_);
  or _55089_ (_03577_, _03380_, _42060_);
  and _55090_ (_03578_, _03577_, _03576_);
  and _55091_ (_03579_, _03578_, _03575_);
  and _55092_ (_03580_, _03579_, _03572_);
  and _55093_ (_03581_, _03580_, _03565_);
  nor _55094_ (_03582_, _03581_, _03446_);
  nor _55095_ (_03583_, _03582_, _03550_);
  and _55096_ (_03584_, _03504_, _03176_);
  and _55097_ (_03585_, _03504_, _03168_);
  nor _55098_ (_03586_, _03585_, _03584_);
  not _55099_ (_03587_, _03586_);
  and _55100_ (_03588_, _03587_, _03583_);
  not _55101_ (_03589_, _03222_);
  not _55102_ (_03590_, _03226_);
  and _55103_ (_03591_, _03489_, _03503_);
  and _55104_ (_03592_, _03489_, _03218_);
  or _55105_ (_03593_, _03592_, _03591_);
  and _55106_ (_03594_, _03593_, _03590_);
  and _55107_ (_03595_, _03489_, _03451_);
  nor _55108_ (_03596_, _03493_, _03595_);
  nor _55109_ (_03597_, _03596_, _03226_);
  nor _55110_ (_03598_, _03597_, _03594_);
  not _55111_ (_03599_, _03215_);
  and _55112_ (_03600_, _03599_, _03181_);
  and _55113_ (_03601_, _03221_, _03176_);
  nor _55114_ (_03602_, _03601_, _03600_);
  and _55115_ (_03603_, _03220_, _03451_);
  and _55116_ (_03604_, _03603_, _03590_);
  and _55117_ (_03605_, _03503_, _03220_);
  and _55118_ (_03606_, _03605_, _03590_);
  nor _55119_ (_03607_, _03606_, _03604_);
  and _55120_ (_03608_, _03607_, _03602_);
  not _55121_ (_03609_, _03229_);
  and _55122_ (_03610_, _03609_, _03221_);
  not _55123_ (_03611_, _03214_);
  and _55124_ (_03612_, _03489_, _03611_);
  and _55125_ (_03613_, _03612_, _03590_);
  nor _55126_ (_03614_, _03613_, _03610_);
  and _55127_ (_03615_, _03590_, _03221_);
  and _55128_ (_03616_, _03220_, _03611_);
  and _55129_ (_03617_, _03616_, _03590_);
  nor _55130_ (_03618_, _03617_, _03615_);
  and _55131_ (_03619_, _03618_, _03614_);
  and _55132_ (_03620_, _03619_, _03608_);
  and _55133_ (_03621_, _03187_, _03452_);
  and _55134_ (_03622_, _03599_, _03191_);
  nor _55135_ (_03623_, _03622_, _03621_);
  and _55136_ (_03624_, _03599_, _03200_);
  and _55137_ (_03625_, _03223_, _03452_);
  nor _55138_ (_03626_, _03625_, _03624_);
  and _55139_ (_03627_, _03626_, _03623_);
  and _55140_ (_03628_, _03202_, _03452_);
  and _55141_ (_03629_, _03504_, _03197_);
  nor _55142_ (_03630_, _03629_, _03628_);
  and _55143_ (_03631_, _03504_, _03195_);
  nor _55144_ (_03632_, _03631_, _03453_);
  and _55145_ (_03633_, _03632_, _03630_);
  and _55146_ (_03634_, _03633_, _03627_);
  and _55147_ (_03635_, _03634_, _03620_);
  and _55148_ (_03636_, _03635_, _03598_);
  and _55149_ (_03637_, _03636_, _02905_);
  nor _55150_ (_03638_, _03637_, \oc8051_golden_model_1.PC [1]);
  and _55151_ (_03639_, _03637_, \oc8051_golden_model_1.PC [1]);
  nor _55152_ (_03640_, _03639_, _03638_);
  nor _55153_ (_03641_, _03636_, _02905_);
  nor _55154_ (_03642_, _03641_, _03637_);
  nor _55155_ (_03643_, _03642_, _03640_);
  nor _55156_ (_03644_, _03636_, _03245_);
  and _55157_ (_03645_, _03636_, _03266_);
  nor _55158_ (_03646_, _03645_, _03644_);
  not _55159_ (_03647_, _03646_);
  not _55160_ (_03648_, _03297_);
  nor _55161_ (_03649_, _03636_, _03648_);
  not _55162_ (_03650_, _03311_);
  and _55163_ (_03651_, _03636_, _03650_);
  nor _55164_ (_03652_, _03651_, _03649_);
  and _55165_ (_03653_, _03652_, _03647_);
  and _55166_ (_03654_, _03653_, _03643_);
  and _55167_ (_03655_, _03654_, _02025_);
  and _55168_ (_03656_, _03652_, _03646_);
  and _55169_ (_03657_, _03656_, _03643_);
  and _55170_ (_03658_, _03657_, _02056_);
  nor _55171_ (_03659_, _03658_, _03655_);
  nor _55172_ (_03660_, _03652_, _03646_);
  and _55173_ (_03661_, _03642_, _03640_);
  and _55174_ (_03662_, _03661_, _03660_);
  and _55175_ (_03663_, _03662_, _02070_);
  nor _55176_ (_03664_, _03652_, _03647_);
  and _55177_ (_03665_, _03664_, _03661_);
  and _55178_ (_03666_, _03665_, _02027_);
  nor _55179_ (_03667_, _03666_, _03663_);
  and _55180_ (_03668_, _03667_, _03659_);
  not _55181_ (_03669_, _03642_);
  nor _55182_ (_03671_, _03669_, _03640_);
  and _55183_ (_03672_, _03671_, _03653_);
  and _55184_ (_03673_, _03672_, _02042_);
  and _55185_ (_03674_, _03669_, _03640_);
  and _55186_ (_03675_, _03674_, _03653_);
  and _55187_ (_03676_, _03675_, _02048_);
  nor _55188_ (_03677_, _03676_, _03673_);
  and _55189_ (_03678_, _03661_, _03653_);
  and _55190_ (_03679_, _03678_, _02053_);
  and _55191_ (_03680_, _03661_, _03656_);
  and _55192_ (_03681_, _03680_, _02020_);
  nor _55193_ (_03682_, _03681_, _03679_);
  and _55194_ (_03683_, _03682_, _03677_);
  and _55195_ (_03684_, _03683_, _03668_);
  and _55196_ (_03685_, _03660_, _03643_);
  and _55197_ (_03686_, _03685_, _02058_);
  and _55198_ (_03687_, _03671_, _03660_);
  and _55199_ (_03688_, _03687_, _02068_);
  nor _55200_ (_03689_, _03688_, _03686_);
  and _55201_ (_03690_, _03674_, _03660_);
  and _55202_ (_03691_, _03690_, _02045_);
  and _55203_ (_03692_, _03664_, _03643_);
  and _55204_ (_03693_, _03692_, _02061_);
  nor _55205_ (_03694_, _03693_, _03691_);
  and _55206_ (_03695_, _03694_, _03689_);
  and _55207_ (_03696_, _03671_, _03664_);
  and _55208_ (_03697_, _03696_, _02030_);
  and _55209_ (_03698_, _03674_, _03664_);
  and _55210_ (_03699_, _03698_, _02032_);
  nor _55211_ (_03700_, _03699_, _03697_);
  and _55212_ (_03701_, _03671_, _03656_);
  and _55213_ (_03702_, _03701_, _02022_);
  and _55214_ (_03703_, _03674_, _03656_);
  and _55215_ (_03704_, _03703_, _02037_);
  nor _55216_ (_03705_, _03704_, _03702_);
  and _55217_ (_03706_, _03705_, _03700_);
  and _55218_ (_03707_, _03706_, _03695_);
  and _55219_ (_03708_, _03707_, _03684_);
  nor _55220_ (_03709_, _03708_, _03589_);
  not _55221_ (_03710_, _03505_);
  nor _55222_ (_03711_, _03615_, _03508_);
  nor _55223_ (_03712_, _03711_, _03581_);
  not _55224_ (_03713_, _03712_);
  and _55225_ (_03714_, _03504_, _03507_);
  and _55226_ (_03715_, _03504_, _03609_);
  or _55227_ (_03716_, _03715_, _03714_);
  and _55228_ (_03717_, _03716_, _03583_);
  and _55229_ (_03718_, _03590_, _03452_);
  and _55230_ (_03719_, _03504_, _03590_);
  nor _55231_ (_03720_, _03719_, _03718_);
  not _55232_ (_03721_, _03711_);
  not _55233_ (_03722_, \oc8051_golden_model_1.SP [3]);
  and _55234_ (_03723_, _03609_, _03452_);
  and _55235_ (_03724_, _03723_, _03722_);
  not _55236_ (_03725_, _03234_);
  and _55237_ (_03726_, _03725_, _03221_);
  nor _55238_ (_03727_, _03726_, _03610_);
  or _55239_ (_03728_, _03727_, _03581_);
  and _55240_ (_03729_, _03507_, _03221_);
  nor _55241_ (_03730_, _03723_, _03715_);
  nand _55242_ (_03731_, _03727_, \oc8051_golden_model_1.PSW [3]);
  and _55243_ (_03732_, _03731_, _03730_);
  or _55244_ (_03733_, _03732_, _03729_);
  and _55245_ (_03734_, _03733_, _03728_);
  or _55246_ (_03735_, _03734_, _03724_);
  not _55247_ (_03736_, _03714_);
  not _55248_ (_03737_, _03729_);
  or _55249_ (_03738_, _03737_, _03581_);
  and _55250_ (_03739_, _03738_, _03736_);
  and _55251_ (_03740_, _03739_, _03735_);
  or _55252_ (_03741_, _03740_, _03721_);
  and _55253_ (_03742_, _03741_, _03720_);
  or _55254_ (_03743_, _03742_, _03717_);
  and _55255_ (_03744_, _03743_, _03713_);
  nor _55256_ (_03745_, _03237_, _03219_);
  not _55257_ (_03746_, _03720_);
  and _55258_ (_03747_, _03746_, _03583_);
  nor _55259_ (_03748_, _03747_, _03745_);
  not _55260_ (_03749_, _03748_);
  nor _55261_ (_03750_, _03749_, _03744_);
  not _55262_ (_03751_, _03237_);
  and _55263_ (_03752_, _03751_, _03452_);
  and _55264_ (_03753_, _03504_, _03751_);
  nor _55265_ (_03754_, _03753_, _03752_);
  not _55266_ (_03755_, _03754_);
  not _55267_ (_03756_, _03581_);
  and _55268_ (_03757_, _03745_, _03756_);
  nor _55269_ (_03758_, _03757_, _03755_);
  not _55270_ (_03759_, _03758_);
  nor _55271_ (_03760_, _03759_, _03750_);
  and _55272_ (_03761_, _03223_, _03221_);
  and _55273_ (_03762_, _03755_, _03583_);
  nor _55274_ (_03763_, _03762_, _03761_);
  not _55275_ (_03764_, _03763_);
  nor _55276_ (_03765_, _03764_, _03760_);
  not _55277_ (_03766_, _03761_);
  nor _55278_ (_03767_, _03766_, _03581_);
  or _55279_ (_03768_, _03767_, _03765_);
  and _55280_ (_03769_, _03768_, _03710_);
  nor _55281_ (_03770_, _03583_, _03710_);
  or _55282_ (_03771_, _03770_, _03769_);
  and _55283_ (_03772_, _03771_, _03589_);
  or _55284_ (_03773_, _03772_, _03587_);
  nor _55285_ (_03774_, _03773_, _03709_);
  nor _55286_ (_03775_, _03774_, _03588_);
  and _55287_ (_03776_, _03221_, _03187_);
  not _55288_ (_03777_, _03776_);
  and _55289_ (_03778_, _03221_, _03181_);
  not _55290_ (_03779_, _03778_);
  and _55291_ (_03780_, _03504_, _03181_);
  nor _55292_ (_03781_, _03780_, _03600_);
  and _55293_ (_03782_, _03781_, _03779_);
  and _55294_ (_03783_, _03221_, _03200_);
  not _55295_ (_03784_, _03783_);
  and _55296_ (_03785_, _03504_, _03200_);
  nor _55297_ (_03786_, _03785_, _03624_);
  and _55298_ (_03787_, _03786_, _03784_);
  and _55299_ (_03788_, _03221_, _03191_);
  not _55300_ (_03789_, _03788_);
  and _55301_ (_03790_, _03504_, _03191_);
  nor _55302_ (_03791_, _03790_, _03622_);
  and _55303_ (_03792_, _03791_, _03789_);
  and _55304_ (_03793_, _03792_, _03787_);
  and _55305_ (_03794_, _03793_, _03782_);
  and _55306_ (_03795_, _03794_, _03777_);
  not _55307_ (_03796_, _03795_);
  nor _55308_ (_03797_, _03796_, _03775_);
  and _55309_ (_03798_, _03504_, _03187_);
  and _55310_ (_03799_, _03796_, _03581_);
  nor _55311_ (_03800_, _03799_, _03798_);
  not _55312_ (_03801_, _03800_);
  nor _55313_ (_03802_, _03801_, _03797_);
  and _55314_ (_03803_, _03798_, \oc8051_golden_model_1.SP [3]);
  or _55315_ (_03804_, _03803_, _03621_);
  nor _55316_ (_03805_, _03804_, _03802_);
  and _55317_ (_03806_, _03583_, _03621_);
  or _55318_ (_03807_, _03806_, _03805_);
  and _55319_ (_03808_, _03807_, _03518_);
  and _55320_ (_03809_, _03517_, _03581_);
  or _55321_ (_03810_, _03809_, _03808_);
  nand _55322_ (_03811_, _03810_, _03516_);
  and _55323_ (_03812_, _03515_, _03722_);
  nor _55324_ (_03813_, _03812_, _03628_);
  nand _55325_ (_03814_, _03813_, _03811_);
  and _55326_ (_03815_, _03221_, _03197_);
  not _55327_ (_03816_, _03628_);
  nor _55328_ (_03817_, _03816_, _03583_);
  nor _55329_ (_03818_, _03817_, _03815_);
  nand _55330_ (_03819_, _03818_, _03814_);
  and _55331_ (_03820_, _03815_, _03581_);
  nor _55332_ (_03821_, _03820_, _03453_);
  and _55333_ (_03822_, _03821_, _03819_);
  not _55334_ (_03823_, _03453_);
  nor _55335_ (_03824_, _03583_, _03823_);
  or _55336_ (_03825_, _03824_, _03822_);
  nand _55337_ (_03826_, _03825_, _03514_);
  nor _55338_ (_03827_, _03514_, _03581_);
  not _55339_ (_03828_, _03827_);
  and _55340_ (_03829_, _03828_, _03826_);
  nor _55341_ (_03830_, _03391_, _42316_);
  nor _55342_ (_03831_, _03370_, _42152_);
  nor _55343_ (_03832_, _03831_, _03830_);
  nor _55344_ (_03833_, _03363_, _41906_);
  nor _55345_ (_03834_, _03374_, _41686_);
  nor _55346_ (_03835_, _03834_, _03833_);
  and _55347_ (_03836_, _03835_, _03832_);
  nor _55348_ (_03837_, _03378_, _42111_);
  nor _55349_ (_03838_, _03380_, _42070_);
  nor _55350_ (_03839_, _03838_, _03837_);
  nor _55351_ (_03840_, _03384_, _42275_);
  nor _55352_ (_03841_, _03393_, _42193_);
  nor _55353_ (_03842_, _03841_, _03840_);
  and _55354_ (_03843_, _03842_, _03839_);
  and _55355_ (_03844_, _03843_, _03836_);
  nor _55356_ (_03845_, _03386_, _41824_);
  nor _55357_ (_03846_, _03404_, _41775_);
  nor _55358_ (_03847_, _03846_, _03845_);
  nor _55359_ (_03848_, _03396_, _41988_);
  nor _55360_ (_03849_, _03409_, _41727_);
  nor _55361_ (_03850_, _03849_, _03848_);
  and _55362_ (_03851_, _03850_, _03847_);
  nor _55363_ (_03852_, _03407_, _42234_);
  nor _55364_ (_03853_, _03402_, _42029_);
  nor _55365_ (_03854_, _03853_, _03852_);
  nor _55366_ (_03855_, _03358_, _41947_);
  nor _55367_ (_03856_, _03398_, _41865_);
  nor _55368_ (_03857_, _03856_, _03855_);
  and _55369_ (_03858_, _03857_, _03854_);
  and _55370_ (_03859_, _03858_, _03851_);
  and _55371_ (_03860_, _03859_, _03844_);
  nor _55372_ (_03861_, _03860_, _03454_);
  and _55373_ (_03862_, _03861_, _03715_);
  not _55374_ (_03863_, _03862_);
  not _55375_ (_03864_, _03861_);
  nor _55376_ (_03865_, _03621_, _03453_);
  and _55377_ (_03866_, _03865_, _03754_);
  and _55378_ (_03867_, _03866_, _03720_);
  nor _55379_ (_03868_, _03628_, _03714_);
  and _55380_ (_03869_, _03586_, _03710_);
  and _55381_ (_03870_, _03869_, _03868_);
  and _55382_ (_03872_, _03870_, _03867_);
  nor _55383_ (_03873_, _03872_, _03864_);
  nor _55384_ (_03874_, _03396_, _41973_);
  nor _55385_ (_03875_, _03386_, _41809_);
  nor _55386_ (_03876_, _03875_, _03874_);
  nor _55387_ (_03877_, _03393_, _42178_);
  nor _55388_ (_03878_, _03380_, _42055_);
  nor _55389_ (_03879_, _03878_, _03877_);
  and _55390_ (_03880_, _03879_, _03876_);
  nor _55391_ (_03881_, _03358_, _41932_);
  nor _55392_ (_03882_, _03363_, _41891_);
  nor _55393_ (_03883_, _03882_, _03881_);
  nor _55394_ (_03884_, _03404_, _41758_);
  nor _55395_ (_03885_, _03409_, _41712_);
  nor _55396_ (_03886_, _03885_, _03884_);
  and _55397_ (_03887_, _03886_, _03883_);
  and _55398_ (_03888_, _03887_, _03880_);
  nor _55399_ (_03889_, _03370_, _42137_);
  nor _55400_ (_03890_, _03378_, _42096_);
  nor _55401_ (_03891_, _03890_, _03889_);
  nor _55402_ (_03892_, _03391_, _42301_);
  nor _55403_ (_03893_, _03402_, _42014_);
  nor _55404_ (_03894_, _03893_, _03892_);
  and _55405_ (_03895_, _03894_, _03891_);
  nor _55406_ (_03896_, _03384_, _42260_);
  nor _55407_ (_03897_, _03407_, _42219_);
  nor _55408_ (_03898_, _03897_, _03896_);
  nor _55409_ (_03899_, _03398_, _41850_);
  nor _55410_ (_03900_, _03374_, _41671_);
  nor _55411_ (_03901_, _03900_, _03899_);
  and _55412_ (_03902_, _03901_, _03898_);
  and _55413_ (_03903_, _03902_, _03895_);
  and _55414_ (_03904_, _03903_, _03888_);
  nor _55415_ (_03905_, _03761_, _03745_);
  and _55416_ (_03906_, _03905_, _03737_);
  and _55417_ (_03907_, _03727_, _03711_);
  and _55418_ (_03908_, _03907_, _03906_);
  nor _55419_ (_03909_, _03815_, _03447_);
  and _55420_ (_03910_, _03909_, _03777_);
  and _55421_ (_03911_, _03910_, _03518_);
  and _55422_ (_03912_, _03911_, _03908_);
  and _55423_ (_03913_, _03912_, _03794_);
  nor _55424_ (_03914_, _03913_, _03904_);
  not _55425_ (_03915_, _03914_);
  and _55426_ (_03916_, _03690_, _01997_);
  and _55427_ (_03917_, _03654_, _01977_);
  nor _55428_ (_03918_, _03917_, _03916_);
  and _55429_ (_03919_, _03672_, _01992_);
  and _55430_ (_03920_, _03680_, _01965_);
  nor _55431_ (_03921_, _03920_, _03919_);
  and _55432_ (_03922_, _03921_, _03918_);
  and _55433_ (_03923_, _03692_, _02005_);
  and _55434_ (_03924_, _03657_, _01979_);
  nor _55435_ (_03925_, _03924_, _03923_);
  and _55436_ (_03926_, _03696_, _01972_);
  and _55437_ (_03927_, _03665_, _02000_);
  nor _55438_ (_03928_, _03927_, _03926_);
  and _55439_ (_03929_, _03928_, _03925_);
  and _55440_ (_03930_, _03929_, _03922_);
  and _55441_ (_03931_, _03675_, _01986_);
  and _55442_ (_03932_, _03678_, _02014_);
  nor _55443_ (_03933_, _03932_, _03931_);
  and _55444_ (_03934_, _03687_, _01989_);
  and _55445_ (_03935_, _03703_, _01970_);
  nor _55446_ (_03936_, _03935_, _03934_);
  and _55447_ (_03937_, _03936_, _03933_);
  and _55448_ (_03938_, _03685_, _02002_);
  and _55449_ (_03939_, _03701_, _01967_);
  nor _55450_ (_03940_, _03939_, _03938_);
  and _55451_ (_03941_, _03662_, _02012_);
  and _55452_ (_03942_, _03698_, _01974_);
  nor _55453_ (_03943_, _03942_, _03941_);
  and _55454_ (_03944_, _03943_, _03940_);
  and _55455_ (_03945_, _03944_, _03937_);
  and _55456_ (_03946_, _03945_, _03930_);
  nor _55457_ (_03947_, _03946_, _03589_);
  not _55458_ (_03948_, _03490_);
  not _55459_ (_03949_, _03202_);
  nor _55460_ (_03950_, _03590_, _03191_);
  and _55461_ (_03951_, _03950_, _03949_);
  nor _55462_ (_03952_, _03951_, _03948_);
  not _55463_ (_03953_, _03952_);
  and _55464_ (_03954_, _03489_, _03027_);
  not _55465_ (_03955_, _03954_);
  nor _55466_ (_03956_, _03590_, _03187_);
  and _55467_ (_03957_, _03956_, _03212_);
  nor _55468_ (_03958_, _03957_, _03955_);
  not _55469_ (_03959_, _03958_);
  and _55470_ (_03960_, _03489_, _03195_);
  not _55471_ (_03961_, _03960_);
  and _55472_ (_03962_, _03489_, _03609_);
  and _55473_ (_03963_, _03490_, _03181_);
  nor _55474_ (_03964_, _03963_, _03962_);
  and _55475_ (_03965_, _03964_, _03961_);
  and _55476_ (_03966_, _03965_, _03959_);
  and _55477_ (_03967_, _03966_, _03953_);
  and _55478_ (_03968_, _03592_, _03187_);
  and _55479_ (_03969_, _03595_, _03168_);
  nor _55480_ (_03970_, _03969_, _03968_);
  and _55481_ (_03971_, _03954_, _03200_);
  and _55482_ (_03972_, _03954_, _03197_);
  nor _55483_ (_03973_, _03972_, _03971_);
  nor _55484_ (_03974_, _03223_, _03181_);
  nor _55485_ (_03975_, _03974_, _03955_);
  not _55486_ (_03976_, _03975_);
  and _55487_ (_03977_, _03976_, _03973_);
  and _55488_ (_03978_, _03977_, _03970_);
  and _55489_ (_03979_, _03954_, _03725_);
  and _55490_ (_03980_, _03592_, _03725_);
  or _55491_ (_03981_, _03980_, _03979_);
  and _55492_ (_03982_, _03954_, _03191_);
  nor _55493_ (_03983_, _03982_, _03981_);
  and _55494_ (_03984_, _03490_, _03200_);
  and _55495_ (_03985_, _03489_, _03507_);
  nor _55496_ (_03986_, _03985_, _03984_);
  and _55497_ (_03987_, _03986_, _03983_);
  and _55498_ (_03988_, _03595_, _03223_);
  not _55499_ (_03989_, _03988_);
  and _55500_ (_03990_, _03954_, _03202_);
  nor _55501_ (_03991_, _03491_, _03990_);
  and _55502_ (_03992_, _03991_, _03989_);
  and _55503_ (_03993_, _03992_, _03987_);
  and _55504_ (_03994_, _03993_, _03978_);
  not _55505_ (_03995_, \oc8051_golden_model_1.SP [2]);
  not _55506_ (_03996_, _03723_);
  nor _55507_ (_03997_, _03798_, _03515_);
  and _55508_ (_03998_, _03997_, _03996_);
  nor _55509_ (_03999_, _03998_, _03995_);
  or _55510_ (_04000_, _03223_, _03168_);
  and _55511_ (_04001_, _04000_, _03592_);
  not _55512_ (_04002_, _04001_);
  and _55513_ (_04003_, _03595_, _03187_);
  and _55514_ (_04004_, _03595_, _03725_);
  nor _55515_ (_04005_, _04004_, _04003_);
  and _55516_ (_04006_, _04005_, _04002_);
  not _55517_ (_04007_, _04006_);
  nor _55518_ (_04008_, _04007_, _03999_);
  and _55519_ (_04009_, _04008_, _03994_);
  and _55520_ (_04010_, _04009_, _03967_);
  not _55521_ (_04011_, _04010_);
  nor _55522_ (_04012_, _04011_, _03947_);
  and _55523_ (_04013_, _04012_, _03915_);
  not _55524_ (_04014_, _04013_);
  nor _55525_ (_04015_, _04014_, _03873_);
  and _55526_ (_04016_, _04015_, _03863_);
  not _55527_ (_04017_, \oc8051_golden_model_1.IRAM[0] [1]);
  or _55528_ (_04018_, _03384_, _42250_);
  or _55529_ (_04019_, _03407_, _42209_);
  and _55530_ (_04020_, _04019_, _04018_);
  or _55531_ (_04021_, _03370_, _42127_);
  or _55532_ (_04022_, _03378_, _42086_);
  and _55533_ (_04023_, _04022_, _04021_);
  and _55534_ (_04024_, _04023_, _04020_);
  or _55535_ (_04025_, _03374_, _41661_);
  or _55536_ (_04026_, _03409_, _41702_);
  and _55537_ (_04027_, _04026_, _04025_);
  or _55538_ (_04028_, _03363_, _41881_);
  or _55539_ (_04029_, _03398_, _41840_);
  and _55540_ (_04030_, _04029_, _04028_);
  and _55541_ (_04031_, _04030_, _04027_);
  and _55542_ (_04032_, _04031_, _04024_);
  or _55543_ (_04033_, _03380_, _42045_);
  or _55544_ (_04034_, _03402_, _42004_);
  and _55545_ (_04035_, _04034_, _04033_);
  or _55546_ (_04036_, _03391_, _42291_);
  or _55547_ (_04037_, _03393_, _42168_);
  and _55548_ (_04038_, _04037_, _04036_);
  and _55549_ (_04039_, _04038_, _04035_);
  or _55550_ (_04040_, _03396_, _41963_);
  or _55551_ (_04041_, _03358_, _41922_);
  and _55552_ (_04042_, _04041_, _04040_);
  or _55553_ (_04043_, _03386_, _41791_);
  or _55554_ (_04044_, _03404_, _41743_);
  and _55555_ (_04045_, _04044_, _04043_);
  and _55556_ (_04046_, _04045_, _04042_);
  and _55557_ (_04047_, _04046_, _04039_);
  and _55558_ (_04048_, _04047_, _04032_);
  nor _55559_ (_04049_, _04048_, _03514_);
  not _55560_ (_04050_, _04049_);
  and _55561_ (_04051_, _03756_, _03446_);
  and _55562_ (_04052_, _04051_, _03453_);
  and _55563_ (_04053_, _03505_, _04051_);
  nor _55564_ (_04054_, _04048_, _03766_);
  not _55565_ (_04055_, _03715_);
  not _55566_ (_04056_, _03726_);
  nor _55567_ (_04057_, _04048_, _04056_);
  and _55568_ (_04058_, _03493_, _03451_);
  nor _55569_ (_04059_, _03605_, _04058_);
  nor _55570_ (_04060_, _04059_, _03234_);
  not _55571_ (_04061_, _04060_);
  not _55572_ (_04062_, _03239_);
  and _55573_ (_04063_, _03605_, _04062_);
  and _55574_ (_04064_, _03591_, _03725_);
  nor _55575_ (_04065_, _04064_, _04063_);
  and _55576_ (_04066_, _03493_, _03503_);
  and _55577_ (_04067_, _04066_, _03725_);
  not _55578_ (_04068_, _04067_);
  nor _55579_ (_04069_, _04004_, _03726_);
  and _55580_ (_04070_, _04069_, _04068_);
  and _55581_ (_04071_, _04070_, _04065_);
  and _55582_ (_04073_, _04071_, _04061_);
  or _55583_ (_04074_, _04073_, _04057_);
  and _55584_ (_04075_, _03489_, _02994_);
  nor _55585_ (_04076_, _04066_, _04075_);
  and _55586_ (_04077_, _04076_, _04059_);
  nor _55587_ (_04078_, _04077_, _03229_);
  nor _55588_ (_04079_, _04078_, _03610_);
  nand _55589_ (_04080_, _04079_, _04074_);
  not _55590_ (_04081_, _03610_);
  or _55591_ (_04082_, _04048_, _04081_);
  nand _55592_ (_04083_, _04082_, _04080_);
  nand _55593_ (_04084_, _04083_, _04055_);
  nand _55594_ (_04085_, _03715_, _04051_);
  nand _55595_ (_04086_, _04085_, _04084_);
  and _55596_ (_04087_, _03723_, _03498_);
  nor _55597_ (_04088_, _04087_, _03729_);
  not _55598_ (_04089_, _04088_);
  nor _55599_ (_04090_, _04077_, _03232_);
  nor _55600_ (_04091_, _04090_, _04089_);
  and _55601_ (_04092_, _04091_, _04086_);
  nor _55602_ (_04093_, _04048_, _03737_);
  or _55603_ (_04094_, _04093_, _04092_);
  and _55604_ (_04095_, _04094_, _03736_);
  and _55605_ (_04096_, _03714_, _04051_);
  or _55606_ (_04097_, _04096_, _04095_);
  and _55607_ (_04098_, _04048_, _03508_);
  nor _55608_ (_04099_, _03606_, _03615_);
  and _55609_ (_04100_, _02994_, _02962_);
  and _55610_ (_04101_, _04100_, _03590_);
  not _55611_ (_04102_, _04101_);
  and _55612_ (_04103_, _04102_, _04099_);
  not _55613_ (_04104_, _04103_);
  nor _55614_ (_04105_, _04104_, _04098_);
  and _55615_ (_04106_, _04105_, _04097_);
  not _55616_ (_04107_, _03615_);
  nor _55617_ (_04108_, _04048_, _04107_);
  or _55618_ (_04109_, _04108_, _04106_);
  nand _55619_ (_04110_, _04109_, _03720_);
  and _55620_ (_04111_, _03746_, _04051_);
  nor _55621_ (_04112_, _04111_, _03745_);
  nand _55622_ (_04113_, _04112_, _04110_);
  and _55623_ (_04114_, _04048_, _03745_);
  and _55624_ (_04115_, _03605_, _03751_);
  nor _55625_ (_04116_, _04115_, _03755_);
  not _55626_ (_04117_, _04116_);
  nor _55627_ (_04118_, _04117_, _04114_);
  and _55628_ (_04119_, _04118_, _04113_);
  and _55629_ (_04120_, _03755_, _04051_);
  nor _55630_ (_04121_, _04120_, _04119_);
  nor _55631_ (_04122_, _04066_, _03591_);
  nor _55632_ (_04123_, _03595_, _03221_);
  and _55633_ (_04124_, _04123_, _04059_);
  and _55634_ (_04125_, _04124_, _04122_);
  nor _55635_ (_04126_, _04125_, _03247_);
  nor _55636_ (_04127_, _04126_, _04121_);
  or _55637_ (_04128_, _04127_, _04054_);
  and _55638_ (_04129_, _04128_, _03710_);
  nor _55639_ (_04130_, _04129_, _04053_);
  nor _55640_ (_04131_, _04077_, _03212_);
  nor _55641_ (_04132_, _04131_, _04130_);
  and _55642_ (_04133_, _03665_, _01864_);
  and _55643_ (_04134_, _03678_, _01900_);
  nor _55644_ (_04135_, _04134_, _04133_);
  and _55645_ (_04136_, _03685_, _01890_);
  and _55646_ (_04137_, _03654_, _01888_);
  nor _55647_ (_04138_, _04137_, _04136_);
  and _55648_ (_04139_, _04138_, _04135_);
  and _55649_ (_04140_, _03698_, _01862_);
  and _55650_ (_04141_, _03675_, _01885_);
  nor _55651_ (_04142_, _04141_, _04140_);
  and _55652_ (_04143_, _03680_, _01869_);
  and _55653_ (_04144_, _03703_, _01871_);
  nor _55654_ (_04145_, _04144_, _04143_);
  and _55655_ (_04146_, _04145_, _04142_);
  and _55656_ (_04147_, _04146_, _04139_);
  and _55657_ (_04148_, _03662_, _01875_);
  and _55658_ (_04149_, _03692_, _01893_);
  nor _55659_ (_04150_, _04149_, _04148_);
  and _55660_ (_04151_, _03672_, _01877_);
  and _55661_ (_04152_, _03701_, _01853_);
  nor _55662_ (_04153_, _04152_, _04151_);
  and _55663_ (_04154_, _04153_, _04150_);
  and _55664_ (_04155_, _03690_, _01879_);
  and _55665_ (_04156_, _03696_, _01859_);
  nor _55666_ (_04157_, _04156_, _04155_);
  and _55667_ (_04158_, _03687_, _01902_);
  and _55668_ (_04159_, _03657_, _01856_);
  nor _55669_ (_04160_, _04159_, _04158_);
  and _55670_ (_04161_, _04160_, _04157_);
  and _55671_ (_04162_, _04161_, _04154_);
  and _55672_ (_04163_, _04162_, _04147_);
  and _55673_ (_04164_, _04163_, _03222_);
  nor _55674_ (_04165_, _04164_, _03585_);
  and _55675_ (_04166_, _04165_, _04132_);
  and _55676_ (_04167_, _03585_, _04051_);
  or _55677_ (_04168_, _04167_, _04166_);
  and _55678_ (_04169_, _03605_, _03176_);
  nor _55679_ (_04170_, _04169_, _03584_);
  and _55680_ (_04171_, _04170_, _04168_);
  and _55681_ (_04172_, _03584_, _04051_);
  or _55682_ (_04174_, _04172_, _04171_);
  not _55683_ (_04175_, _03181_);
  nor _55684_ (_04176_, _04058_, _03591_);
  nor _55685_ (_04177_, _04176_, _04175_);
  not _55686_ (_04178_, _04177_);
  and _55687_ (_04179_, _03963_, _02994_);
  not _55688_ (_04180_, _04179_);
  and _55689_ (_04181_, _04066_, _03181_);
  and _55690_ (_04182_, _03605_, _03181_);
  nor _55691_ (_04183_, _04182_, _04181_);
  and _55692_ (_04184_, _04183_, _04180_);
  and _55693_ (_04185_, _04184_, _04178_);
  and _55694_ (_04186_, _04185_, _04174_);
  and _55695_ (_04187_, _03792_, _03782_);
  not _55696_ (_04188_, _04048_);
  nor _55697_ (_04189_, _04188_, _04187_);
  not _55698_ (_04190_, _03200_);
  nor _55699_ (_04191_, _04077_, _04190_);
  not _55700_ (_04192_, _04191_);
  not _55701_ (_04193_, _03191_);
  nor _55702_ (_04194_, _03605_, _04075_);
  nor _55703_ (_04195_, _04194_, _04193_);
  not _55704_ (_04196_, _04195_);
  and _55705_ (_04197_, _04066_, _03191_);
  and _55706_ (_04198_, _03494_, _03191_);
  and _55707_ (_04199_, _04198_, _02994_);
  nor _55708_ (_04200_, _04199_, _04197_);
  and _55709_ (_04201_, _04200_, _04196_);
  and _55710_ (_04202_, _04201_, _04192_);
  not _55711_ (_04203_, _04202_);
  nor _55712_ (_04204_, _04203_, _04189_);
  and _55713_ (_04205_, _04204_, _04186_);
  nor _55714_ (_04206_, _04188_, _03787_);
  not _55715_ (_04207_, _03187_);
  nor _55716_ (_04208_, _03605_, _03221_);
  and _55717_ (_04209_, _04208_, _04122_);
  nor _55718_ (_04210_, _04209_, _04207_);
  and _55719_ (_04211_, _04058_, _03187_);
  nor _55720_ (_04212_, _04211_, _04003_);
  not _55721_ (_04213_, _04212_);
  nor _55722_ (_04214_, _04213_, _04210_);
  not _55723_ (_04215_, _04214_);
  nor _55724_ (_04216_, _04215_, _04206_);
  and _55725_ (_04217_, _04216_, _04205_);
  nor _55726_ (_04218_, _04048_, _03777_);
  or _55727_ (_04219_, _04218_, _04217_);
  and _55728_ (_04220_, _03798_, _03498_);
  nor _55729_ (_04221_, _04220_, _03621_);
  and _55730_ (_04222_, _04221_, _04219_);
  and _55731_ (_04223_, _03621_, _04051_);
  or _55732_ (_04224_, _04223_, _04222_);
  and _55733_ (_04225_, _03591_, _03202_);
  and _55734_ (_04226_, _04066_, _03202_);
  nor _55735_ (_04227_, _04226_, _04225_);
  not _55736_ (_04228_, _04227_);
  nor _55737_ (_04229_, _04124_, _03949_);
  nor _55738_ (_04230_, _04229_, _04228_);
  and _55739_ (_04231_, _04230_, _04224_);
  nor _55740_ (_04232_, _04048_, _03518_);
  or _55741_ (_04233_, _04232_, _04231_);
  and _55742_ (_04234_, _03515_, _03498_);
  nor _55743_ (_04235_, _04234_, _03628_);
  and _55744_ (_04236_, _04235_, _04233_);
  and _55745_ (_04237_, _03628_, _04051_);
  or _55746_ (_04238_, _04237_, _04236_);
  and _55747_ (_04239_, _02994_, _03197_);
  and _55748_ (_04240_, _04239_, _02962_);
  not _55749_ (_04241_, _04240_);
  and _55750_ (_04242_, _03605_, _03197_);
  nor _55751_ (_04243_, _04242_, _03815_);
  and _55752_ (_04244_, _04243_, _04241_);
  and _55753_ (_04245_, _04244_, _04238_);
  not _55754_ (_04246_, _03815_);
  nor _55755_ (_04247_, _04048_, _04246_);
  or _55756_ (_04248_, _04247_, _04245_);
  and _55757_ (_04249_, _04248_, _03823_);
  or _55758_ (_04250_, _04249_, _04052_);
  and _55759_ (_04251_, _03960_, _02994_);
  not _55760_ (_04252_, _04251_);
  and _55761_ (_04253_, _03493_, _03195_);
  and _55762_ (_04254_, _04253_, _02994_);
  not _55763_ (_04255_, _04254_);
  and _55764_ (_04256_, _03605_, _03195_);
  nor _55765_ (_04257_, _04256_, _03447_);
  and _55766_ (_04258_, _04257_, _04255_);
  and _55767_ (_04259_, _04258_, _04252_);
  nand _55768_ (_04260_, _04259_, _04250_);
  nand _55769_ (_04261_, _04260_, _04050_);
  or _55770_ (_04262_, _04261_, _04017_);
  nor _55771_ (_04263_, _03715_, _03505_);
  and _55772_ (_04264_, _03868_, _03586_);
  and _55773_ (_04265_, _04264_, _04263_);
  and _55774_ (_04266_, _04265_, _03867_);
  not _55775_ (_04267_, _04266_);
  and _55776_ (_04268_, _04267_, _03487_);
  not _55777_ (_04269_, _04268_);
  nor _55778_ (_04270_, _03414_, _03913_);
  not _55779_ (_04271_, _04270_);
  and _55780_ (_04272_, _03692_, _01949_);
  and _55781_ (_04273_, _03654_, _01917_);
  nor _55782_ (_04275_, _04273_, _04272_);
  and _55783_ (_04276_, _03672_, _01933_);
  and _55784_ (_04277_, _03680_, _01924_);
  nor _55785_ (_04278_, _04277_, _04276_);
  and _55786_ (_04279_, _04278_, _04275_);
  and _55787_ (_04280_, _03685_, _01946_);
  and _55788_ (_04281_, _03657_, _01944_);
  nor _55789_ (_04282_, _04281_, _04280_);
  and _55790_ (_04283_, _03687_, _01958_);
  and _55791_ (_04284_, _03665_, _01919_);
  nor _55792_ (_04285_, _04284_, _04283_);
  and _55793_ (_04286_, _04285_, _04282_);
  and _55794_ (_04287_, _04286_, _04279_);
  and _55795_ (_04288_, _03675_, _01930_);
  and _55796_ (_04289_, _03678_, _01956_);
  nor _55797_ (_04290_, _04289_, _04288_);
  and _55798_ (_04291_, _03696_, _01914_);
  and _55799_ (_04292_, _03703_, _01926_);
  nor _55800_ (_04293_, _04292_, _04291_);
  and _55801_ (_04294_, _04293_, _04290_);
  and _55802_ (_04295_, _03662_, _01941_);
  and _55803_ (_04296_, _03701_, _01909_);
  nor _55804_ (_04297_, _04296_, _04295_);
  and _55805_ (_04298_, _03690_, _01937_);
  and _55806_ (_04299_, _03698_, _01912_);
  nor _55807_ (_04300_, _04299_, _04298_);
  and _55808_ (_04301_, _04300_, _04297_);
  and _55809_ (_04302_, _04301_, _04294_);
  and _55810_ (_04303_, _04302_, _04287_);
  nor _55811_ (_04304_, _04303_, _03589_);
  and _55812_ (_04305_, _03493_, _03027_);
  and _55813_ (_04306_, _04305_, _03200_);
  and _55814_ (_04307_, _04305_, _03609_);
  nor _55815_ (_04308_, _04307_, _04306_);
  and _55816_ (_04309_, _04305_, _03168_);
  and _55817_ (_04310_, _04305_, _03202_);
  nor _55818_ (_04311_, _04310_, _04309_);
  and _55819_ (_04312_, _04311_, _04308_);
  and _55820_ (_04313_, _03954_, _03609_);
  nor _55821_ (_04314_, _03982_, _04313_);
  and _55822_ (_04315_, _04305_, _03191_);
  nor _55823_ (_04316_, _04315_, _03979_);
  and _55824_ (_04317_, _04316_, _04314_);
  and _55825_ (_04318_, _04317_, _04312_);
  and _55826_ (_04319_, _04318_, _03959_);
  and _55827_ (_04320_, _04305_, _03195_);
  not _55828_ (_04321_, _04320_);
  and _55829_ (_04322_, _04305_, _03197_);
  and _55830_ (_04323_, _03985_, _03027_);
  nor _55831_ (_04324_, _04323_, _04322_);
  and _55832_ (_04325_, _04324_, _04321_);
  and _55833_ (_04326_, _04305_, _03590_);
  nor _55834_ (_04327_, _03990_, _04326_);
  and _55835_ (_04328_, _04327_, _03973_);
  and _55836_ (_04329_, _03954_, _03195_);
  nor _55837_ (_04330_, _04329_, _03975_);
  and _55838_ (_04331_, _04330_, _04328_);
  and _55839_ (_04332_, _04331_, _04325_);
  not _55840_ (_04333_, _04305_);
  and _55841_ (_04334_, _03234_, _03247_);
  nor _55842_ (_04335_, _03181_, _03187_);
  and _55843_ (_04336_, _04335_, _03232_);
  and _55844_ (_04337_, _04336_, _04334_);
  nor _55845_ (_04338_, _04337_, _04333_);
  nor _55846_ (_04339_, _03998_, _03496_);
  nor _55847_ (_04340_, _04339_, _04338_);
  and _55848_ (_04341_, _04340_, _04332_);
  and _55849_ (_04342_, _04341_, _04319_);
  not _55850_ (_04343_, _04342_);
  nor _55851_ (_04344_, _04343_, _04304_);
  and _55852_ (_04345_, _04344_, _04271_);
  and _55853_ (_04346_, _04345_, _04269_);
  not _55854_ (_04347_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _55855_ (_04348_, _04260_, _04050_);
  or _55856_ (_04349_, _04348_, _04347_);
  and _55857_ (_04350_, _04349_, _04346_);
  nand _55858_ (_04351_, _04350_, _04262_);
  not _55859_ (_04352_, \oc8051_golden_model_1.IRAM[3] [1]);
  or _55860_ (_04353_, _04348_, _04352_);
  not _55861_ (_04354_, _04346_);
  not _55862_ (_04355_, \oc8051_golden_model_1.IRAM[2] [1]);
  or _55863_ (_04356_, _04261_, _04355_);
  and _55864_ (_04357_, _04356_, _04354_);
  nand _55865_ (_04358_, _04357_, _04353_);
  nand _55866_ (_04359_, _04358_, _04351_);
  nand _55867_ (_04360_, _04359_, _04016_);
  not _55868_ (_04361_, _04016_);
  not _55869_ (_04362_, \oc8051_golden_model_1.IRAM[7] [1]);
  or _55870_ (_04363_, _04348_, _04362_);
  not _55871_ (_04364_, \oc8051_golden_model_1.IRAM[6] [1]);
  or _55872_ (_04365_, _04261_, _04364_);
  and _55873_ (_04366_, _04365_, _04354_);
  nand _55874_ (_04367_, _04366_, _04363_);
  not _55875_ (_04368_, \oc8051_golden_model_1.IRAM[4] [1]);
  or _55876_ (_04369_, _04261_, _04368_);
  not _55877_ (_04370_, \oc8051_golden_model_1.IRAM[5] [1]);
  or _55878_ (_04371_, _04348_, _04370_);
  and _55879_ (_04372_, _04371_, _04346_);
  nand _55880_ (_04373_, _04372_, _04369_);
  nand _55881_ (_04374_, _04373_, _04367_);
  nand _55882_ (_04376_, _04374_, _04361_);
  nand _55883_ (_04377_, _04376_, _04360_);
  nand _55884_ (_04378_, _04377_, _03829_);
  not _55885_ (_04379_, _03829_);
  not _55886_ (_04380_, \oc8051_golden_model_1.IRAM[11] [1]);
  or _55887_ (_04381_, _04348_, _04380_);
  nand _55888_ (_04382_, _04348_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _55889_ (_04383_, _04382_, _04354_);
  nand _55890_ (_04384_, _04383_, _04381_);
  not _55891_ (_04385_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _55892_ (_04386_, _04261_, _04385_);
  nand _55893_ (_04387_, _04261_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _55894_ (_04388_, _04387_, _04346_);
  nand _55895_ (_04389_, _04388_, _04386_);
  nand _55896_ (_04390_, _04389_, _04384_);
  nand _55897_ (_04391_, _04390_, _04016_);
  not _55898_ (_04392_, \oc8051_golden_model_1.IRAM[15] [1]);
  or _55899_ (_04393_, _04348_, _04392_);
  nand _55900_ (_04394_, _04348_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _55901_ (_04395_, _04394_, _04354_);
  nand _55902_ (_04396_, _04395_, _04393_);
  not _55903_ (_04397_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _55904_ (_04398_, _04261_, _04397_);
  nand _55905_ (_04399_, _04261_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _55906_ (_04400_, _04399_, _04346_);
  nand _55907_ (_04401_, _04400_, _04398_);
  nand _55908_ (_04402_, _04401_, _04396_);
  nand _55909_ (_04403_, _04402_, _04361_);
  nand _55910_ (_04404_, _04403_, _04391_);
  nand _55911_ (_04405_, _04404_, _04379_);
  nand _55912_ (_04406_, _04405_, _04378_);
  and _55913_ (_04407_, _04406_, _03513_);
  or _55914_ (_04408_, _04407_, _03512_);
  and _55915_ (_04409_, _03612_, _03725_);
  and _55916_ (_04410_, _04409_, _03446_);
  and _55917_ (_04411_, _03414_, _04410_);
  or _55918_ (_04412_, _04411_, _04408_);
  and _55919_ (_04413_, _03500_, _03980_);
  not _55920_ (_04414_, _04413_);
  and _55921_ (_04415_, _03490_, _03609_);
  and _55922_ (_04416_, _03494_, _03609_);
  nor _55923_ (_04417_, _04416_, _04415_);
  and _55924_ (_04418_, _04417_, _04414_);
  not _55925_ (_04419_, _04418_);
  nor _55926_ (_04420_, _04419_, _04412_);
  and _55927_ (_04421_, _03610_, _03446_);
  nor _55928_ (_04422_, _03511_, _03229_);
  and _55929_ (_04423_, _04406_, _04422_);
  nor _55930_ (_04424_, _04423_, _04421_);
  and _55931_ (_04425_, _04424_, _04420_);
  and _55932_ (_04426_, _04421_, _03415_);
  nor _55933_ (_04427_, _04426_, _04425_);
  and _55934_ (_04428_, _03715_, _03446_);
  and _55935_ (_04429_, _03486_, _04428_);
  nor _55936_ (_04430_, _04429_, _04427_);
  and _55937_ (_04431_, _03723_, _03446_);
  nor _55938_ (_04432_, _03501_, _03230_);
  nor _55939_ (_04433_, _04432_, _04431_);
  and _55940_ (_04434_, _04433_, _04430_);
  and _55941_ (_04435_, _04431_, _03415_);
  nor _55942_ (_04436_, _04435_, _04434_);
  and _55943_ (_04437_, _03490_, _03507_);
  and _55944_ (_04438_, _03494_, _03507_);
  nor _55945_ (_04439_, _04438_, _04437_);
  not _55946_ (_04440_, _04439_);
  nor _55947_ (_04441_, _04440_, _04436_);
  and _55948_ (_04442_, _03729_, _03446_);
  nor _55949_ (_04443_, _03511_, _03232_);
  and _55950_ (_04444_, _04406_, _04443_);
  nor _55951_ (_04445_, _04444_, _04442_);
  and _55952_ (_04446_, _04445_, _04441_);
  and _55953_ (_04447_, _04442_, _03415_);
  nor _55954_ (_04448_, _04447_, _04446_);
  and _55955_ (_04449_, _03714_, _03446_);
  and _55956_ (_04450_, _03486_, _04449_);
  nor _55957_ (_04451_, _04450_, _04448_);
  and _55958_ (_04452_, _04451_, _03510_);
  nor _55959_ (_04453_, _04452_, _03509_);
  and _55960_ (_04454_, _03719_, _03446_);
  and _55961_ (_04455_, _04454_, _03486_);
  or _55962_ (_04456_, _04455_, _04453_);
  nor _55963_ (_04457_, _03501_, _03227_);
  and _55964_ (_04458_, _03745_, _03213_);
  nor _55965_ (_04459_, _04458_, _04457_);
  not _55966_ (_04460_, _04459_);
  nor _55967_ (_04461_, _04460_, _04456_);
  and _55968_ (_04462_, _03505_, _03446_);
  nor _55969_ (_04463_, _03511_, _03237_);
  and _55970_ (_04464_, _04406_, _04463_);
  nor _55971_ (_04465_, _04464_, _04462_);
  and _55972_ (_04466_, _04465_, _04461_);
  nor _55973_ (_04467_, _04466_, _03506_);
  nor _55974_ (_04468_, _04467_, _03224_);
  and _55975_ (_04469_, _03501_, _03224_);
  nor _55976_ (_04470_, _04469_, _04468_);
  and _55977_ (_04471_, _03446_, _03168_);
  and _55978_ (_04472_, _04471_, _03494_);
  not _55979_ (_04473_, _04309_);
  or _55980_ (_04474_, _03592_, _03954_);
  and _55981_ (_04475_, _04474_, _03168_);
  nor _55982_ (_04477_, _04475_, _03969_);
  and _55983_ (_04478_, _04477_, _04473_);
  nor _55984_ (_04479_, _04478_, _03454_);
  nor _55985_ (_04480_, _04479_, _04472_);
  nor _55986_ (_04481_, _03511_, _03212_);
  and _55987_ (_04482_, _04481_, _03446_);
  and _55988_ (_04483_, _04471_, _03221_);
  nor _55989_ (_04484_, _04483_, _04482_);
  and _55990_ (_04485_, _04484_, _04480_);
  nor _55991_ (_04486_, _04485_, _03415_);
  and _55992_ (_04487_, _03592_, _03176_);
  and _55993_ (_04488_, _03493_, _03218_);
  and _55994_ (_04489_, _04488_, _03176_);
  or _55995_ (_04490_, _04489_, _04487_);
  not _55996_ (_04491_, _04490_);
  and _55997_ (_04492_, _04058_, _03176_);
  and _55998_ (_04493_, _03595_, _03176_);
  nor _55999_ (_04494_, _04493_, _04492_);
  and _56000_ (_04495_, _04494_, _04491_);
  not _56001_ (_04496_, _04495_);
  nor _56002_ (_04497_, _04496_, _04486_);
  not _56003_ (_04498_, _04497_);
  nor _56004_ (_04499_, _04498_, _04470_);
  and _56005_ (_04500_, _03601_, _03446_);
  not _56006_ (_04501_, _03176_);
  nor _56007_ (_04502_, _03511_, _04501_);
  and _56008_ (_04503_, _04406_, _04502_);
  nor _56009_ (_04504_, _04503_, _04500_);
  and _56010_ (_04505_, _04504_, _04499_);
  and _56011_ (_04506_, _04500_, _03415_);
  nor _56012_ (_04507_, _04506_, _04505_);
  nor _56013_ (_04508_, _04507_, _03178_);
  and _56014_ (_04509_, _03501_, _03178_);
  nor _56015_ (_04510_, _04509_, _04508_);
  and _56016_ (_04511_, _03780_, _03446_);
  and _56017_ (_04512_, _03600_, _03446_);
  nor _56018_ (_04513_, _04512_, _04511_);
  and _56019_ (_04514_, _03790_, _03446_);
  and _56020_ (_04515_, _03622_, _03446_);
  nor _56021_ (_04516_, _04515_, _04514_);
  and _56022_ (_04517_, _04516_, _04513_);
  nor _56023_ (_04518_, _04517_, _03415_);
  nor _56024_ (_04519_, _04518_, _03192_);
  not _56025_ (_04520_, _04519_);
  nor _56026_ (_04521_, _04520_, _04510_);
  and _56027_ (_04522_, _03501_, _03192_);
  nor _56028_ (_04523_, _04522_, _04521_);
  nor _56029_ (_04524_, _03786_, _03454_);
  and _56030_ (_04525_, _04524_, _03414_);
  or _56031_ (_04526_, _04525_, _03188_);
  nor _56032_ (_04527_, _04526_, _04523_);
  nor _56033_ (_04528_, _04527_, _03502_);
  nor _56034_ (_04529_, _04528_, _03495_);
  and _56035_ (_04530_, _04529_, _03492_);
  and _56036_ (_04531_, _03815_, _03446_);
  not _56037_ (_04532_, _03197_);
  nor _56038_ (_04533_, _03511_, _04532_);
  and _56039_ (_04534_, _04406_, _04533_);
  nor _56040_ (_04535_, _04534_, _04531_);
  and _56041_ (_04536_, _04535_, _04530_);
  and _56042_ (_04537_, _04531_, _03415_);
  nor _56043_ (_04538_, _04537_, _04536_);
  and _56044_ (_04539_, _03446_, _03453_);
  nor _56045_ (_04540_, _03629_, _03198_);
  nor _56046_ (_04541_, _03501_, _04540_);
  nor _56047_ (_04542_, _04541_, _04539_);
  not _56048_ (_04543_, _04542_);
  nor _56049_ (_04544_, _04543_, _04538_);
  nor _56050_ (_04545_, _04544_, _03488_);
  and _56051_ (_04546_, _03490_, _03195_);
  and _56052_ (_04547_, _03494_, _03195_);
  nor _56053_ (_04548_, _04547_, _04546_);
  not _56054_ (_04549_, _04548_);
  nor _56055_ (_04550_, _04549_, _04545_);
  not _56056_ (_04551_, _03195_);
  nor _56057_ (_04552_, _03511_, _04551_);
  and _56058_ (_04553_, _04406_, _04552_);
  nor _56059_ (_04554_, _04553_, _03448_);
  and _56060_ (_04555_, _04554_, _04550_);
  nor _56061_ (_04556_, _04555_, _03449_);
  not _56062_ (_04557_, _04556_);
  not _56063_ (_04558_, _04539_);
  and _56064_ (_04559_, _03188_, _03498_);
  nor _56065_ (_04560_, _04485_, _04188_);
  and _56066_ (_04561_, _03719_, _04051_);
  not _56067_ (_04562_, _04454_);
  not _56068_ (_04563_, \oc8051_golden_model_1.IRAM[0] [0]);
  or _56069_ (_04564_, _04261_, _04563_);
  not _56070_ (_04565_, \oc8051_golden_model_1.IRAM[1] [0]);
  or _56071_ (_04566_, _04348_, _04565_);
  and _56072_ (_04567_, _04566_, _04346_);
  nand _56073_ (_04568_, _04567_, _04564_);
  not _56074_ (_04569_, \oc8051_golden_model_1.IRAM[3] [0]);
  or _56075_ (_04570_, _04348_, _04569_);
  not _56076_ (_04571_, \oc8051_golden_model_1.IRAM[2] [0]);
  or _56077_ (_04572_, _04261_, _04571_);
  and _56078_ (_04573_, _04572_, _04354_);
  nand _56079_ (_04574_, _04573_, _04570_);
  nand _56080_ (_04575_, _04574_, _04568_);
  nand _56081_ (_04576_, _04575_, _04016_);
  not _56082_ (_04578_, \oc8051_golden_model_1.IRAM[7] [0]);
  or _56083_ (_04579_, _04348_, _04578_);
  not _56084_ (_04580_, \oc8051_golden_model_1.IRAM[6] [0]);
  or _56085_ (_04581_, _04261_, _04580_);
  and _56086_ (_04582_, _04581_, _04354_);
  nand _56087_ (_04583_, _04582_, _04579_);
  not _56088_ (_04584_, \oc8051_golden_model_1.IRAM[4] [0]);
  or _56089_ (_04585_, _04261_, _04584_);
  not _56090_ (_04586_, \oc8051_golden_model_1.IRAM[5] [0]);
  or _56091_ (_04587_, _04348_, _04586_);
  and _56092_ (_04588_, _04587_, _04346_);
  nand _56093_ (_04589_, _04588_, _04585_);
  nand _56094_ (_04590_, _04589_, _04583_);
  nand _56095_ (_04591_, _04590_, _04361_);
  nand _56096_ (_04592_, _04591_, _04576_);
  nand _56097_ (_04593_, _04592_, _03829_);
  not _56098_ (_04594_, \oc8051_golden_model_1.IRAM[11] [0]);
  or _56099_ (_04595_, _04348_, _04594_);
  nand _56100_ (_04596_, _04348_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _56101_ (_04597_, _04596_, _04354_);
  nand _56102_ (_04598_, _04597_, _04595_);
  not _56103_ (_04599_, \oc8051_golden_model_1.IRAM[8] [0]);
  or _56104_ (_04600_, _04261_, _04599_);
  nand _56105_ (_04601_, _04261_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _56106_ (_04602_, _04601_, _04346_);
  nand _56107_ (_04603_, _04602_, _04600_);
  nand _56108_ (_04604_, _04603_, _04598_);
  nand _56109_ (_04605_, _04604_, _04016_);
  not _56110_ (_04606_, \oc8051_golden_model_1.IRAM[15] [0]);
  or _56111_ (_04607_, _04348_, _04606_);
  nand _56112_ (_04608_, _04348_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _56113_ (_04609_, _04608_, _04354_);
  nand _56114_ (_04610_, _04609_, _04607_);
  not _56115_ (_04611_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _56116_ (_04612_, _04261_, _04611_);
  nand _56117_ (_04613_, _04261_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _56118_ (_04614_, _04613_, _04346_);
  nand _56119_ (_04615_, _04614_, _04612_);
  nand _56120_ (_04616_, _04615_, _04610_);
  nand _56121_ (_04617_, _04616_, _04361_);
  nand _56122_ (_04618_, _04617_, _04605_);
  nand _56123_ (_04619_, _04618_, _04379_);
  and _56124_ (_04620_, _04619_, _04593_);
  and _56125_ (_04621_, _04620_, _03513_);
  nor _56126_ (_04622_, _03603_, _03030_);
  and _56127_ (_04623_, _04622_, _04059_);
  nor _56128_ (_04624_, _04623_, _03239_);
  not _56129_ (_04625_, _04624_);
  nor _56130_ (_04626_, _04625_, _04621_);
  and _56131_ (_04627_, _04048_, _04410_);
  or _56132_ (_04628_, _04627_, _04626_);
  and _56133_ (_04629_, _03980_, \oc8051_golden_model_1.SP [0]);
  and _56134_ (_04630_, _04100_, _03609_);
  nor _56135_ (_04631_, _04630_, _04629_);
  not _56136_ (_04632_, _04631_);
  nor _56137_ (_04633_, _04632_, _04628_);
  nand _56138_ (_04634_, _04619_, _04593_);
  and _56139_ (_04635_, _04422_, _04634_);
  nor _56140_ (_04636_, _04635_, _04421_);
  and _56141_ (_04637_, _04636_, _04633_);
  and _56142_ (_04638_, _04421_, _04188_);
  nor _56143_ (_04639_, _04638_, _04637_);
  nor _56144_ (_04640_, _04639_, _04428_);
  not _56145_ (_04641_, _04640_);
  and _56146_ (_04642_, _04641_, _04085_);
  nor _56147_ (_04643_, _03230_, _03498_);
  nor _56148_ (_04644_, _04643_, _04642_);
  and _56149_ (_04645_, _04431_, _04048_);
  and _56150_ (_04646_, _04100_, _03507_);
  nor _56151_ (_04647_, _04646_, _04645_);
  and _56152_ (_04648_, _04647_, _04644_);
  and _56153_ (_04649_, _04443_, _04634_);
  not _56154_ (_04650_, _04649_);
  and _56155_ (_04651_, _04650_, _04648_);
  and _56156_ (_04652_, _04442_, _04048_);
  nor _56157_ (_04653_, _04652_, _04449_);
  and _56158_ (_04654_, _04653_, _04651_);
  nor _56159_ (_04655_, _04654_, _04096_);
  nor _56160_ (_04656_, _04655_, _03508_);
  and _56161_ (_04657_, _03508_, _03498_);
  or _56162_ (_04658_, _04657_, _04656_);
  and _56163_ (_04659_, _04658_, _04562_);
  nor _56164_ (_04660_, _04659_, _04561_);
  nor _56165_ (_04661_, _03227_, _03498_);
  and _56166_ (_04662_, _04100_, _03751_);
  nor _56167_ (_04663_, _04662_, _04661_);
  not _56168_ (_04664_, _04663_);
  nor _56169_ (_04665_, _04664_, _04660_);
  and _56170_ (_04666_, _04463_, _04634_);
  nor _56171_ (_04667_, _04666_, _04462_);
  and _56172_ (_04668_, _04667_, _04665_);
  nor _56173_ (_04669_, _04668_, _04053_);
  nor _56174_ (_04670_, _04669_, _03224_);
  and _56175_ (_04671_, _03224_, _03498_);
  nor _56176_ (_04672_, _04671_, _04670_);
  and _56177_ (_04673_, _04100_, _03176_);
  or _56178_ (_04674_, _04673_, _04672_);
  nor _56179_ (_04675_, _04674_, _04560_);
  and _56180_ (_04676_, _04502_, _04634_);
  not _56181_ (_04677_, _04676_);
  and _56182_ (_04679_, _04677_, _04675_);
  and _56183_ (_04680_, _04500_, _04048_);
  nor _56184_ (_04681_, _04680_, _03178_);
  and _56185_ (_04682_, _04681_, _04679_);
  and _56186_ (_04683_, _03178_, _03498_);
  nor _56187_ (_04684_, _04683_, _04682_);
  nor _56188_ (_04685_, _04517_, _04188_);
  nor _56189_ (_04686_, _04685_, _03192_);
  not _56190_ (_04687_, _04686_);
  nor _56191_ (_04688_, _04687_, _04684_);
  and _56192_ (_04689_, _03192_, _03498_);
  nor _56193_ (_04690_, _04689_, _04688_);
  and _56194_ (_04691_, _04524_, _04048_);
  or _56195_ (_04692_, _04691_, _03188_);
  nor _56196_ (_04693_, _04692_, _04690_);
  nor _56197_ (_04694_, _04693_, _04559_);
  nor _56198_ (_04695_, _04694_, _04240_);
  and _56199_ (_04696_, _04533_, _04634_);
  nor _56200_ (_04697_, _04696_, _04531_);
  and _56201_ (_04698_, _04697_, _04695_);
  and _56202_ (_04699_, _04531_, _04188_);
  nor _56203_ (_04700_, _04699_, _04698_);
  nor _56204_ (_04701_, _04540_, _03498_);
  nor _56205_ (_04702_, _04701_, _04700_);
  and _56206_ (_04703_, _04702_, _04558_);
  nor _56207_ (_04704_, _04703_, _04052_);
  and _56208_ (_04705_, _04100_, _03195_);
  nor _56209_ (_04706_, _04705_, _04704_);
  and _56210_ (_04707_, _04552_, _04634_);
  nor _56211_ (_04708_, _04707_, _03448_);
  and _56212_ (_04709_, _04708_, _04706_);
  and _56213_ (_04710_, _03448_, _04188_);
  nor _56214_ (_04711_, _04710_, _04709_);
  nor _56215_ (_04712_, _04483_, _04472_);
  not _56216_ (_04713_, _03448_);
  and _56217_ (_04714_, _03593_, _03176_);
  not _56218_ (_04715_, _04714_);
  and _56219_ (_04716_, _03493_, _03176_);
  and _56220_ (_04717_, _04716_, _03027_);
  nor _56221_ (_04718_, _04717_, _04546_);
  and _56222_ (_04719_, _04718_, _04715_);
  and _56223_ (_04720_, _04719_, _04325_);
  or _56224_ (_04721_, _03593_, _03595_);
  and _56225_ (_04722_, _04721_, _03751_);
  not _56226_ (_04723_, _03221_);
  and _56227_ (_04724_, _04622_, _04723_);
  nor _56228_ (_04725_, _04724_, _03239_);
  not _56229_ (_04726_, _03494_);
  and _56230_ (_04727_, _03511_, _04726_);
  nor _56231_ (_04728_, _04727_, _03239_);
  or _56232_ (_04729_, _04728_, _04725_);
  nor _56233_ (_04730_, _04729_, _04722_);
  and _56234_ (_04731_, _04730_, _04720_);
  and _56235_ (_04732_, _04716_, _03218_);
  nor _56236_ (_04733_, _04732_, _04493_);
  nor _56237_ (_04734_, _04502_, _04492_);
  and _56238_ (_04735_, _04540_, _03193_);
  and _56239_ (_04736_, _04735_, _04734_);
  and _56240_ (_04737_, _04736_, _04733_);
  nor _56241_ (_04738_, _04463_, _04443_);
  nor _56242_ (_04739_, _04552_, _04422_);
  and _56243_ (_04740_, _04739_, _04738_);
  nor _56244_ (_04741_, _03491_, _03972_);
  nor _56245_ (_04742_, _04307_, _03962_);
  and _56246_ (_04743_, _04742_, _04741_);
  and _56247_ (_04744_, _04743_, _04740_);
  not _56248_ (_04745_, _03495_);
  and _56249_ (_04746_, _03612_, _03751_);
  nor _56250_ (_04747_, _04416_, _04746_);
  and _56251_ (_04748_, _04747_, _04745_);
  and _56252_ (_04749_, _04305_, _03751_);
  or _56253_ (_04750_, _04488_, _04305_);
  and _56254_ (_04751_, _04750_, _03507_);
  nor _56255_ (_04752_, _04751_, _04749_);
  and _56256_ (_04753_, _03494_, _03751_);
  and _56257_ (_04754_, _03612_, _03176_);
  nor _56258_ (_04755_, _04754_, _04753_);
  and _56259_ (_04756_, _04755_, _04752_);
  and _56260_ (_04757_, _04756_, _04748_);
  and _56261_ (_04758_, _04757_, _04744_);
  and _56262_ (_04759_, _04058_, _03507_);
  nor _56263_ (_04760_, _04329_, _04759_);
  nor _56264_ (_04761_, _04547_, _04437_);
  and _56265_ (_04762_, _04761_, _04760_);
  not _56266_ (_04763_, _03980_);
  nor _56267_ (_04764_, _04533_, _03508_);
  and _56268_ (_04765_, _04764_, _04763_);
  not _56269_ (_04766_, _03227_);
  nor _56270_ (_04767_, _04766_, _03224_);
  not _56271_ (_04768_, _03230_);
  nor _56272_ (_04769_, _04768_, _03178_);
  and _56273_ (_04770_, _04769_, _04767_);
  and _56274_ (_04771_, _04770_, _04765_);
  and _56275_ (_04772_, _04771_, _04762_);
  and _56276_ (_04773_, _04772_, _04758_);
  and _56277_ (_04774_, _04773_, _04737_);
  and _56278_ (_04775_, _04774_, _04731_);
  and _56279_ (_04776_, _04775_, _04713_);
  nor _56280_ (_04777_, _04500_, _04442_);
  and _56281_ (_04778_, _04777_, _04776_);
  and _56282_ (_04780_, _04778_, _04712_);
  nor _56283_ (_04781_, _04482_, _04479_);
  nor _56284_ (_04782_, _03714_, _03453_);
  and _56285_ (_04783_, _04782_, _04246_);
  and _56286_ (_04784_, _04783_, _04263_);
  nor _56287_ (_04785_, _04784_, _03454_);
  nor _56288_ (_04786_, _04785_, _04524_);
  and _56289_ (_04787_, _04786_, _04781_);
  nor _56290_ (_04788_, _04431_, _04410_);
  nor _56291_ (_04789_, _04454_, _04421_);
  and _56292_ (_04790_, _04789_, _04788_);
  and _56293_ (_04791_, _04790_, _04787_);
  and _56294_ (_04792_, _04791_, _04517_);
  and _56295_ (_04793_, _04792_, _04780_);
  and _56296_ (_04794_, _43868_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not _56297_ (_04795_, _04794_);
  nor _56298_ (_04796_, _04795_, _04793_);
  not _56299_ (_04797_, _04796_);
  nor _56300_ (_04798_, _04797_, _04711_);
  and _56301_ (_04799_, _04798_, _04557_);
  not _56302_ (_04800_, _03904_);
  and _56303_ (_04801_, _03448_, _04800_);
  and _56304_ (_04802_, _03861_, _03453_);
  and _56305_ (_04803_, _03493_, _03197_);
  and _56306_ (_04804_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _56307_ (_04805_, _04804_, \oc8051_golden_model_1.SP [2]);
  nor _56308_ (_04806_, _04804_, \oc8051_golden_model_1.SP [2]);
  nor _56309_ (_04807_, _04806_, _04805_);
  and _56310_ (_04808_, _04807_, _03188_);
  and _56311_ (_04809_, _04500_, _04800_);
  and _56312_ (_04810_, _03861_, _03505_);
  and _56313_ (_04811_, _04807_, _03508_);
  and _56314_ (_04812_, _04421_, _04800_);
  not _56315_ (_04813_, _04807_);
  and _56316_ (_04814_, _04813_, _03980_);
  and _56317_ (_04815_, _03493_, _03609_);
  nor _56318_ (_04816_, _04815_, _04814_);
  and _56319_ (_04817_, _03904_, _04410_);
  not _56320_ (_04818_, _04725_);
  not _56321_ (_04819_, \oc8051_golden_model_1.IRAM[0] [2]);
  or _56322_ (_04820_, _04261_, _04819_);
  not _56323_ (_04821_, \oc8051_golden_model_1.IRAM[1] [2]);
  or _56324_ (_04822_, _04348_, _04821_);
  and _56325_ (_04823_, _04822_, _04346_);
  nand _56326_ (_04824_, _04823_, _04820_);
  not _56327_ (_04825_, \oc8051_golden_model_1.IRAM[3] [2]);
  or _56328_ (_04826_, _04348_, _04825_);
  not _56329_ (_04827_, \oc8051_golden_model_1.IRAM[2] [2]);
  or _56330_ (_04828_, _04261_, _04827_);
  and _56331_ (_04829_, _04828_, _04354_);
  nand _56332_ (_04830_, _04829_, _04826_);
  nand _56333_ (_04831_, _04830_, _04824_);
  nand _56334_ (_04832_, _04831_, _04016_);
  not _56335_ (_04833_, \oc8051_golden_model_1.IRAM[7] [2]);
  or _56336_ (_04834_, _04348_, _04833_);
  not _56337_ (_04835_, \oc8051_golden_model_1.IRAM[6] [2]);
  or _56338_ (_04836_, _04261_, _04835_);
  and _56339_ (_04837_, _04836_, _04354_);
  nand _56340_ (_04838_, _04837_, _04834_);
  not _56341_ (_04839_, \oc8051_golden_model_1.IRAM[4] [2]);
  or _56342_ (_04840_, _04261_, _04839_);
  not _56343_ (_04841_, \oc8051_golden_model_1.IRAM[5] [2]);
  or _56344_ (_04842_, _04348_, _04841_);
  and _56345_ (_04843_, _04842_, _04346_);
  nand _56346_ (_04844_, _04843_, _04840_);
  nand _56347_ (_04845_, _04844_, _04838_);
  nand _56348_ (_04846_, _04845_, _04361_);
  nand _56349_ (_04847_, _04846_, _04832_);
  nand _56350_ (_04848_, _04847_, _03829_);
  not _56351_ (_04849_, \oc8051_golden_model_1.IRAM[11] [2]);
  or _56352_ (_04850_, _04348_, _04849_);
  not _56353_ (_04851_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _56354_ (_04852_, _04261_, _04851_);
  and _56355_ (_04853_, _04852_, _04354_);
  nand _56356_ (_04854_, _04853_, _04850_);
  nand _56357_ (_04855_, _04348_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand _56358_ (_04856_, _04261_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _56359_ (_04857_, _04856_, _04346_);
  nand _56360_ (_04858_, _04857_, _04855_);
  nand _56361_ (_04859_, _04858_, _04854_);
  nand _56362_ (_04860_, _04859_, _04016_);
  not _56363_ (_04861_, \oc8051_golden_model_1.IRAM[15] [2]);
  or _56364_ (_04862_, _04348_, _04861_);
  not _56365_ (_04863_, \oc8051_golden_model_1.IRAM[14] [2]);
  or _56366_ (_04864_, _04261_, _04863_);
  and _56367_ (_04865_, _04864_, _04354_);
  nand _56368_ (_04866_, _04865_, _04862_);
  nand _56369_ (_04867_, _04348_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand _56370_ (_04868_, _04261_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _56371_ (_04869_, _04868_, _04346_);
  nand _56372_ (_04870_, _04869_, _04867_);
  nand _56373_ (_04871_, _04870_, _04866_);
  nand _56374_ (_04872_, _04871_, _04361_);
  nand _56375_ (_04873_, _04872_, _04860_);
  nand _56376_ (_04874_, _04873_, _04379_);
  nand _56377_ (_04875_, _04874_, _04848_);
  nor _56378_ (_04876_, _04875_, _03029_);
  nor _56379_ (_04877_, _04876_, _04818_);
  nor _56380_ (_04878_, _04877_, _04817_);
  and _56381_ (_04879_, _04878_, _04816_);
  and _56382_ (_04880_, _04875_, _04422_);
  nor _56383_ (_04881_, _04880_, _04421_);
  and _56384_ (_04882_, _04881_, _04879_);
  nor _56385_ (_04883_, _04882_, _04812_);
  nor _56386_ (_04884_, _04883_, _04428_);
  nor _56387_ (_04885_, _04884_, _03862_);
  nor _56388_ (_04886_, _04807_, _03230_);
  nor _56389_ (_04887_, _04886_, _04885_);
  and _56390_ (_04888_, _03493_, _03507_);
  and _56391_ (_04889_, _04431_, _03904_);
  nor _56392_ (_04890_, _04889_, _04888_);
  and _56393_ (_04891_, _04890_, _04887_);
  and _56394_ (_04892_, _04875_, _04443_);
  nor _56395_ (_04893_, _04892_, _04442_);
  and _56396_ (_04894_, _04893_, _04891_);
  and _56397_ (_04895_, _04442_, _04800_);
  nor _56398_ (_04896_, _04895_, _04894_);
  and _56399_ (_04897_, _03860_, _04449_);
  nor _56400_ (_04898_, _04897_, _04896_);
  and _56401_ (_04899_, _04898_, _03510_);
  nor _56402_ (_04900_, _04899_, _04811_);
  and _56403_ (_04901_, _04454_, _03860_);
  or _56404_ (_04902_, _04901_, _04900_);
  and _56405_ (_04903_, _03493_, _03751_);
  nor _56406_ (_04904_, _04807_, _03227_);
  nor _56407_ (_04905_, _04904_, _04903_);
  not _56408_ (_04906_, _04905_);
  nor _56409_ (_04907_, _04906_, _04902_);
  and _56410_ (_04908_, _04875_, _04463_);
  nor _56411_ (_04909_, _04908_, _04462_);
  and _56412_ (_04910_, _04909_, _04907_);
  nor _56413_ (_04911_, _04910_, _04810_);
  nor _56414_ (_04912_, _04911_, _03224_);
  and _56415_ (_04913_, _04807_, _03224_);
  nor _56416_ (_04914_, _04913_, _04912_);
  nor _56417_ (_04915_, _04485_, _04800_);
  nor _56418_ (_04916_, _04915_, _04716_);
  not _56419_ (_04917_, _04916_);
  nor _56420_ (_04918_, _04917_, _04914_);
  and _56421_ (_04919_, _04875_, _04502_);
  nor _56422_ (_04920_, _04919_, _04500_);
  and _56423_ (_04921_, _04920_, _04918_);
  nor _56424_ (_04922_, _04921_, _04809_);
  nor _56425_ (_04923_, _04922_, _03178_);
  and _56426_ (_04924_, _04807_, _03178_);
  nor _56427_ (_04925_, _04924_, _04923_);
  nor _56428_ (_04926_, _04517_, _04800_);
  nor _56429_ (_04927_, _04926_, _03192_);
  not _56430_ (_04928_, _04927_);
  nor _56431_ (_04929_, _04928_, _04925_);
  and _56432_ (_04930_, _04807_, _03192_);
  nor _56433_ (_04931_, _04930_, _04929_);
  and _56434_ (_04932_, _04524_, _03904_);
  or _56435_ (_04933_, _04932_, _03188_);
  nor _56436_ (_04934_, _04933_, _04931_);
  nor _56437_ (_04935_, _04934_, _04808_);
  nor _56438_ (_04936_, _04935_, _04803_);
  and _56439_ (_04937_, _04875_, _04533_);
  nor _56440_ (_04938_, _04937_, _04531_);
  and _56441_ (_04939_, _04938_, _04936_);
  and _56442_ (_04940_, _04531_, _04800_);
  nor _56443_ (_04941_, _04940_, _04939_);
  nor _56444_ (_04942_, _04807_, _04540_);
  nor _56445_ (_04943_, _04942_, _04539_);
  not _56446_ (_04944_, _04943_);
  nor _56447_ (_04945_, _04944_, _04941_);
  nor _56448_ (_04946_, _04945_, _04802_);
  nor _56449_ (_04947_, _04946_, _04253_);
  and _56450_ (_04948_, _04875_, _04552_);
  nor _56451_ (_04949_, _04948_, _03448_);
  and _56452_ (_04950_, _04949_, _04947_);
  nor _56453_ (_04951_, _04950_, _04801_);
  not _56454_ (_04952_, _04951_);
  not _56455_ (_04953_, \oc8051_golden_model_1.IRAM[0] [3]);
  or _56456_ (_04954_, _04261_, _04953_);
  not _56457_ (_04955_, \oc8051_golden_model_1.IRAM[1] [3]);
  or _56458_ (_04956_, _04348_, _04955_);
  and _56459_ (_04957_, _04956_, _04346_);
  nand _56460_ (_04958_, _04957_, _04954_);
  not _56461_ (_04959_, \oc8051_golden_model_1.IRAM[3] [3]);
  or _56462_ (_04960_, _04348_, _04959_);
  not _56463_ (_04961_, \oc8051_golden_model_1.IRAM[2] [3]);
  or _56464_ (_04962_, _04261_, _04961_);
  and _56465_ (_04963_, _04962_, _04354_);
  nand _56466_ (_04964_, _04963_, _04960_);
  nand _56467_ (_04965_, _04964_, _04958_);
  nand _56468_ (_04966_, _04965_, _04016_);
  not _56469_ (_04967_, \oc8051_golden_model_1.IRAM[7] [3]);
  or _56470_ (_04968_, _04348_, _04967_);
  not _56471_ (_04969_, \oc8051_golden_model_1.IRAM[6] [3]);
  or _56472_ (_04970_, _04261_, _04969_);
  and _56473_ (_04971_, _04970_, _04354_);
  nand _56474_ (_04972_, _04971_, _04968_);
  not _56475_ (_04973_, \oc8051_golden_model_1.IRAM[4] [3]);
  or _56476_ (_04974_, _04261_, _04973_);
  not _56477_ (_04975_, \oc8051_golden_model_1.IRAM[5] [3]);
  or _56478_ (_04976_, _04348_, _04975_);
  and _56479_ (_04977_, _04976_, _04346_);
  nand _56480_ (_04978_, _04977_, _04974_);
  nand _56481_ (_04979_, _04978_, _04972_);
  nand _56482_ (_04980_, _04979_, _04361_);
  nand _56483_ (_04981_, _04980_, _04966_);
  nand _56484_ (_04982_, _04981_, _03829_);
  nand _56485_ (_04983_, _04261_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _56486_ (_04984_, _04348_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _56487_ (_04985_, _04984_, _04354_);
  nand _56488_ (_04986_, _04985_, _04983_);
  nand _56489_ (_04987_, _04348_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand _56490_ (_04988_, _04261_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _56491_ (_04989_, _04988_, _04346_);
  nand _56492_ (_04990_, _04989_, _04987_);
  nand _56493_ (_04991_, _04990_, _04986_);
  nand _56494_ (_04992_, _04991_, _04016_);
  nand _56495_ (_04993_, _04261_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _56496_ (_04994_, _04348_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _56497_ (_04995_, _04994_, _04354_);
  nand _56498_ (_04996_, _04995_, _04993_);
  nand _56499_ (_04997_, _04348_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand _56500_ (_04998_, _04261_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _56501_ (_04999_, _04998_, _04346_);
  nand _56502_ (_05000_, _04999_, _04997_);
  nand _56503_ (_05001_, _05000_, _04996_);
  nand _56504_ (_05002_, _05001_, _04361_);
  nand _56505_ (_05003_, _05002_, _04992_);
  nand _56506_ (_05004_, _05003_, _04379_);
  nand _56507_ (_05005_, _05004_, _04982_);
  and _56508_ (_05006_, _05005_, _04502_);
  and _56509_ (_05007_, _05005_, _04463_);
  nor _56510_ (_05008_, _04805_, \oc8051_golden_model_1.SP [3]);
  and _56511_ (_05009_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _56512_ (_05010_, _05009_, \oc8051_golden_model_1.SP [3]);
  and _56513_ (_05011_, _05010_, \oc8051_golden_model_1.SP [0]);
  nor _56514_ (_05012_, _05011_, _05008_);
  and _56515_ (_05013_, _05012_, _04766_);
  and _56516_ (_05014_, _03549_, _04428_);
  and _56517_ (_05015_, _05005_, _04422_);
  and _56518_ (_05016_, _05012_, _03980_);
  and _56519_ (_05017_, _05005_, _03513_);
  not _56520_ (_05018_, \oc8051_golden_model_1.PSW [3]);
  and _56521_ (_05019_, _03240_, _05018_);
  nor _56522_ (_05020_, _05019_, _04410_);
  not _56523_ (_05021_, _05020_);
  nor _56524_ (_05022_, _05021_, _05017_);
  and _56525_ (_05023_, _04409_, _04051_);
  nor _56526_ (_05024_, _05023_, _05022_);
  nor _56527_ (_05025_, _05024_, _03980_);
  or _56528_ (_05026_, _05025_, _04422_);
  nor _56529_ (_05027_, _05026_, _05016_);
  or _56530_ (_05028_, _05027_, _04421_);
  nor _56531_ (_05029_, _05028_, _05015_);
  and _56532_ (_05030_, _04421_, _03756_);
  or _56533_ (_05031_, _05030_, _04428_);
  nor _56534_ (_05032_, _05031_, _05029_);
  nor _56535_ (_05033_, _05032_, _05014_);
  nor _56536_ (_05034_, _05033_, _04768_);
  nor _56537_ (_05035_, _05012_, _03230_);
  nor _56538_ (_05036_, _05035_, _04431_);
  not _56539_ (_05037_, _05036_);
  nor _56540_ (_05038_, _05037_, _05034_);
  and _56541_ (_05039_, _04431_, _03756_);
  nor _56542_ (_05040_, _05039_, _04443_);
  not _56543_ (_05041_, _05040_);
  nor _56544_ (_05042_, _05041_, _05038_);
  and _56545_ (_05043_, _05005_, _04443_);
  nor _56546_ (_05044_, _05043_, _04442_);
  not _56547_ (_05045_, _05044_);
  nor _56548_ (_05046_, _05045_, _05042_);
  and _56549_ (_05047_, _04442_, _03756_);
  or _56550_ (_05048_, _05047_, _04449_);
  nor _56551_ (_05049_, _05048_, _05046_);
  and _56552_ (_05050_, _03549_, _04449_);
  nor _56553_ (_05051_, _05050_, _05049_);
  and _56554_ (_05052_, _05051_, _03510_);
  and _56555_ (_05053_, _05012_, _03508_);
  nor _56556_ (_05054_, _05053_, _05052_);
  nor _56557_ (_05055_, _05054_, _04454_);
  nor _56558_ (_05056_, _04562_, _03583_);
  or _56559_ (_05057_, _05056_, _05055_);
  and _56560_ (_05058_, _05057_, _03227_);
  or _56561_ (_05059_, _05058_, _04463_);
  nor _56562_ (_05060_, _05059_, _05013_);
  or _56563_ (_05061_, _05060_, _04462_);
  nor _56564_ (_05062_, _05061_, _05007_);
  not _56565_ (_05063_, _04462_);
  nor _56566_ (_05064_, _05063_, _03583_);
  nor _56567_ (_05065_, _05064_, _05062_);
  nor _56568_ (_05066_, _05065_, _03224_);
  and _56569_ (_05067_, _05012_, _03224_);
  not _56570_ (_05068_, _05067_);
  and _56571_ (_05069_, _05068_, _04485_);
  not _56572_ (_05070_, _05069_);
  nor _56573_ (_05071_, _05070_, _05066_);
  nor _56574_ (_05072_, _04485_, _03756_);
  nor _56575_ (_05073_, _05072_, _05071_);
  nor _56576_ (_05074_, _05073_, _04502_);
  or _56577_ (_05075_, _05074_, _04500_);
  nor _56578_ (_05076_, _05075_, _05006_);
  and _56579_ (_05077_, _04500_, _03756_);
  nor _56580_ (_05078_, _05077_, _05076_);
  nor _56581_ (_05079_, _05078_, _03178_);
  and _56582_ (_05080_, _05012_, _03178_);
  not _56583_ (_05081_, _05080_);
  and _56584_ (_05082_, _05081_, _04517_);
  not _56585_ (_05083_, _05082_);
  nor _56586_ (_05084_, _05083_, _05079_);
  nor _56587_ (_05085_, _04517_, _03756_);
  nor _56588_ (_05086_, _05085_, _03192_);
  not _56589_ (_05087_, _05086_);
  nor _56590_ (_05088_, _05087_, _05084_);
  and _56591_ (_05089_, _05012_, _03192_);
  or _56592_ (_05090_, _05089_, _04524_);
  nor _56593_ (_05091_, _05090_, _05088_);
  and _56594_ (_05092_, _04524_, _03581_);
  or _56595_ (_05093_, _05092_, _03188_);
  nor _56596_ (_05094_, _05093_, _05091_);
  and _56597_ (_05095_, _05012_, _03188_);
  nor _56598_ (_05096_, _05095_, _04533_);
  not _56599_ (_05097_, _05096_);
  nor _56600_ (_05098_, _05097_, _05094_);
  and _56601_ (_05099_, _05005_, _04533_);
  nor _56602_ (_05100_, _05099_, _04531_);
  not _56603_ (_05101_, _05100_);
  nor _56604_ (_05102_, _05101_, _05098_);
  not _56605_ (_05103_, _04540_);
  and _56606_ (_05104_, _04531_, _03756_);
  nor _56607_ (_05105_, _05104_, _05103_);
  not _56608_ (_05106_, _05105_);
  nor _56609_ (_05107_, _05106_, _05102_);
  nor _56610_ (_05108_, _05012_, _04540_);
  nor _56611_ (_05109_, _05108_, _04539_);
  not _56612_ (_05110_, _05109_);
  nor _56613_ (_05111_, _05110_, _05107_);
  not _56614_ (_05112_, _03549_);
  and _56615_ (_05113_, _04539_, _05112_);
  nor _56616_ (_05114_, _05113_, _04552_);
  not _56617_ (_05115_, _05114_);
  nor _56618_ (_05116_, _05115_, _05111_);
  and _56619_ (_05117_, _05005_, _04552_);
  nor _56620_ (_05118_, _05117_, _03448_);
  not _56621_ (_05119_, _05118_);
  nor _56622_ (_05120_, _05119_, _05116_);
  and _56623_ (_05121_, _03827_, _03446_);
  nor _56624_ (_05122_, _05121_, _05120_);
  nor _56625_ (_05123_, _04797_, _05122_);
  and _56626_ (_05124_, _05123_, _04952_);
  and _56627_ (_05125_, _05124_, _04799_);
  or _56628_ (_05126_, _05125_, \oc8051_golden_model_1.IRAM[15] [7]);
  and _56629_ (_05127_, _05009_, _03498_);
  nor _56630_ (_05128_, _04807_, _03499_);
  nor _56631_ (_05129_, _05128_, _05127_);
  and _56632_ (_05130_, _05127_, _03722_);
  nor _56633_ (_05131_, _05010_, _05008_);
  nor _56634_ (_05132_, _05131_, _05130_);
  not _56635_ (_05133_, _05132_);
  and _56636_ (_05134_, _04769_, _04763_);
  and _56637_ (_05135_, _05134_, _04767_);
  and _56638_ (_05136_, _05135_, _04735_);
  nor _56639_ (_05137_, _05136_, _04795_);
  and _56640_ (_05138_, _05137_, _05133_);
  and _56641_ (_05139_, _05138_, _05129_);
  and _56642_ (_05140_, _05139_, _03497_);
  not _56643_ (_05141_, _05140_);
  and _56644_ (_05142_, _05141_, _05126_);
  not _56645_ (_05143_, _05125_);
  not _56646_ (_05144_, \oc8051_golden_model_1.IRAM[0] [7]);
  or _56647_ (_05145_, _04261_, _05144_);
  not _56648_ (_05146_, \oc8051_golden_model_1.IRAM[1] [7]);
  or _56649_ (_05147_, _04348_, _05146_);
  and _56650_ (_05148_, _05147_, _04346_);
  nand _56651_ (_05149_, _05148_, _05145_);
  not _56652_ (_05150_, \oc8051_golden_model_1.IRAM[3] [7]);
  or _56653_ (_05151_, _04348_, _05150_);
  not _56654_ (_05152_, \oc8051_golden_model_1.IRAM[2] [7]);
  or _56655_ (_05153_, _04261_, _05152_);
  and _56656_ (_05154_, _05153_, _04354_);
  nand _56657_ (_05155_, _05154_, _05151_);
  nand _56658_ (_05156_, _05155_, _05149_);
  nand _56659_ (_05157_, _05156_, _04016_);
  not _56660_ (_05158_, \oc8051_golden_model_1.IRAM[7] [7]);
  or _56661_ (_05159_, _04348_, _05158_);
  not _56662_ (_05160_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _56663_ (_05161_, _04261_, _05160_);
  and _56664_ (_05162_, _05161_, _04354_);
  nand _56665_ (_05163_, _05162_, _05159_);
  not _56666_ (_05164_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _56667_ (_05165_, _04261_, _05164_);
  not _56668_ (_05166_, \oc8051_golden_model_1.IRAM[5] [7]);
  or _56669_ (_05167_, _04348_, _05166_);
  and _56670_ (_05168_, _05167_, _04346_);
  nand _56671_ (_05169_, _05168_, _05165_);
  nand _56672_ (_05170_, _05169_, _05163_);
  nand _56673_ (_05171_, _05170_, _04361_);
  nand _56674_ (_05172_, _05171_, _05157_);
  nand _56675_ (_05173_, _05172_, _03829_);
  not _56676_ (_05174_, \oc8051_golden_model_1.IRAM[11] [7]);
  or _56677_ (_05175_, _04348_, _05174_);
  not _56678_ (_05176_, \oc8051_golden_model_1.IRAM[10] [7]);
  or _56679_ (_05177_, _04261_, _05176_);
  and _56680_ (_05178_, _05177_, _04354_);
  nand _56681_ (_05179_, _05178_, _05175_);
  not _56682_ (_05180_, \oc8051_golden_model_1.IRAM[8] [7]);
  or _56683_ (_05181_, _04261_, _05180_);
  not _56684_ (_05182_, \oc8051_golden_model_1.IRAM[9] [7]);
  or _56685_ (_05183_, _04348_, _05182_);
  and _56686_ (_05184_, _05183_, _04346_);
  nand _56687_ (_05185_, _05184_, _05181_);
  nand _56688_ (_05186_, _05185_, _05179_);
  nand _56689_ (_05187_, _05186_, _04016_);
  not _56690_ (_05188_, \oc8051_golden_model_1.IRAM[15] [7]);
  or _56691_ (_05189_, _04348_, _05188_);
  not _56692_ (_05190_, \oc8051_golden_model_1.IRAM[14] [7]);
  or _56693_ (_05191_, _04261_, _05190_);
  and _56694_ (_05192_, _05191_, _04354_);
  nand _56695_ (_05193_, _05192_, _05189_);
  not _56696_ (_05194_, \oc8051_golden_model_1.IRAM[12] [7]);
  or _56697_ (_05195_, _04261_, _05194_);
  not _56698_ (_05196_, \oc8051_golden_model_1.IRAM[13] [7]);
  or _56699_ (_05197_, _04348_, _05196_);
  and _56700_ (_05198_, _05197_, _04346_);
  nand _56701_ (_05199_, _05198_, _05195_);
  nand _56702_ (_05200_, _05199_, _05193_);
  nand _56703_ (_05201_, _05200_, _04361_);
  nand _56704_ (_05202_, _05201_, _05187_);
  nand _56705_ (_05203_, _05202_, _04379_);
  nand _56706_ (_05204_, _05203_, _05173_);
  or _56707_ (_05205_, _05204_, _03454_);
  and _56708_ (_05206_, _03549_, _03454_);
  and _56709_ (_05207_, _05206_, _03860_);
  and _56710_ (_05208_, _05207_, _03486_);
  and _56711_ (_05209_, _05208_, _03581_);
  nor _56712_ (_05210_, _03414_, _04048_);
  and _56713_ (_05211_, _05210_, _04800_);
  and _56714_ (_05212_, _05211_, _05209_);
  and _56715_ (_05213_, _05212_, \oc8051_golden_model_1.PCON [7]);
  not _56716_ (_05214_, _05213_);
  and _56717_ (_05215_, _03414_, _04188_);
  and _56718_ (_05216_, _05215_, _03904_);
  and _56719_ (_05217_, _05216_, _03756_);
  not _56720_ (_05218_, _03486_);
  and _56721_ (_05219_, _05218_, _03860_);
  and _56722_ (_05220_, _05219_, _05206_);
  and _56723_ (_05221_, _05220_, _05217_);
  and _56724_ (_05222_, _05221_, \oc8051_golden_model_1.SBUF [7]);
  and _56725_ (_05223_, _03414_, _04048_);
  and _56726_ (_05224_, _05223_, _03904_);
  and _56727_ (_05225_, _05224_, _03756_);
  not _56728_ (_05226_, _03860_);
  and _56729_ (_05227_, _03486_, _05226_);
  and _56730_ (_05228_, _05227_, _05206_);
  and _56731_ (_05229_, _05228_, _05225_);
  and _56732_ (_05230_, _05229_, \oc8051_golden_model_1.IE [7]);
  nor _56733_ (_05231_, _05230_, _05222_);
  and _56734_ (_05232_, _05231_, _05214_);
  and _56735_ (_05233_, _03904_, _03581_);
  and _56736_ (_05234_, _05233_, _05223_);
  and _56737_ (_05235_, _05234_, _05228_);
  and _56738_ (_05236_, _05235_, \oc8051_golden_model_1.P2 [7]);
  nor _56739_ (_05237_, _03486_, _03860_);
  and _56740_ (_05238_, _05237_, _05206_);
  and _56741_ (_05239_, _05238_, _05234_);
  and _56742_ (_05240_, _05239_, \oc8051_golden_model_1.P3 [7]);
  nor _56743_ (_05241_, _05240_, _05236_);
  and _56744_ (_05242_, _05241_, _05232_);
  nor _56745_ (_05243_, _03549_, _03446_);
  and _56746_ (_05244_, _05243_, _05219_);
  and _56747_ (_05245_, _05244_, _05234_);
  and _56748_ (_05246_, _05245_, \oc8051_golden_model_1.PSW [7]);
  and _56749_ (_05247_, _05243_, _05237_);
  and _56750_ (_05248_, _05247_, _05234_);
  and _56751_ (_05249_, _05248_, \oc8051_golden_model_1.B [7]);
  nor _56752_ (_05250_, _05249_, _05246_);
  and _56753_ (_05251_, _05238_, _05225_);
  and _56754_ (_05252_, _05251_, \oc8051_golden_model_1.IP [7]);
  and _56755_ (_05253_, _05243_, _05227_);
  and _56756_ (_05254_, _05253_, _05234_);
  and _56757_ (_05255_, _05254_, \oc8051_golden_model_1.ACC [7]);
  nor _56758_ (_05256_, _05255_, _05252_);
  and _56759_ (_05257_, _05256_, _05250_);
  and _56760_ (_05258_, _05225_, _05208_);
  and _56761_ (_05259_, _05258_, \oc8051_golden_model_1.TCON [7]);
  not _56762_ (_05260_, _05208_);
  nor _56763_ (_05261_, _03904_, _03581_);
  nand _56764_ (_05262_, _05261_, _05223_);
  nor _56765_ (_05263_, _05262_, _05260_);
  and _56766_ (_05264_, _05263_, \oc8051_golden_model_1.TH0 [7]);
  nor _56767_ (_05265_, _05264_, _05259_);
  and _56768_ (_05266_, _05234_, _05220_);
  and _56769_ (_05267_, _05266_, \oc8051_golden_model_1.P1 [7]);
  not _56770_ (_05268_, _05210_);
  nand _56771_ (_05269_, _03904_, _03756_);
  or _56772_ (_05270_, _05269_, _05268_);
  nor _56773_ (_05271_, _05270_, _05260_);
  and _56774_ (_05272_, _05271_, \oc8051_golden_model_1.TL1 [7]);
  nor _56775_ (_05273_, _05272_, _05267_);
  and _56776_ (_05274_, _05273_, _05265_);
  and _56777_ (_05275_, _05225_, _05220_);
  and _56778_ (_05276_, _05275_, \oc8051_golden_model_1.SCON [7]);
  nand _56779_ (_05277_, _05261_, _05215_);
  nor _56780_ (_05278_, _05277_, _05260_);
  and _56781_ (_05279_, _05278_, \oc8051_golden_model_1.TH1 [7]);
  nor _56782_ (_05280_, _05279_, _05276_);
  nor _56783_ (_05281_, _03414_, _04188_);
  not _56784_ (_05282_, _05281_);
  or _56785_ (_05283_, _05282_, _05269_);
  nor _56786_ (_05284_, _05283_, _05260_);
  and _56787_ (_05285_, _05284_, \oc8051_golden_model_1.TL0 [7]);
  and _56788_ (_05286_, _05217_, _05208_);
  and _56789_ (_05287_, _05286_, \oc8051_golden_model_1.TMOD [7]);
  nor _56790_ (_05288_, _05287_, _05285_);
  and _56791_ (_05289_, _05288_, _05280_);
  and _56792_ (_05290_, _05289_, _05274_);
  and _56793_ (_05291_, _05290_, _05257_);
  and _56794_ (_05292_, _05291_, _05242_);
  and _56795_ (_05293_, _05234_, _05208_);
  and _56796_ (_05294_, _05293_, \oc8051_golden_model_1.P0 [7]);
  not _56797_ (_05295_, _05294_);
  and _56798_ (_05296_, _05210_, _03904_);
  and _56799_ (_05297_, _05296_, _05209_);
  and _56800_ (_05298_, _05297_, \oc8051_golden_model_1.DPH [7]);
  not _56801_ (_05299_, _05298_);
  and _56802_ (_05300_, _05216_, _05209_);
  and _56803_ (_05301_, _05300_, \oc8051_golden_model_1.SP [7]);
  and _56804_ (_05302_, _05281_, _03904_);
  and _56805_ (_05303_, _05302_, _05209_);
  and _56806_ (_05304_, _05303_, \oc8051_golden_model_1.DPL [7]);
  nor _56807_ (_05305_, _05304_, _05301_);
  and _56808_ (_05306_, _05305_, _05299_);
  and _56809_ (_05307_, _05306_, _05295_);
  and _56810_ (_05308_, _05307_, _05292_);
  and _56811_ (_05309_, _05308_, _05205_);
  not _56812_ (_05310_, _05309_);
  not _56813_ (_05311_, \oc8051_golden_model_1.IRAM[0] [6]);
  or _56814_ (_05312_, _04261_, _05311_);
  not _56815_ (_05313_, \oc8051_golden_model_1.IRAM[1] [6]);
  or _56816_ (_05314_, _04348_, _05313_);
  and _56817_ (_05315_, _05314_, _04346_);
  nand _56818_ (_05316_, _05315_, _05312_);
  not _56819_ (_05317_, \oc8051_golden_model_1.IRAM[3] [6]);
  or _56820_ (_05318_, _04348_, _05317_);
  not _56821_ (_05319_, \oc8051_golden_model_1.IRAM[2] [6]);
  or _56822_ (_05320_, _04261_, _05319_);
  and _56823_ (_05321_, _05320_, _04354_);
  nand _56824_ (_05322_, _05321_, _05318_);
  nand _56825_ (_05323_, _05322_, _05316_);
  nand _56826_ (_05324_, _05323_, _04016_);
  not _56827_ (_05325_, \oc8051_golden_model_1.IRAM[7] [6]);
  or _56828_ (_05326_, _04348_, _05325_);
  not _56829_ (_05327_, \oc8051_golden_model_1.IRAM[6] [6]);
  or _56830_ (_05328_, _04261_, _05327_);
  and _56831_ (_05329_, _05328_, _04354_);
  nand _56832_ (_05330_, _05329_, _05326_);
  not _56833_ (_05331_, \oc8051_golden_model_1.IRAM[4] [6]);
  or _56834_ (_05332_, _04261_, _05331_);
  not _56835_ (_05333_, \oc8051_golden_model_1.IRAM[5] [6]);
  or _56836_ (_05334_, _04348_, _05333_);
  and _56837_ (_05335_, _05334_, _04346_);
  nand _56838_ (_05336_, _05335_, _05332_);
  nand _56839_ (_05337_, _05336_, _05330_);
  nand _56840_ (_05338_, _05337_, _04361_);
  nand _56841_ (_05339_, _05338_, _05324_);
  nand _56842_ (_05340_, _05339_, _03829_);
  nand _56843_ (_05341_, _04261_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _56844_ (_05342_, _04348_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _56845_ (_05343_, _05342_, _04354_);
  nand _56846_ (_05344_, _05343_, _05341_);
  nand _56847_ (_05345_, _04348_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand _56848_ (_05346_, _04261_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _56849_ (_05347_, _05346_, _04346_);
  nand _56850_ (_05348_, _05347_, _05345_);
  nand _56851_ (_05349_, _05348_, _05344_);
  nand _56852_ (_05350_, _05349_, _04016_);
  nand _56853_ (_05351_, _04261_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _56854_ (_05352_, _04348_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _56855_ (_05353_, _05352_, _04354_);
  nand _56856_ (_05354_, _05353_, _05351_);
  nand _56857_ (_05355_, _04348_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand _56858_ (_05356_, _04261_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _56859_ (_05357_, _05356_, _04346_);
  nand _56860_ (_05358_, _05357_, _05355_);
  nand _56861_ (_05359_, _05358_, _05354_);
  nand _56862_ (_05360_, _05359_, _04361_);
  nand _56863_ (_05361_, _05360_, _05350_);
  nand _56864_ (_05362_, _05361_, _04379_);
  nand _56865_ (_05363_, _05362_, _05340_);
  or _56866_ (_05364_, _05363_, _03454_);
  and _56867_ (_05365_, _05297_, \oc8051_golden_model_1.DPH [6]);
  not _56868_ (_05366_, _05365_);
  and _56869_ (_05367_, _05263_, \oc8051_golden_model_1.TH0 [6]);
  and _56870_ (_05368_, _05271_, \oc8051_golden_model_1.TL1 [6]);
  nor _56871_ (_05369_, _05368_, _05367_);
  and _56872_ (_05370_, _05369_, _05366_);
  and _56873_ (_05371_, _05300_, \oc8051_golden_model_1.SP [6]);
  and _56874_ (_05372_, _05303_, \oc8051_golden_model_1.DPL [6]);
  nor _56875_ (_05373_, _05372_, _05371_);
  and _56876_ (_05374_, _05212_, \oc8051_golden_model_1.PCON [6]);
  not _56877_ (_05375_, _05374_);
  and _56878_ (_05376_, _05221_, \oc8051_golden_model_1.SBUF [6]);
  and _56879_ (_05377_, _05229_, \oc8051_golden_model_1.IE [6]);
  nor _56880_ (_05378_, _05377_, _05376_);
  and _56881_ (_05379_, _05378_, _05375_);
  and _56882_ (_05380_, _05379_, _05373_);
  and _56883_ (_05381_, _05380_, _05370_);
  and _56884_ (_05382_, _05284_, \oc8051_golden_model_1.TL0 [6]);
  and _56885_ (_05383_, _05275_, \oc8051_golden_model_1.SCON [6]);
  nor _56886_ (_05384_, _05383_, _05382_);
  and _56887_ (_05385_, _05278_, \oc8051_golden_model_1.TH1 [6]);
  not _56888_ (_05386_, _05385_);
  and _56889_ (_05387_, _05258_, \oc8051_golden_model_1.TCON [6]);
  and _56890_ (_05388_, _05286_, \oc8051_golden_model_1.TMOD [6]);
  nor _56891_ (_05389_, _05388_, _05387_);
  and _56892_ (_05390_, _05389_, _05386_);
  and _56893_ (_05391_, _05390_, _05384_);
  and _56894_ (_05392_, _05251_, \oc8051_golden_model_1.IP [6]);
  and _56895_ (_05393_, _05248_, \oc8051_golden_model_1.B [6]);
  nor _56896_ (_05394_, _05393_, _05392_);
  and _56897_ (_05395_, _05245_, \oc8051_golden_model_1.PSW [6]);
  and _56898_ (_05396_, _05254_, \oc8051_golden_model_1.ACC [6]);
  nor _56899_ (_05397_, _05396_, _05395_);
  and _56900_ (_05398_, _05397_, _05394_);
  and _56901_ (_05399_, _05293_, \oc8051_golden_model_1.P0 [6]);
  not _56902_ (_05400_, _05399_);
  and _56903_ (_05401_, _05266_, \oc8051_golden_model_1.P1 [6]);
  not _56904_ (_05402_, _05401_);
  and _56905_ (_05403_, _05235_, \oc8051_golden_model_1.P2 [6]);
  and _56906_ (_05404_, _05239_, \oc8051_golden_model_1.P3 [6]);
  nor _56907_ (_05405_, _05404_, _05403_);
  and _56908_ (_05406_, _05405_, _05402_);
  and _56909_ (_05407_, _05406_, _05400_);
  and _56910_ (_05408_, _05407_, _05398_);
  and _56911_ (_05409_, _05408_, _05391_);
  and _56912_ (_05410_, _05409_, _05381_);
  and _56913_ (_05411_, _05410_, _05364_);
  not _56914_ (_05412_, _05411_);
  not _56915_ (_05413_, \oc8051_golden_model_1.IRAM[0] [5]);
  or _56916_ (_05414_, _04261_, _05413_);
  not _56917_ (_05415_, \oc8051_golden_model_1.IRAM[1] [5]);
  or _56918_ (_05416_, _04348_, _05415_);
  and _56919_ (_05417_, _05416_, _04346_);
  nand _56920_ (_05418_, _05417_, _05414_);
  not _56921_ (_05419_, \oc8051_golden_model_1.IRAM[3] [5]);
  or _56922_ (_05420_, _04348_, _05419_);
  not _56923_ (_05421_, \oc8051_golden_model_1.IRAM[2] [5]);
  or _56924_ (_05422_, _04261_, _05421_);
  and _56925_ (_05423_, _05422_, _04354_);
  nand _56926_ (_05424_, _05423_, _05420_);
  nand _56927_ (_05425_, _05424_, _05418_);
  nand _56928_ (_05426_, _05425_, _04016_);
  not _56929_ (_05427_, \oc8051_golden_model_1.IRAM[7] [5]);
  or _56930_ (_05428_, _04348_, _05427_);
  not _56931_ (_05429_, \oc8051_golden_model_1.IRAM[6] [5]);
  or _56932_ (_05430_, _04261_, _05429_);
  and _56933_ (_05431_, _05430_, _04354_);
  nand _56934_ (_05432_, _05431_, _05428_);
  not _56935_ (_05433_, \oc8051_golden_model_1.IRAM[4] [5]);
  or _56936_ (_05434_, _04261_, _05433_);
  not _56937_ (_05435_, \oc8051_golden_model_1.IRAM[5] [5]);
  or _56938_ (_05436_, _04348_, _05435_);
  and _56939_ (_05437_, _05436_, _04346_);
  nand _56940_ (_05438_, _05437_, _05434_);
  nand _56941_ (_05439_, _05438_, _05432_);
  nand _56942_ (_05440_, _05439_, _04361_);
  nand _56943_ (_05441_, _05440_, _05426_);
  nand _56944_ (_05442_, _05441_, _03829_);
  nand _56945_ (_05443_, _04261_, \oc8051_golden_model_1.IRAM[11] [5]);
  not _56946_ (_05444_, \oc8051_golden_model_1.IRAM[10] [5]);
  or _56947_ (_05445_, _04261_, _05444_);
  and _56948_ (_05446_, _05445_, _04354_);
  nand _56949_ (_05447_, _05446_, _05443_);
  nand _56950_ (_05448_, _04348_, \oc8051_golden_model_1.IRAM[8] [5]);
  not _56951_ (_05449_, \oc8051_golden_model_1.IRAM[9] [5]);
  or _56952_ (_05450_, _04348_, _05449_);
  and _56953_ (_05451_, _05450_, _04346_);
  nand _56954_ (_05452_, _05451_, _05448_);
  nand _56955_ (_05453_, _05452_, _05447_);
  nand _56956_ (_05454_, _05453_, _04016_);
  nand _56957_ (_05455_, _04261_, \oc8051_golden_model_1.IRAM[15] [5]);
  not _56958_ (_05456_, \oc8051_golden_model_1.IRAM[14] [5]);
  or _56959_ (_05457_, _04261_, _05456_);
  and _56960_ (_05458_, _05457_, _04354_);
  nand _56961_ (_05459_, _05458_, _05455_);
  nand _56962_ (_05460_, _04348_, \oc8051_golden_model_1.IRAM[12] [5]);
  not _56963_ (_05461_, \oc8051_golden_model_1.IRAM[13] [5]);
  or _56964_ (_05462_, _04348_, _05461_);
  and _56965_ (_05463_, _05462_, _04346_);
  nand _56966_ (_05464_, _05463_, _05460_);
  nand _56967_ (_05465_, _05464_, _05459_);
  nand _56968_ (_05466_, _05465_, _04361_);
  nand _56969_ (_05467_, _05466_, _05454_);
  nand _56970_ (_05468_, _05467_, _04379_);
  nand _56971_ (_05469_, _05468_, _05442_);
  or _56972_ (_05470_, _05469_, _03454_);
  and _56973_ (_05471_, _05297_, \oc8051_golden_model_1.DPH [5]);
  not _56974_ (_05472_, _05471_);
  and _56975_ (_05473_, _05300_, \oc8051_golden_model_1.SP [5]);
  and _56976_ (_05474_, _05303_, \oc8051_golden_model_1.DPL [5]);
  nor _56977_ (_05475_, _05474_, _05473_);
  and _56978_ (_05476_, _05475_, _05472_);
  and _56979_ (_05477_, _05258_, \oc8051_golden_model_1.TCON [5]);
  not _56980_ (_05478_, _05477_);
  and _56981_ (_05479_, _05284_, \oc8051_golden_model_1.TL0 [5]);
  and _56982_ (_05480_, _05275_, \oc8051_golden_model_1.SCON [5]);
  nor _56983_ (_05481_, _05480_, _05479_);
  and _56984_ (_05482_, _05481_, _05478_);
  and _56985_ (_05483_, _05263_, \oc8051_golden_model_1.TH0 [5]);
  and _56986_ (_05484_, _05278_, \oc8051_golden_model_1.TH1 [5]);
  nor _56987_ (_05485_, _05484_, _05483_);
  and _56988_ (_05486_, _05286_, \oc8051_golden_model_1.TMOD [5]);
  and _56989_ (_05487_, _05271_, \oc8051_golden_model_1.TL1 [5]);
  nor _56990_ (_05488_, _05487_, _05486_);
  and _56991_ (_05489_, _05488_, _05485_);
  and _56992_ (_05490_, _05489_, _05482_);
  and _56993_ (_05491_, _05490_, _05476_);
  and _56994_ (_05492_, _05212_, \oc8051_golden_model_1.PCON [5]);
  not _56995_ (_05493_, _05492_);
  and _56996_ (_05494_, _05221_, \oc8051_golden_model_1.SBUF [5]);
  and _56997_ (_05495_, _05229_, \oc8051_golden_model_1.IE [5]);
  nor _56998_ (_05496_, _05495_, _05494_);
  and _56999_ (_05497_, _05496_, _05493_);
  and _57000_ (_05498_, _05293_, \oc8051_golden_model_1.P0 [5]);
  not _57001_ (_05499_, _05498_);
  and _57002_ (_05500_, _05245_, \oc8051_golden_model_1.PSW [5]);
  and _57003_ (_05501_, _05254_, \oc8051_golden_model_1.ACC [5]);
  nor _57004_ (_05502_, _05501_, _05500_);
  and _57005_ (_05503_, _05251_, \oc8051_golden_model_1.IP [5]);
  and _57006_ (_05504_, _05248_, \oc8051_golden_model_1.B [5]);
  nor _57007_ (_05505_, _05504_, _05503_);
  and _57008_ (_05506_, _05505_, _05502_);
  and _57009_ (_05507_, _05266_, \oc8051_golden_model_1.P1 [5]);
  not _57010_ (_05508_, _05507_);
  and _57011_ (_05509_, _05235_, \oc8051_golden_model_1.P2 [5]);
  and _57012_ (_05510_, _05239_, \oc8051_golden_model_1.P3 [5]);
  nor _57013_ (_05511_, _05510_, _05509_);
  and _57014_ (_05512_, _05511_, _05508_);
  and _57015_ (_05513_, _05512_, _05506_);
  and _57016_ (_05514_, _05513_, _05499_);
  and _57017_ (_05515_, _05514_, _05497_);
  and _57018_ (_05516_, _05515_, _05491_);
  and _57019_ (_05517_, _05516_, _05470_);
  not _57020_ (_05518_, _05517_);
  or _57021_ (_05519_, _05005_, _03454_);
  and _57022_ (_05520_, _05297_, \oc8051_golden_model_1.DPH [3]);
  not _57023_ (_05521_, _05520_);
  and _57024_ (_05522_, _05300_, \oc8051_golden_model_1.SP [3]);
  and _57025_ (_05523_, _05303_, \oc8051_golden_model_1.DPL [3]);
  nor _57026_ (_05524_, _05523_, _05522_);
  and _57027_ (_05525_, _05524_, _05521_);
  and _57028_ (_05526_, _05258_, \oc8051_golden_model_1.TCON [3]);
  not _57029_ (_05527_, _05526_);
  and _57030_ (_05528_, _05284_, \oc8051_golden_model_1.TL0 [3]);
  and _57031_ (_05529_, _05275_, \oc8051_golden_model_1.SCON [3]);
  nor _57032_ (_05530_, _05529_, _05528_);
  and _57033_ (_05531_, _05530_, _05527_);
  and _57034_ (_05532_, _05263_, \oc8051_golden_model_1.TH0 [3]);
  and _57035_ (_05533_, _05278_, \oc8051_golden_model_1.TH1 [3]);
  nor _57036_ (_05534_, _05533_, _05532_);
  and _57037_ (_05535_, _05286_, \oc8051_golden_model_1.TMOD [3]);
  and _57038_ (_05536_, _05271_, \oc8051_golden_model_1.TL1 [3]);
  nor _57039_ (_05537_, _05536_, _05535_);
  and _57040_ (_05538_, _05537_, _05534_);
  and _57041_ (_05539_, _05538_, _05531_);
  and _57042_ (_05540_, _05539_, _05525_);
  and _57043_ (_05541_, _05212_, \oc8051_golden_model_1.PCON [3]);
  not _57044_ (_05542_, _05541_);
  and _57045_ (_05543_, _05221_, \oc8051_golden_model_1.SBUF [3]);
  and _57046_ (_05544_, _05229_, \oc8051_golden_model_1.IE [3]);
  nor _57047_ (_05545_, _05544_, _05543_);
  and _57048_ (_05546_, _05545_, _05542_);
  and _57049_ (_05547_, _05293_, \oc8051_golden_model_1.P0 [3]);
  not _57050_ (_05548_, _05547_);
  and _57051_ (_05549_, _05245_, \oc8051_golden_model_1.PSW [3]);
  and _57052_ (_05550_, _05248_, \oc8051_golden_model_1.B [3]);
  nor _57053_ (_05551_, _05550_, _05549_);
  and _57054_ (_05552_, _05251_, \oc8051_golden_model_1.IP [3]);
  and _57055_ (_05553_, _05254_, \oc8051_golden_model_1.ACC [3]);
  nor _57056_ (_05554_, _05553_, _05552_);
  and _57057_ (_05555_, _05554_, _05551_);
  and _57058_ (_05556_, _05266_, \oc8051_golden_model_1.P1 [3]);
  not _57059_ (_05557_, _05556_);
  and _57060_ (_05558_, _05235_, \oc8051_golden_model_1.P2 [3]);
  and _57061_ (_05559_, _05239_, \oc8051_golden_model_1.P3 [3]);
  nor _57062_ (_05560_, _05559_, _05558_);
  and _57063_ (_05561_, _05560_, _05557_);
  and _57064_ (_05562_, _05561_, _05555_);
  and _57065_ (_05563_, _05562_, _05548_);
  and _57066_ (_05564_, _05563_, _05546_);
  and _57067_ (_05565_, _05564_, _05540_);
  and _57068_ (_05566_, _05565_, _05519_);
  not _57069_ (_05567_, _05566_);
  or _57070_ (_05568_, _04406_, _03454_);
  and _57071_ (_05569_, _05300_, \oc8051_golden_model_1.SP [1]);
  not _57072_ (_05570_, _05569_);
  and _57073_ (_05571_, _05303_, \oc8051_golden_model_1.DPL [1]);
  and _57074_ (_05572_, _05258_, \oc8051_golden_model_1.TCON [1]);
  nor _57075_ (_05573_, _05572_, _05571_);
  and _57076_ (_05574_, _05573_, _05570_);
  and _57077_ (_05575_, _05293_, \oc8051_golden_model_1.P0 [1]);
  not _57078_ (_05576_, _05575_);
  and _57079_ (_05577_, _05266_, \oc8051_golden_model_1.P1 [1]);
  not _57080_ (_05578_, _05577_);
  and _57081_ (_05579_, _05235_, \oc8051_golden_model_1.P2 [1]);
  and _57082_ (_05580_, _05239_, \oc8051_golden_model_1.P3 [1]);
  nor _57083_ (_05581_, _05580_, _05579_);
  and _57084_ (_05582_, _05581_, _05578_);
  and _57085_ (_05583_, _05582_, _05576_);
  and _57086_ (_05584_, _05583_, _05574_);
  and _57087_ (_05585_, _05271_, \oc8051_golden_model_1.TL1 [1]);
  and _57088_ (_05586_, _05278_, \oc8051_golden_model_1.TH1 [1]);
  nor _57089_ (_05587_, _05586_, _05585_);
  and _57090_ (_05588_, _05286_, \oc8051_golden_model_1.TMOD [1]);
  and _57091_ (_05589_, _05275_, \oc8051_golden_model_1.SCON [1]);
  nor _57092_ (_05590_, _05589_, _05588_);
  and _57093_ (_05591_, _05590_, _05587_);
  and _57094_ (_05592_, _05297_, \oc8051_golden_model_1.DPH [1]);
  not _57095_ (_05593_, _05592_);
  and _57096_ (_05594_, _05284_, \oc8051_golden_model_1.TL0 [1]);
  and _57097_ (_05595_, _05263_, \oc8051_golden_model_1.TH0 [1]);
  nor _57098_ (_05596_, _05595_, _05594_);
  and _57099_ (_05597_, _05596_, _05593_);
  and _57100_ (_05598_, _05597_, _05591_);
  and _57101_ (_05599_, _05212_, \oc8051_golden_model_1.PCON [1]);
  not _57102_ (_05600_, _05599_);
  and _57103_ (_05601_, _05251_, \oc8051_golden_model_1.IP [1]);
  not _57104_ (_05602_, _05601_);
  and _57105_ (_05603_, _05245_, \oc8051_golden_model_1.PSW [1]);
  and _57106_ (_05604_, _05248_, \oc8051_golden_model_1.B [1]);
  nor _57107_ (_05605_, _05604_, _05603_);
  and _57108_ (_05606_, _05605_, _05602_);
  and _57109_ (_05607_, _05221_, \oc8051_golden_model_1.SBUF [1]);
  not _57110_ (_05608_, _05607_);
  and _57111_ (_05609_, _05229_, \oc8051_golden_model_1.IE [1]);
  and _57112_ (_05610_, _05254_, \oc8051_golden_model_1.ACC [1]);
  nor _57113_ (_05611_, _05610_, _05609_);
  and _57114_ (_05612_, _05611_, _05608_);
  and _57115_ (_05613_, _05612_, _05606_);
  and _57116_ (_05614_, _05613_, _05600_);
  and _57117_ (_05615_, _05614_, _05598_);
  and _57118_ (_05616_, _05615_, _05584_);
  and _57119_ (_05617_, _05616_, _05568_);
  not _57120_ (_05618_, _05617_);
  or _57121_ (_05619_, _04634_, _03454_);
  and _57122_ (_05620_, _05297_, \oc8051_golden_model_1.DPH [0]);
  not _57123_ (_05621_, _05620_);
  and _57124_ (_05622_, _05300_, \oc8051_golden_model_1.SP [0]);
  and _57125_ (_05623_, _05303_, \oc8051_golden_model_1.DPL [0]);
  nor _57126_ (_05624_, _05623_, _05622_);
  and _57127_ (_05625_, _05624_, _05621_);
  and _57128_ (_05626_, _05258_, \oc8051_golden_model_1.TCON [0]);
  not _57129_ (_05627_, _05626_);
  and _57130_ (_05628_, _05284_, \oc8051_golden_model_1.TL0 [0]);
  and _57131_ (_05629_, _05275_, \oc8051_golden_model_1.SCON [0]);
  nor _57132_ (_05630_, _05629_, _05628_);
  and _57133_ (_05631_, _05630_, _05627_);
  and _57134_ (_05632_, _05263_, \oc8051_golden_model_1.TH0 [0]);
  and _57135_ (_05633_, _05278_, \oc8051_golden_model_1.TH1 [0]);
  nor _57136_ (_05634_, _05633_, _05632_);
  and _57137_ (_05635_, _05286_, \oc8051_golden_model_1.TMOD [0]);
  and _57138_ (_05636_, _05271_, \oc8051_golden_model_1.TL1 [0]);
  nor _57139_ (_05637_, _05636_, _05635_);
  and _57140_ (_05638_, _05637_, _05634_);
  and _57141_ (_05639_, _05638_, _05631_);
  and _57142_ (_05640_, _05639_, _05625_);
  and _57143_ (_05641_, _05212_, \oc8051_golden_model_1.PCON [0]);
  not _57144_ (_05642_, _05641_);
  and _57145_ (_05643_, _05221_, \oc8051_golden_model_1.SBUF [0]);
  and _57146_ (_05644_, _05229_, \oc8051_golden_model_1.IE [0]);
  nor _57147_ (_05645_, _05644_, _05643_);
  and _57148_ (_05646_, _05645_, _05642_);
  and _57149_ (_05647_, _05293_, \oc8051_golden_model_1.P0 [0]);
  not _57150_ (_05648_, _05647_);
  and _57151_ (_05649_, _05251_, \oc8051_golden_model_1.IP [0]);
  and _57152_ (_05650_, _05248_, \oc8051_golden_model_1.B [0]);
  nor _57153_ (_05651_, _05650_, _05649_);
  and _57154_ (_05652_, _05245_, \oc8051_golden_model_1.PSW [0]);
  and _57155_ (_05653_, _05254_, \oc8051_golden_model_1.ACC [0]);
  nor _57156_ (_05654_, _05653_, _05652_);
  and _57157_ (_05655_, _05654_, _05651_);
  and _57158_ (_05656_, _05266_, \oc8051_golden_model_1.P1 [0]);
  not _57159_ (_05657_, _05656_);
  and _57160_ (_05658_, _05235_, \oc8051_golden_model_1.P2 [0]);
  and _57161_ (_05659_, _05239_, \oc8051_golden_model_1.P3 [0]);
  nor _57162_ (_05660_, _05659_, _05658_);
  and _57163_ (_05661_, _05660_, _05657_);
  and _57164_ (_05662_, _05661_, _05655_);
  and _57165_ (_05663_, _05662_, _05648_);
  and _57166_ (_05664_, _05663_, _05646_);
  and _57167_ (_05665_, _05664_, _05640_);
  nand _57168_ (_05666_, _05665_, _05619_);
  and _57169_ (_05667_, _05666_, _05618_);
  or _57170_ (_05668_, _04875_, _03454_);
  and _57171_ (_05669_, _05300_, \oc8051_golden_model_1.SP [2]);
  not _57172_ (_05670_, _05669_);
  and _57173_ (_05671_, _05303_, \oc8051_golden_model_1.DPL [2]);
  and _57174_ (_05672_, _05258_, \oc8051_golden_model_1.TCON [2]);
  nor _57175_ (_05673_, _05672_, _05671_);
  and _57176_ (_05674_, _05673_, _05670_);
  and _57177_ (_05675_, _05293_, \oc8051_golden_model_1.P0 [2]);
  not _57178_ (_05676_, _05675_);
  and _57179_ (_05677_, _05266_, \oc8051_golden_model_1.P1 [2]);
  not _57180_ (_05678_, _05677_);
  and _57181_ (_05679_, _05235_, \oc8051_golden_model_1.P2 [2]);
  and _57182_ (_05680_, _05239_, \oc8051_golden_model_1.P3 [2]);
  nor _57183_ (_05681_, _05680_, _05679_);
  and _57184_ (_05682_, _05681_, _05678_);
  and _57185_ (_05683_, _05682_, _05676_);
  and _57186_ (_05684_, _05683_, _05674_);
  and _57187_ (_05685_, _05271_, \oc8051_golden_model_1.TL1 [2]);
  and _57188_ (_05686_, _05278_, \oc8051_golden_model_1.TH1 [2]);
  nor _57189_ (_05687_, _05686_, _05685_);
  and _57190_ (_05688_, _05286_, \oc8051_golden_model_1.TMOD [2]);
  and _57191_ (_05689_, _05275_, \oc8051_golden_model_1.SCON [2]);
  nor _57192_ (_05690_, _05689_, _05688_);
  and _57193_ (_05691_, _05690_, _05687_);
  and _57194_ (_05692_, _05297_, \oc8051_golden_model_1.DPH [2]);
  not _57195_ (_05693_, _05692_);
  and _57196_ (_05694_, _05284_, \oc8051_golden_model_1.TL0 [2]);
  and _57197_ (_05695_, _05263_, \oc8051_golden_model_1.TH0 [2]);
  nor _57198_ (_05696_, _05695_, _05694_);
  and _57199_ (_05697_, _05696_, _05693_);
  and _57200_ (_05698_, _05697_, _05691_);
  and _57201_ (_05699_, _05212_, \oc8051_golden_model_1.PCON [2]);
  not _57202_ (_05700_, _05699_);
  and _57203_ (_05701_, _05251_, \oc8051_golden_model_1.IP [2]);
  not _57204_ (_05702_, _05701_);
  and _57205_ (_05703_, _05245_, \oc8051_golden_model_1.PSW [2]);
  and _57206_ (_05704_, _05254_, \oc8051_golden_model_1.ACC [2]);
  nor _57207_ (_05705_, _05704_, _05703_);
  and _57208_ (_05706_, _05705_, _05702_);
  and _57209_ (_05707_, _05221_, \oc8051_golden_model_1.SBUF [2]);
  not _57210_ (_05708_, _05707_);
  and _57211_ (_05709_, _05229_, \oc8051_golden_model_1.IE [2]);
  and _57212_ (_05710_, _05248_, \oc8051_golden_model_1.B [2]);
  nor _57213_ (_05711_, _05710_, _05709_);
  and _57214_ (_05712_, _05711_, _05708_);
  and _57215_ (_05713_, _05712_, _05706_);
  and _57216_ (_05714_, _05713_, _05700_);
  and _57217_ (_05715_, _05714_, _05698_);
  and _57218_ (_05716_, _05715_, _05684_);
  and _57219_ (_05717_, _05716_, _05668_);
  not _57220_ (_05718_, _05717_);
  and _57221_ (_05719_, _05718_, _05667_);
  and _57222_ (_05720_, _05719_, _05567_);
  not _57223_ (_05721_, \oc8051_golden_model_1.IRAM[0] [4]);
  or _57224_ (_05722_, _04261_, _05721_);
  not _57225_ (_05723_, \oc8051_golden_model_1.IRAM[1] [4]);
  or _57226_ (_05724_, _04348_, _05723_);
  and _57227_ (_05725_, _05724_, _04346_);
  nand _57228_ (_05726_, _05725_, _05722_);
  not _57229_ (_05727_, \oc8051_golden_model_1.IRAM[3] [4]);
  or _57230_ (_05728_, _04348_, _05727_);
  not _57231_ (_05729_, \oc8051_golden_model_1.IRAM[2] [4]);
  or _57232_ (_05730_, _04261_, _05729_);
  and _57233_ (_05731_, _05730_, _04354_);
  nand _57234_ (_05732_, _05731_, _05728_);
  nand _57235_ (_05733_, _05732_, _05726_);
  nand _57236_ (_05734_, _05733_, _04016_);
  not _57237_ (_05735_, \oc8051_golden_model_1.IRAM[7] [4]);
  or _57238_ (_05736_, _04348_, _05735_);
  not _57239_ (_05737_, \oc8051_golden_model_1.IRAM[6] [4]);
  or _57240_ (_05738_, _04261_, _05737_);
  and _57241_ (_05739_, _05738_, _04354_);
  nand _57242_ (_05740_, _05739_, _05736_);
  not _57243_ (_05741_, \oc8051_golden_model_1.IRAM[4] [4]);
  or _57244_ (_05742_, _04261_, _05741_);
  not _57245_ (_05743_, \oc8051_golden_model_1.IRAM[5] [4]);
  or _57246_ (_05744_, _04348_, _05743_);
  and _57247_ (_05745_, _05744_, _04346_);
  nand _57248_ (_05746_, _05745_, _05742_);
  nand _57249_ (_05747_, _05746_, _05740_);
  nand _57250_ (_05748_, _05747_, _04361_);
  nand _57251_ (_05749_, _05748_, _05734_);
  nand _57252_ (_05750_, _05749_, _03829_);
  nand _57253_ (_05751_, _04261_, \oc8051_golden_model_1.IRAM[11] [4]);
  not _57254_ (_05752_, \oc8051_golden_model_1.IRAM[10] [4]);
  or _57255_ (_05753_, _04261_, _05752_);
  and _57256_ (_05754_, _05753_, _04354_);
  nand _57257_ (_05755_, _05754_, _05751_);
  nand _57258_ (_05756_, _04348_, \oc8051_golden_model_1.IRAM[8] [4]);
  not _57259_ (_05757_, \oc8051_golden_model_1.IRAM[9] [4]);
  or _57260_ (_05758_, _04348_, _05757_);
  and _57261_ (_05759_, _05758_, _04346_);
  nand _57262_ (_05760_, _05759_, _05756_);
  nand _57263_ (_05761_, _05760_, _05755_);
  nand _57264_ (_05762_, _05761_, _04016_);
  nand _57265_ (_05763_, _04261_, \oc8051_golden_model_1.IRAM[15] [4]);
  not _57266_ (_05764_, \oc8051_golden_model_1.IRAM[14] [4]);
  or _57267_ (_05765_, _04261_, _05764_);
  and _57268_ (_05766_, _05765_, _04354_);
  nand _57269_ (_05767_, _05766_, _05763_);
  nand _57270_ (_05768_, _04348_, \oc8051_golden_model_1.IRAM[12] [4]);
  not _57271_ (_05769_, \oc8051_golden_model_1.IRAM[13] [4]);
  or _57272_ (_05770_, _04348_, _05769_);
  and _57273_ (_05771_, _05770_, _04346_);
  nand _57274_ (_05772_, _05771_, _05768_);
  nand _57275_ (_05773_, _05772_, _05767_);
  nand _57276_ (_05774_, _05773_, _04361_);
  nand _57277_ (_05775_, _05774_, _05762_);
  nand _57278_ (_05776_, _05775_, _04379_);
  nand _57279_ (_05777_, _05776_, _05750_);
  or _57280_ (_05778_, _05777_, _03454_);
  and _57281_ (_05779_, _05278_, \oc8051_golden_model_1.TH1 [4]);
  and _57282_ (_05780_, _05221_, \oc8051_golden_model_1.SBUF [4]);
  nor _57283_ (_05781_, _05780_, _05779_);
  and _57284_ (_05782_, _05286_, \oc8051_golden_model_1.TMOD [4]);
  and _57285_ (_05783_, _05275_, \oc8051_golden_model_1.SCON [4]);
  nor _57286_ (_05784_, _05783_, _05782_);
  and _57287_ (_05785_, _05784_, _05781_);
  and _57288_ (_05786_, _05303_, \oc8051_golden_model_1.DPL [4]);
  not _57289_ (_05787_, _05786_);
  and _57290_ (_05788_, _05284_, \oc8051_golden_model_1.TL0 [4]);
  and _57291_ (_05789_, _05229_, \oc8051_golden_model_1.IE [4]);
  nor _57292_ (_05790_, _05789_, _05788_);
  and _57293_ (_05791_, _05790_, _05787_);
  and _57294_ (_05792_, _05300_, \oc8051_golden_model_1.SP [4]);
  and _57295_ (_05793_, _05297_, \oc8051_golden_model_1.DPH [4]);
  nor _57296_ (_05794_, _05793_, _05792_);
  and _57297_ (_05795_, _05794_, _05791_);
  and _57298_ (_05796_, _05795_, _05785_);
  not _57299_ (_05797_, _05796_);
  and _57300_ (_05798_, _05266_, \oc8051_golden_model_1.P1 [4]);
  and _57301_ (_05799_, _05258_, \oc8051_golden_model_1.TCON [4]);
  and _57302_ (_05800_, _05235_, \oc8051_golden_model_1.P2 [4]);
  and _57303_ (_05801_, _05239_, \oc8051_golden_model_1.P3 [4]);
  or _57304_ (_05802_, _05801_, _05800_);
  or _57305_ (_05803_, _05802_, _05799_);
  or _57306_ (_05804_, _05803_, _05798_);
  and _57307_ (_05805_, _05212_, \oc8051_golden_model_1.PCON [4]);
  not _57308_ (_05806_, _05805_);
  and _57309_ (_05807_, _05245_, \oc8051_golden_model_1.PSW [4]);
  and _57310_ (_05808_, _05248_, \oc8051_golden_model_1.B [4]);
  nor _57311_ (_05809_, _05808_, _05807_);
  and _57312_ (_05810_, _05251_, \oc8051_golden_model_1.IP [4]);
  and _57313_ (_05811_, _05254_, \oc8051_golden_model_1.ACC [4]);
  nor _57314_ (_05812_, _05811_, _05810_);
  and _57315_ (_05813_, _05812_, _05809_);
  and _57316_ (_05814_, _05813_, _05806_);
  and _57317_ (_05815_, _05293_, \oc8051_golden_model_1.P0 [4]);
  not _57318_ (_05816_, _05815_);
  and _57319_ (_05817_, _05263_, \oc8051_golden_model_1.TH0 [4]);
  and _57320_ (_05818_, _05271_, \oc8051_golden_model_1.TL1 [4]);
  nor _57321_ (_05819_, _05818_, _05817_);
  and _57322_ (_05820_, _05819_, _05816_);
  nand _57323_ (_05821_, _05820_, _05814_);
  or _57324_ (_05822_, _05821_, _05804_);
  nor _57325_ (_05823_, _05822_, _05797_);
  and _57326_ (_05824_, _05823_, _05778_);
  not _57327_ (_05825_, _05824_);
  and _57328_ (_05826_, _05825_, _05720_);
  and _57329_ (_05827_, _05826_, _05518_);
  and _57330_ (_05828_, _05827_, _05412_);
  nor _57331_ (_05829_, _05828_, _05310_);
  and _57332_ (_05830_, _05828_, _05310_);
  nor _57333_ (_05831_, _05830_, _05829_);
  and _57334_ (_05832_, _05831_, _03448_);
  not _57335_ (_05833_, _05204_);
  and _57336_ (_05834_, _05777_, _05469_);
  and _57337_ (_05835_, _04406_, _04634_);
  and _57338_ (_05836_, _04875_, _05005_);
  and _57339_ (_05837_, _05836_, _05835_);
  and _57340_ (_05838_, _05837_, _05834_);
  and _57341_ (_05839_, _05838_, _05363_);
  or _57342_ (_05840_, _05839_, _05833_);
  nand _57343_ (_05841_, _05839_, _05833_);
  and _57344_ (_05842_, _05841_, _05840_);
  and _57345_ (_05843_, _03595_, _03197_);
  nor _57346_ (_05844_, _04322_, _05843_);
  and _57347_ (_05845_, _04474_, _03197_);
  not _57348_ (_05846_, _05845_);
  and _57349_ (_05847_, _05846_, _05844_);
  and _57350_ (_05848_, _05847_, _04745_);
  or _57351_ (_05849_, _05848_, _05842_);
  not _57352_ (_05850_, _04511_);
  and _57353_ (_05851_, _03654_, _01716_);
  and _57354_ (_05852_, _03657_, _01688_);
  nor _57355_ (_05853_, _05852_, _05851_);
  and _57356_ (_05854_, _03685_, _01719_);
  and _57357_ (_05855_, _03698_, _01673_);
  nor _57358_ (_05856_, _05855_, _05854_);
  and _57359_ (_05857_, _05856_, _05853_);
  and _57360_ (_05858_, _03701_, _01663_);
  and _57361_ (_05859_, _03703_, _01632_);
  nor _57362_ (_05860_, _05859_, _05858_);
  and _57363_ (_05861_, _03672_, _01697_);
  and _57364_ (_05862_, _03678_, _01735_);
  nor _57365_ (_05863_, _05862_, _05861_);
  and _57366_ (_05864_, _05863_, _05860_);
  and _57367_ (_05865_, _05864_, _05857_);
  and _57368_ (_05866_, _03662_, _01708_);
  and _57369_ (_05867_, _03692_, _01723_);
  nor _57370_ (_05868_, _05867_, _05866_);
  and _57371_ (_05869_, _03687_, _01731_);
  and _57372_ (_05870_, _03690_, _01704_);
  nor _57373_ (_05871_, _05870_, _05869_);
  and _57374_ (_05872_, _05871_, _05868_);
  and _57375_ (_05873_, _03675_, _01713_);
  and _57376_ (_05874_, _03680_, _01668_);
  nor _57377_ (_05875_, _05874_, _05873_);
  and _57378_ (_05876_, _03696_, _01678_);
  and _57379_ (_05877_, _03665_, _01684_);
  nor _57380_ (_05878_, _05877_, _05876_);
  and _57381_ (_05879_, _05878_, _05875_);
  and _57382_ (_05880_, _05879_, _05872_);
  and _57383_ (_05881_, _05880_, _05865_);
  and _57384_ (_05882_, _05881_, _05309_);
  nor _57385_ (_05883_, _05881_, _05309_);
  nor _57386_ (_05884_, _05883_, _05882_);
  and _57387_ (_05885_, _05884_, _04512_);
  not _57388_ (_05886_, _03601_);
  not _57389_ (_05887_, _04754_);
  not _57390_ (_05888_, _04502_);
  nor _57391_ (_05889_, _04717_, _04714_);
  and _57392_ (_05890_, _03494_, _03176_);
  nor _57393_ (_05891_, _05890_, _04493_);
  and _57394_ (_05892_, _05891_, _05889_);
  and _57395_ (_05893_, _05892_, _05888_);
  and _57396_ (_05894_, _05893_, _05887_);
  and _57397_ (_05895_, _05894_, _05886_);
  or _57398_ (_05896_, _05895_, _03454_);
  not _57399_ (_05897_, _03224_);
  nor _57400_ (_05898_, _03487_, _04051_);
  and _57401_ (_05899_, _03864_, _03583_);
  and _57402_ (_05900_, _05899_, _05898_);
  and _57403_ (_05901_, _05244_, _05900_);
  and _57404_ (_05902_, _05901_, \oc8051_golden_model_1.PSW [7]);
  and _57405_ (_05903_, _05253_, _05900_);
  and _57406_ (_05904_, _05903_, \oc8051_golden_model_1.ACC [7]);
  nor _57407_ (_05905_, _05904_, _05902_);
  nor _57408_ (_05906_, _03861_, _03583_);
  and _57409_ (_05907_, _05906_, _05898_);
  and _57410_ (_05908_, _05907_, _05238_);
  and _57411_ (_05909_, _05908_, \oc8051_golden_model_1.IP [7]);
  and _57412_ (_05910_, _05247_, _05900_);
  and _57413_ (_05911_, _05910_, \oc8051_golden_model_1.B [7]);
  nor _57414_ (_05912_, _05911_, _05909_);
  and _57415_ (_05913_, _05912_, _05905_);
  and _57416_ (_05914_, _05209_, \oc8051_golden_model_1.P0INREG [7]);
  not _57417_ (_05915_, _05914_);
  and _57418_ (_05916_, _05220_, _05900_);
  and _57419_ (_05917_, _05916_, \oc8051_golden_model_1.P1INREG [7]);
  and _57420_ (_05918_, _05228_, _05900_);
  and _57421_ (_05919_, _05918_, \oc8051_golden_model_1.P2INREG [7]);
  nor _57422_ (_05920_, _05919_, _05917_);
  and _57423_ (_05921_, _05920_, _05915_);
  and _57424_ (_05922_, _05907_, _05220_);
  and _57425_ (_05923_, _05922_, \oc8051_golden_model_1.SCON [7]);
  and _57426_ (_05924_, _05907_, _05228_);
  and _57427_ (_05925_, _05924_, \oc8051_golden_model_1.IE [7]);
  nor _57428_ (_05926_, _05925_, _05923_);
  and _57429_ (_05927_, _05907_, _05208_);
  and _57430_ (_05928_, _05927_, \oc8051_golden_model_1.TCON [7]);
  and _57431_ (_05929_, _05238_, _05900_);
  and _57432_ (_05930_, _05929_, \oc8051_golden_model_1.P3INREG [7]);
  nor _57433_ (_05931_, _05930_, _05928_);
  and _57434_ (_05932_, _05931_, _05926_);
  and _57435_ (_05933_, _05932_, _05921_);
  and _57436_ (_05934_, _05933_, _05913_);
  and _57437_ (_05935_, _05934_, _05205_);
  nor _57438_ (_05936_, _05935_, _05211_);
  and _57439_ (_05937_, _05211_, \oc8051_golden_model_1.PSW [7]);
  nor _57440_ (_05938_, _05937_, _05936_);
  nor _57441_ (_05939_, _05938_, _05063_);
  not _57442_ (_05940_, _04449_);
  and _57443_ (_05941_, _05918_, \oc8051_golden_model_1.P2 [7]);
  and _57444_ (_05942_, _05929_, \oc8051_golden_model_1.P3 [7]);
  or _57445_ (_05943_, _05942_, _05941_);
  nor _57446_ (_05944_, _05943_, _05928_);
  and _57447_ (_05945_, _05209_, \oc8051_golden_model_1.P0 [7]);
  and _57448_ (_05946_, _05916_, \oc8051_golden_model_1.P1 [7]);
  nor _57449_ (_05947_, _05946_, _05945_);
  and _57450_ (_05948_, _05947_, _05926_);
  and _57451_ (_05949_, _05948_, _05913_);
  and _57452_ (_05950_, _05949_, _05944_);
  and _57453_ (_05951_, _05950_, _05205_);
  nor _57454_ (_05952_, _05951_, _05211_);
  or _57455_ (_05953_, _05952_, _05940_);
  not _57456_ (_05954_, _04428_);
  and _57457_ (_05955_, _05824_, _05517_);
  not _57458_ (_05956_, _05666_);
  and _57459_ (_05957_, _05956_, _05617_);
  and _57460_ (_05958_, _05717_, _05566_);
  and _57461_ (_05959_, _05958_, _05957_);
  and _57462_ (_05960_, _05959_, _05955_);
  and _57463_ (_05961_, _05960_, _05411_);
  nor _57464_ (_05962_, _05961_, _05310_);
  and _57465_ (_05963_, _05961_, _05310_);
  nor _57466_ (_05964_, _05963_, _05962_);
  and _57467_ (_05965_, _05964_, _04421_);
  not _57468_ (_05966_, _04422_);
  nor _57469_ (_05967_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _57470_ (_05968_, _05967_, _03995_);
  nor _57471_ (_05969_, _05968_, _03722_);
  nor _57472_ (_05970_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _57473_ (_05971_, _05970_, _03722_);
  and _57474_ (_05972_, _05971_, _03498_);
  nor _57475_ (_05973_, _05972_, _05969_);
  nor _57476_ (_05974_, _05973_, _03997_);
  not _57477_ (_05975_, _05974_);
  not _57478_ (_05976_, _04463_);
  nand _57479_ (_05977_, _05005_, _05976_);
  and _57480_ (_05978_, _04463_, _03581_);
  not _57481_ (_05979_, _05978_);
  and _57482_ (_05980_, _05979_, _03997_);
  nand _57483_ (_05981_, _05980_, _05977_);
  and _57484_ (_05982_, _05981_, _05975_);
  nor _57485_ (_05983_, _05967_, _03995_);
  nor _57486_ (_05984_, _05983_, _05968_);
  nor _57487_ (_05985_, _05984_, _03997_);
  not _57488_ (_05986_, _05985_);
  nand _57489_ (_05987_, _04875_, _05976_);
  and _57490_ (_05988_, _04463_, _03904_);
  not _57491_ (_05989_, _05988_);
  and _57492_ (_05990_, _05989_, _03997_);
  nand _57493_ (_05991_, _05990_, _05987_);
  and _57494_ (_05992_, _05991_, _05986_);
  or _57495_ (_05993_, _04463_, _04620_);
  not _57496_ (_05994_, _03997_);
  and _57497_ (_05995_, _04463_, _04048_);
  nor _57498_ (_05997_, _05995_, _05994_);
  nand _57499_ (_05998_, _05997_, _05993_);
  nor _57500_ (_06000_, _03997_, \oc8051_golden_model_1.SP [0]);
  not _57501_ (_06001_, _06000_);
  nand _57502_ (_06003_, _06001_, _05998_);
  or _57503_ (_06004_, _06003_, _05144_);
  nor _57504_ (_06006_, _03500_, _03997_);
  not _57505_ (_06007_, _06006_);
  or _57506_ (_06009_, _04406_, _04463_);
  or _57507_ (_06010_, _05976_, _03414_);
  and _57508_ (_06012_, _06010_, _03997_);
  nand _57509_ (_06013_, _06012_, _06009_);
  and _57510_ (_06015_, _06013_, _06007_);
  not _57511_ (_06016_, _06015_);
  and _57512_ (_06018_, _06001_, _05998_);
  or _57513_ (_06019_, _06018_, _05146_);
  and _57514_ (_06021_, _06019_, _06016_);
  nand _57515_ (_06022_, _06021_, _06004_);
  or _57516_ (_06024_, _06003_, _05152_);
  or _57517_ (_06025_, _06018_, _05150_);
  and _57518_ (_06027_, _06025_, _06015_);
  nand _57519_ (_06028_, _06027_, _06024_);
  nand _57520_ (_06030_, _06028_, _06022_);
  nand _57521_ (_06031_, _06030_, _05992_);
  not _57522_ (_06033_, _05992_);
  or _57523_ (_06034_, _06003_, _05164_);
  or _57524_ (_06035_, _06018_, _05166_);
  and _57525_ (_06036_, _06035_, _06016_);
  nand _57526_ (_06037_, _06036_, _06034_);
  or _57527_ (_06038_, _06003_, _05160_);
  or _57528_ (_06039_, _06018_, _05158_);
  and _57529_ (_06040_, _06039_, _06015_);
  nand _57530_ (_06041_, _06040_, _06038_);
  nand _57531_ (_06042_, _06041_, _06037_);
  nand _57532_ (_06043_, _06042_, _06033_);
  nand _57533_ (_06044_, _06043_, _06031_);
  nand _57534_ (_06045_, _06044_, _05982_);
  not _57535_ (_06046_, _05982_);
  or _57536_ (_06047_, _06003_, _05176_);
  or _57537_ (_06048_, _06018_, _05174_);
  and _57538_ (_06049_, _06048_, _06015_);
  nand _57539_ (_06050_, _06049_, _06047_);
  or _57540_ (_06051_, _06003_, _05180_);
  or _57541_ (_06052_, _06018_, _05182_);
  and _57542_ (_06053_, _06052_, _06016_);
  nand _57543_ (_06054_, _06053_, _06051_);
  nand _57544_ (_06055_, _06054_, _06050_);
  nand _57545_ (_06056_, _06055_, _05992_);
  or _57546_ (_06057_, _06003_, _05194_);
  or _57547_ (_06058_, _06018_, _05196_);
  and _57548_ (_06059_, _06058_, _06016_);
  nand _57549_ (_06060_, _06059_, _06057_);
  or _57550_ (_06061_, _06003_, _05190_);
  or _57551_ (_06062_, _06018_, _05188_);
  and _57552_ (_06063_, _06062_, _06015_);
  nand _57553_ (_06064_, _06063_, _06061_);
  nand _57554_ (_06065_, _06064_, _06060_);
  nand _57555_ (_06066_, _06065_, _06033_);
  nand _57556_ (_06067_, _06066_, _06056_);
  nand _57557_ (_06068_, _06067_, _06046_);
  and _57558_ (_06069_, _06068_, _06045_);
  or _57559_ (_06070_, _06069_, _05966_);
  not _57560_ (_06071_, _04421_);
  or _57561_ (_06072_, _03229_, _03219_);
  not _57562_ (_06073_, _06072_);
  and _57563_ (_06074_, _06073_, _05842_);
  not _57564_ (_06075_, \oc8051_golden_model_1.ACC [7]);
  nor _57565_ (_06076_, _03980_, _06075_);
  and _57566_ (_06077_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and _57567_ (_06078_, _06077_, \oc8051_golden_model_1.PC [6]);
  and _57568_ (_06079_, _06078_, _03295_);
  and _57569_ (_06080_, _06079_, \oc8051_golden_model_1.PC [7]);
  nor _57570_ (_06081_, _06079_, \oc8051_golden_model_1.PC [7]);
  nor _57571_ (_06082_, _06081_, _06080_);
  and _57572_ (_06083_, _06082_, _03980_);
  or _57573_ (_06084_, _06083_, _06076_);
  and _57574_ (_06085_, _06084_, _06072_);
  or _57575_ (_06086_, _06085_, _04422_);
  or _57576_ (_06087_, _06086_, _06074_);
  and _57577_ (_06088_, _06087_, _06071_);
  and _57578_ (_06089_, _06088_, _06070_);
  or _57579_ (_06090_, _06089_, _05965_);
  and _57580_ (_06092_, _06090_, _05954_);
  not _57581_ (_06094_, _05211_);
  nand _57582_ (_06095_, _05951_, _06094_);
  and _57583_ (_06097_, _06095_, _04428_);
  or _57584_ (_06098_, _06097_, _04768_);
  or _57585_ (_06100_, _06098_, _06092_);
  nor _57586_ (_06101_, _06082_, _03230_);
  nor _57587_ (_06103_, _06101_, _04431_);
  and _57588_ (_06104_, _06103_, _06100_);
  and _57589_ (_06106_, _05833_, _04431_);
  or _57590_ (_06107_, _06106_, _04449_);
  or _57591_ (_06109_, _06107_, _06104_);
  and _57592_ (_06110_, _06109_, _05953_);
  or _57593_ (_06112_, _06110_, _03508_);
  not _57594_ (_06113_, _05259_);
  nor _57595_ (_06115_, _05272_, _05264_);
  and _57596_ (_06116_, _06115_, _05288_);
  and _57597_ (_06118_, _06116_, _06113_);
  and _57598_ (_06119_, _06118_, _05306_);
  and _57599_ (_06121_, _05280_, _05232_);
  and _57600_ (_06122_, _05235_, \oc8051_golden_model_1.P2INREG [7]);
  and _57601_ (_06124_, _05239_, \oc8051_golden_model_1.P3INREG [7]);
  nor _57602_ (_06125_, _06124_, _06122_);
  and _57603_ (_06126_, _05266_, \oc8051_golden_model_1.P1INREG [7]);
  and _57604_ (_06127_, _05293_, \oc8051_golden_model_1.P0INREG [7]);
  nor _57605_ (_06128_, _06127_, _06126_);
  and _57606_ (_06129_, _06128_, _06125_);
  and _57607_ (_06130_, _06129_, _05257_);
  and _57608_ (_06131_, _06130_, _06121_);
  and _57609_ (_06132_, _06131_, _06119_);
  and _57610_ (_06133_, _06132_, _05205_);
  nand _57611_ (_06134_, _06133_, _03508_);
  and _57612_ (_06135_, _06134_, _04562_);
  and _57613_ (_06136_, _06135_, _06112_);
  nor _57614_ (_06137_, _05951_, _06094_);
  not _57615_ (_06138_, _06137_);
  and _57616_ (_06139_, _06138_, _06095_);
  and _57617_ (_06140_, _06139_, _04454_);
  or _57618_ (_06141_, _06140_, _06136_);
  and _57619_ (_06142_, _06141_, _03227_);
  not _57620_ (_06143_, _06082_);
  nor _57621_ (_06144_, _06143_, _03227_);
  or _57622_ (_06145_, _06144_, _03745_);
  or _57623_ (_06146_, _06145_, _06142_);
  nand _57624_ (_06147_, _06133_, _03745_);
  and _57625_ (_06148_, _06147_, _06146_);
  or _57626_ (_06149_, _06148_, _04463_);
  and _57627_ (_06150_, _06069_, _03446_);
  nand _57628_ (_06151_, _06132_, _04463_);
  or _57629_ (_06152_, _06151_, _06150_);
  and _57630_ (_06153_, _06152_, _05063_);
  and _57631_ (_06154_, _06153_, _06149_);
  or _57632_ (_06155_, _06154_, _05939_);
  and _57633_ (_06156_, _06155_, _05897_);
  nand _57634_ (_06157_, _06082_, _03224_);
  nand _57635_ (_06158_, _06157_, _04480_);
  or _57636_ (_06159_, _06158_, _06156_);
  or _57637_ (_06160_, _05833_, _04480_);
  and _57638_ (_06161_, _06160_, _06159_);
  or _57639_ (_06162_, _06161_, _04482_);
  not _57640_ (_06163_, _04483_);
  not _57641_ (_06164_, _04482_);
  or _57642_ (_06165_, _06069_, _06164_);
  and _57643_ (_06166_, _06165_, _06163_);
  and _57644_ (_06167_, _06166_, _06162_);
  not _57645_ (_06168_, _05894_);
  and _57646_ (_06169_, _03446_, _03222_);
  not _57647_ (_06170_, _06169_);
  not _57648_ (_06171_, _05881_);
  nor _57649_ (_06172_, _06171_, _05204_);
  and _57650_ (_06173_, _03946_, _03708_);
  and _57651_ (_06174_, _03654_, _02224_);
  and _57652_ (_06175_, _03657_, _02202_);
  nor _57653_ (_06176_, _06175_, _06174_);
  and _57654_ (_06177_, _03687_, _02221_);
  and _57655_ (_06178_, _03698_, _02196_);
  nor _57656_ (_06179_, _06178_, _06177_);
  and _57657_ (_06180_, _06179_, _06176_);
  and _57658_ (_06181_, _03701_, _02187_);
  and _57659_ (_06182_, _03703_, _02190_);
  nor _57660_ (_06183_, _06182_, _06181_);
  and _57661_ (_06184_, _03675_, _02213_);
  and _57662_ (_06185_, _03678_, _02217_);
  nor _57663_ (_06186_, _06185_, _06184_);
  and _57664_ (_06187_, _06186_, _06183_);
  and _57665_ (_06188_, _06187_, _06180_);
  and _57666_ (_06189_, _03690_, _02233_);
  and _57667_ (_06190_, _03692_, _02228_);
  nor _57668_ (_06191_, _06190_, _06189_);
  and _57669_ (_06192_, _03685_, _02226_);
  and _57670_ (_06193_, _03662_, _02235_);
  nor _57671_ (_06194_, _06193_, _06192_);
  and _57672_ (_06195_, _06194_, _06191_);
  and _57673_ (_06196_, _03672_, _02210_);
  and _57674_ (_06197_, _03680_, _02185_);
  nor _57675_ (_06198_, _06197_, _06196_);
  and _57676_ (_06199_, _03696_, _02193_);
  and _57677_ (_06200_, _03665_, _02200_);
  nor _57678_ (_06201_, _06200_, _06199_);
  and _57679_ (_06202_, _06201_, _06198_);
  and _57680_ (_06203_, _06202_, _06195_);
  and _57681_ (_06204_, _06203_, _06188_);
  and _57682_ (_06205_, _06204_, _06171_);
  and _57683_ (_06206_, _03685_, _02114_);
  and _57684_ (_06207_, _03703_, _02080_);
  nor _57685_ (_06208_, _06207_, _06206_);
  and _57686_ (_06209_, _03692_, _02117_);
  and _57687_ (_06210_, _03680_, _02075_);
  nor _57688_ (_06211_, _06210_, _06209_);
  and _57689_ (_06212_, _06211_, _06208_);
  and _57690_ (_06213_, _03665_, _02090_);
  and _57691_ (_06214_, _03701_, _02077_);
  nor _57692_ (_06215_, _06214_, _06213_);
  and _57693_ (_06216_, _03654_, _02087_);
  and _57694_ (_06217_, _03678_, _02125_);
  nor _57695_ (_06218_, _06217_, _06216_);
  and _57696_ (_06219_, _06218_, _06215_);
  and _57697_ (_06220_, _06219_, _06212_);
  and _57698_ (_06221_, _03675_, _02101_);
  and _57699_ (_06222_, _03657_, _02112_);
  nor _57700_ (_06223_, _06222_, _06221_);
  and _57701_ (_06224_, _03687_, _02098_);
  and _57702_ (_06225_, _03696_, _02084_);
  nor _57703_ (_06226_, _06225_, _06224_);
  and _57704_ (_06227_, _06226_, _06223_);
  and _57705_ (_06228_, _03690_, _02104_);
  and _57706_ (_06229_, _03698_, _02082_);
  nor _57707_ (_06230_, _06229_, _06228_);
  and _57708_ (_06231_, _03662_, _02109_);
  and _57709_ (_06232_, _03672_, _02123_);
  nor _57710_ (_06233_, _06232_, _06231_);
  and _57711_ (_06234_, _06233_, _06230_);
  and _57712_ (_06235_, _06234_, _06227_);
  and _57713_ (_06236_, _06235_, _06220_);
  and _57714_ (_06237_, _03685_, _02170_);
  and _57715_ (_06238_, _03657_, _02139_);
  nor _57716_ (_06239_, _06238_, _06237_);
  and _57717_ (_06240_, _03687_, _02154_);
  and _57718_ (_06241_, _03698_, _02144_);
  nor _57719_ (_06242_, _06241_, _06240_);
  and _57720_ (_06243_, _06242_, _06239_);
  and _57721_ (_06244_, _03675_, _02178_);
  and _57722_ (_06245_, _03672_, _02160_);
  nor _57723_ (_06246_, _06245_, _06244_);
  and _57724_ (_06247_, _03692_, _02173_);
  and _57725_ (_06248_, _03654_, _02146_);
  nor _57726_ (_06249_, _06248_, _06247_);
  and _57727_ (_06250_, _06249_, _06246_);
  and _57728_ (_06251_, _06250_, _06243_);
  and _57729_ (_06252_, _03690_, _02165_);
  and _57730_ (_06253_, _03662_, _02157_);
  nor _57731_ (_06254_, _06253_, _06252_);
  and _57732_ (_06255_, _03665_, _02168_);
  and _57733_ (_06256_, _03701_, _02132_);
  nor _57734_ (_06257_, _06256_, _06255_);
  and _57735_ (_06258_, _06257_, _06254_);
  and _57736_ (_06259_, _03696_, _02137_);
  and _57737_ (_06260_, _03678_, _02180_);
  nor _57738_ (_06261_, _06260_, _06259_);
  and _57739_ (_06262_, _03680_, _02135_);
  and _57740_ (_06263_, _03703_, _02130_);
  nor _57741_ (_06264_, _06263_, _06262_);
  and _57742_ (_06265_, _06264_, _06261_);
  and _57743_ (_06266_, _06265_, _06258_);
  and _57744_ (_06267_, _06266_, _06251_);
  and _57745_ (_06268_, _06267_, _06236_);
  and _57746_ (_06269_, _06268_, _06205_);
  nor _57747_ (_06270_, _04303_, _04163_);
  and _57748_ (_06271_, _06270_, _06269_);
  and _57749_ (_06272_, _06271_, _06173_);
  and _57750_ (_06273_, _06272_, \oc8051_golden_model_1.DPH [7]);
  not _57751_ (_06274_, _04163_);
  and _57752_ (_06275_, _04303_, _06274_);
  not _57753_ (_06276_, _03708_);
  and _57754_ (_06277_, _03946_, _06276_);
  and _57755_ (_06278_, _06277_, _06269_);
  and _57756_ (_06279_, _06278_, _06275_);
  and _57757_ (_06280_, _06279_, \oc8051_golden_model_1.TMOD [7]);
  nor _57758_ (_06281_, _06280_, _06273_);
  not _57759_ (_06282_, _04303_);
  and _57760_ (_06283_, _06282_, _04163_);
  and _57761_ (_06284_, _06283_, _06278_);
  and _57762_ (_06285_, _06284_, \oc8051_golden_model_1.TL0 [7]);
  nor _57763_ (_06286_, _03946_, _03708_);
  and _57764_ (_06287_, _06286_, _06269_);
  and _57765_ (_06288_, _06287_, _06275_);
  and _57766_ (_06289_, _06288_, \oc8051_golden_model_1.TH1 [7]);
  nor _57767_ (_06290_, _06289_, _06285_);
  and _57768_ (_06291_, _06290_, _06281_);
  and _57769_ (_06292_, _04303_, _04163_);
  and _57770_ (_06293_, _06292_, _06277_);
  nor _57771_ (_06294_, _06267_, _06236_);
  and _57772_ (_06295_, _06294_, _06205_);
  and _57773_ (_06296_, _06295_, _06293_);
  and _57774_ (_06297_, _06296_, \oc8051_golden_model_1.IP [7]);
  not _57775_ (_06298_, _06236_);
  and _57776_ (_06299_, _06267_, _06298_);
  and _57777_ (_06300_, _06292_, _06173_);
  nor _57778_ (_06301_, _06204_, _05881_);
  and _57779_ (_06302_, _06301_, _06300_);
  and _57780_ (_06303_, _06302_, _06299_);
  and _57781_ (_06304_, _06303_, \oc8051_golden_model_1.PSW [7]);
  nor _57782_ (_06305_, _06304_, _06297_);
  not _57783_ (_06306_, _06267_);
  and _57784_ (_06307_, _06306_, _06236_);
  and _57785_ (_06308_, _06307_, _06302_);
  and _57786_ (_06309_, _06308_, \oc8051_golden_model_1.ACC [7]);
  and _57787_ (_06310_, _06302_, _06294_);
  and _57788_ (_06311_, _06310_, \oc8051_golden_model_1.B [7]);
  nor _57789_ (_06312_, _06311_, _06309_);
  and _57790_ (_06313_, _06312_, _06305_);
  and _57791_ (_06314_, _06307_, _06205_);
  and _57792_ (_06315_, _06314_, _06293_);
  and _57793_ (_06316_, _06315_, \oc8051_golden_model_1.IE [7]);
  and _57794_ (_06317_, _06299_, _06205_);
  and _57795_ (_06318_, _06277_, _06275_);
  and _57796_ (_06319_, _06318_, _06317_);
  and _57797_ (_06320_, _06319_, \oc8051_golden_model_1.SBUF [7]);
  and _57798_ (_06321_, _06317_, _06293_);
  and _57799_ (_06322_, _06321_, \oc8051_golden_model_1.SCON [7]);
  or _57800_ (_06323_, _06322_, _06320_);
  nor _57801_ (_06324_, _06323_, _06316_);
  and _57802_ (_06325_, _06324_, _06313_);
  and _57803_ (_06326_, _06325_, _06291_);
  and _57804_ (_06327_, _06292_, _06287_);
  and _57805_ (_06328_, _06327_, \oc8051_golden_model_1.TH0 [7]);
  and _57806_ (_06329_, _06277_, _06271_);
  and _57807_ (_06330_, _06329_, \oc8051_golden_model_1.TL1 [7]);
  nor _57808_ (_06331_, _06330_, _06328_);
  not _57809_ (_06332_, _03946_);
  and _57810_ (_06333_, _06332_, _03708_);
  and _57811_ (_06334_, _06333_, _06271_);
  and _57812_ (_06335_, _06334_, \oc8051_golden_model_1.PCON [7]);
  and _57813_ (_06336_, _06292_, _06278_);
  and _57814_ (_06337_, _06336_, \oc8051_golden_model_1.TCON [7]);
  nor _57815_ (_06338_, _06337_, _06335_);
  and _57816_ (_06339_, _06338_, _06331_);
  and _57817_ (_06340_, _06317_, _06300_);
  and _57818_ (_06341_, _06340_, \oc8051_golden_model_1.P1INREG [7]);
  not _57819_ (_06342_, _06341_);
  and _57820_ (_06343_, _06300_, _06269_);
  and _57821_ (_06344_, _06343_, \oc8051_golden_model_1.P0INREG [7]);
  not _57822_ (_06345_, _06344_);
  and _57823_ (_06346_, _06314_, _06300_);
  and _57824_ (_06347_, _06346_, \oc8051_golden_model_1.P2INREG [7]);
  and _57825_ (_06348_, _06300_, _06295_);
  and _57826_ (_06349_, _06348_, \oc8051_golden_model_1.P3INREG [7]);
  nor _57827_ (_06350_, _06349_, _06347_);
  and _57828_ (_06351_, _06350_, _06345_);
  and _57829_ (_06352_, _06351_, _06342_);
  and _57830_ (_06353_, _06269_, _06173_);
  and _57831_ (_06354_, _06353_, _06275_);
  and _57832_ (_06355_, _06354_, \oc8051_golden_model_1.SP [7]);
  and _57833_ (_06356_, _06353_, _06283_);
  and _57834_ (_06357_, _06356_, \oc8051_golden_model_1.DPL [7]);
  nor _57835_ (_06358_, _06357_, _06355_);
  and _57836_ (_06359_, _06358_, _06352_);
  and _57837_ (_06360_, _06359_, _06339_);
  and _57838_ (_06361_, _06360_, _06326_);
  not _57839_ (_06362_, _06361_);
  nor _57840_ (_06363_, _06362_, _06172_);
  nor _57841_ (_06364_, _06363_, _06170_);
  or _57842_ (_06365_, _06364_, _06168_);
  or _57843_ (_06366_, _06365_, _06167_);
  and _57844_ (_06367_, _06366_, _05896_);
  and _57845_ (_06368_, _06171_, _04500_);
  or _57846_ (_06369_, _06368_, _03178_);
  or _57847_ (_06370_, _06369_, _06367_);
  and _57848_ (_06371_, _06143_, _03178_);
  nor _57849_ (_06372_, _06371_, _04512_);
  and _57850_ (_06373_, _06372_, _06370_);
  or _57851_ (_06374_, _06373_, _05885_);
  and _57852_ (_06375_, _06374_, _05850_);
  nor _57853_ (_06376_, _05309_, _06075_);
  and _57854_ (_06377_, _05309_, _06075_);
  nor _57855_ (_06378_, _06377_, _06376_);
  and _57856_ (_06379_, _06378_, _04511_);
  or _57857_ (_06380_, _06379_, _04515_);
  or _57858_ (_06381_, _06380_, _06375_);
  not _57859_ (_06382_, _04514_);
  not _57860_ (_06383_, _04515_);
  or _57861_ (_06384_, _05883_, _06383_);
  and _57862_ (_06385_, _06384_, _06382_);
  and _57863_ (_06386_, _06385_, _06381_);
  and _57864_ (_06387_, _06376_, _04514_);
  or _57865_ (_06388_, _06387_, _03192_);
  or _57866_ (_06389_, _06388_, _06386_);
  and _57867_ (_06390_, _03624_, _03446_);
  and _57868_ (_06391_, _06143_, _03192_);
  nor _57869_ (_06392_, _06391_, _06390_);
  and _57870_ (_06393_, _06392_, _06389_);
  and _57871_ (_06394_, _03785_, _03446_);
  not _57872_ (_06395_, _06390_);
  nor _57873_ (_06396_, _05882_, _06395_);
  or _57874_ (_06397_, _06396_, _06394_);
  or _57875_ (_06398_, _06397_, _06393_);
  not _57876_ (_06399_, _03188_);
  nand _57877_ (_06400_, _06377_, _06394_);
  and _57878_ (_06401_, _06400_, _06399_);
  and _57879_ (_06402_, _06401_, _06398_);
  nand _57880_ (_06403_, _06082_, _03188_);
  nand _57881_ (_06404_, _06403_, _05848_);
  or _57882_ (_06405_, _06404_, _06402_);
  and _57883_ (_06406_, _06405_, _05849_);
  or _57884_ (_06407_, _06406_, _04533_);
  not _57885_ (_06408_, _04531_);
  not _57886_ (_06409_, _04533_);
  not _57887_ (_06410_, _06069_);
  or _57888_ (_06411_, _06003_, _05311_);
  or _57889_ (_06412_, _06018_, _05313_);
  and _57890_ (_06413_, _06412_, _06016_);
  nand _57891_ (_06414_, _06413_, _06411_);
  or _57892_ (_06415_, _06003_, _05319_);
  or _57893_ (_06416_, _06018_, _05317_);
  and _57894_ (_06417_, _06416_, _06015_);
  nand _57895_ (_06418_, _06417_, _06415_);
  nand _57896_ (_06419_, _06418_, _06414_);
  nand _57897_ (_06420_, _06419_, _05992_);
  or _57898_ (_06421_, _06003_, _05331_);
  or _57899_ (_06422_, _06018_, _05333_);
  and _57900_ (_06423_, _06422_, _06016_);
  nand _57901_ (_06424_, _06423_, _06421_);
  or _57902_ (_06425_, _06003_, _05327_);
  or _57903_ (_06426_, _06018_, _05325_);
  and _57904_ (_06427_, _06426_, _06015_);
  nand _57905_ (_06428_, _06427_, _06425_);
  nand _57906_ (_06429_, _06428_, _06424_);
  nand _57907_ (_06430_, _06429_, _06033_);
  and _57908_ (_06431_, _06430_, _05982_);
  and _57909_ (_06432_, _06431_, _06420_);
  or _57910_ (_06433_, _06003_, \oc8051_golden_model_1.IRAM[10] [6]);
  or _57911_ (_06434_, _06018_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _57912_ (_06435_, _06434_, _06433_);
  nand _57913_ (_06436_, _06435_, _06015_);
  or _57914_ (_06437_, _06003_, \oc8051_golden_model_1.IRAM[8] [6]);
  or _57915_ (_06438_, _06018_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand _57916_ (_06439_, _06438_, _06437_);
  nand _57917_ (_06440_, _06439_, _06016_);
  nand _57918_ (_06441_, _06440_, _06436_);
  nand _57919_ (_06442_, _06441_, _05992_);
  or _57920_ (_06443_, _06003_, \oc8051_golden_model_1.IRAM[14] [6]);
  or _57921_ (_06444_, _06018_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _57922_ (_06445_, _06444_, _06443_);
  nand _57923_ (_06446_, _06445_, _06015_);
  or _57924_ (_06447_, _06003_, \oc8051_golden_model_1.IRAM[12] [6]);
  or _57925_ (_06448_, _06018_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand _57926_ (_06449_, _06448_, _06447_);
  nand _57927_ (_06450_, _06449_, _06016_);
  nand _57928_ (_06451_, _06450_, _06446_);
  nand _57929_ (_06452_, _06451_, _06033_);
  and _57930_ (_06453_, _06452_, _06046_);
  and _57931_ (_06454_, _06453_, _06442_);
  or _57932_ (_06455_, _06454_, _06432_);
  not _57933_ (_06456_, _06455_);
  or _57934_ (_06457_, _06003_, _04017_);
  or _57935_ (_06458_, _06018_, _04347_);
  and _57936_ (_06459_, _06458_, _06016_);
  nand _57937_ (_06460_, _06459_, _06457_);
  or _57938_ (_06461_, _06003_, _04355_);
  or _57939_ (_06462_, _06018_, _04352_);
  and _57940_ (_06463_, _06462_, _06015_);
  nand _57941_ (_06464_, _06463_, _06461_);
  nand _57942_ (_06465_, _06464_, _06460_);
  nand _57943_ (_06466_, _06465_, _05992_);
  or _57944_ (_06467_, _06003_, _04368_);
  or _57945_ (_06468_, _06018_, _04370_);
  and _57946_ (_06469_, _06468_, _06016_);
  nand _57947_ (_06470_, _06469_, _06467_);
  or _57948_ (_06471_, _06003_, _04364_);
  or _57949_ (_06472_, _06018_, _04362_);
  and _57950_ (_06473_, _06472_, _06015_);
  nand _57951_ (_06474_, _06473_, _06471_);
  nand _57952_ (_06475_, _06474_, _06470_);
  nand _57953_ (_06476_, _06475_, _06033_);
  and _57954_ (_06477_, _06476_, _05982_);
  and _57955_ (_06478_, _06477_, _06466_);
  or _57956_ (_06479_, _06003_, \oc8051_golden_model_1.IRAM[10] [1]);
  or _57957_ (_06480_, _06018_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _57958_ (_06481_, _06480_, _06479_);
  nand _57959_ (_06482_, _06481_, _06015_);
  or _57960_ (_06483_, _06003_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _57961_ (_06484_, _06018_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand _57962_ (_06485_, _06484_, _06483_);
  nand _57963_ (_06486_, _06485_, _06016_);
  nand _57964_ (_06487_, _06486_, _06482_);
  nand _57965_ (_06488_, _06487_, _05992_);
  or _57966_ (_06489_, _06003_, \oc8051_golden_model_1.IRAM[14] [1]);
  or _57967_ (_06490_, _06018_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _57968_ (_06491_, _06490_, _06489_);
  nand _57969_ (_06492_, _06491_, _06015_);
  or _57970_ (_06493_, _06003_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _57971_ (_06494_, _06018_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand _57972_ (_06495_, _06494_, _06493_);
  nand _57973_ (_06496_, _06495_, _06016_);
  nand _57974_ (_06497_, _06496_, _06492_);
  nand _57975_ (_06498_, _06497_, _06033_);
  and _57976_ (_06499_, _06498_, _06046_);
  and _57977_ (_06500_, _06499_, _06488_);
  or _57978_ (_06501_, _06500_, _06478_);
  or _57979_ (_06502_, _06003_, _04563_);
  or _57980_ (_06503_, _06018_, _04565_);
  and _57981_ (_06504_, _06503_, _06016_);
  nand _57982_ (_06505_, _06504_, _06502_);
  or _57983_ (_06506_, _06003_, _04571_);
  or _57984_ (_06507_, _06018_, _04569_);
  and _57985_ (_06508_, _06507_, _06015_);
  nand _57986_ (_06509_, _06508_, _06506_);
  nand _57987_ (_06510_, _06509_, _06505_);
  nand _57988_ (_06511_, _06510_, _05992_);
  or _57989_ (_06512_, _06003_, _04584_);
  or _57990_ (_06513_, _06018_, _04586_);
  and _57991_ (_06514_, _06513_, _06016_);
  nand _57992_ (_06515_, _06514_, _06512_);
  or _57993_ (_06516_, _06003_, _04580_);
  or _57994_ (_06517_, _06018_, _04578_);
  and _57995_ (_06518_, _06517_, _06015_);
  nand _57996_ (_06519_, _06518_, _06516_);
  nand _57997_ (_06520_, _06519_, _06515_);
  nand _57998_ (_06521_, _06520_, _06033_);
  and _57999_ (_06522_, _06521_, _05982_);
  and _58000_ (_06523_, _06522_, _06511_);
  or _58001_ (_06524_, _06003_, \oc8051_golden_model_1.IRAM[10] [0]);
  or _58002_ (_06525_, _06018_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _58003_ (_06526_, _06525_, _06524_);
  nand _58004_ (_06527_, _06526_, _06015_);
  or _58005_ (_06528_, _06003_, \oc8051_golden_model_1.IRAM[8] [0]);
  or _58006_ (_06529_, _06018_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand _58007_ (_06530_, _06529_, _06528_);
  nand _58008_ (_06531_, _06530_, _06016_);
  nand _58009_ (_06532_, _06531_, _06527_);
  nand _58010_ (_06533_, _06532_, _05992_);
  or _58011_ (_06534_, _06003_, \oc8051_golden_model_1.IRAM[14] [0]);
  or _58012_ (_06535_, _06018_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand _58013_ (_06536_, _06535_, _06534_);
  nand _58014_ (_06537_, _06536_, _06015_);
  or _58015_ (_06538_, _06003_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _58016_ (_06539_, _06018_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand _58017_ (_06540_, _06539_, _06538_);
  nand _58018_ (_06541_, _06540_, _06016_);
  nand _58019_ (_06542_, _06541_, _06537_);
  nand _58020_ (_06543_, _06542_, _06033_);
  and _58021_ (_06544_, _06543_, _06046_);
  and _58022_ (_06545_, _06544_, _06533_);
  or _58023_ (_06546_, _06545_, _06523_);
  nor _58024_ (_06547_, _06546_, _06501_);
  or _58025_ (_06548_, _06003_, _04953_);
  or _58026_ (_06549_, _06018_, _04955_);
  and _58027_ (_06550_, _06549_, _06016_);
  nand _58028_ (_06551_, _06550_, _06548_);
  or _58029_ (_06552_, _06003_, _04961_);
  or _58030_ (_06553_, _06018_, _04959_);
  and _58031_ (_06554_, _06553_, _06015_);
  nand _58032_ (_06555_, _06554_, _06552_);
  nand _58033_ (_06556_, _06555_, _06551_);
  nand _58034_ (_06557_, _06556_, _05992_);
  or _58035_ (_06558_, _06003_, _04973_);
  or _58036_ (_06559_, _06018_, _04975_);
  and _58037_ (_06560_, _06559_, _06016_);
  nand _58038_ (_06561_, _06560_, _06558_);
  or _58039_ (_06562_, _06003_, _04969_);
  or _58040_ (_06563_, _06018_, _04967_);
  and _58041_ (_06564_, _06563_, _06015_);
  nand _58042_ (_06565_, _06564_, _06562_);
  nand _58043_ (_06566_, _06565_, _06561_);
  nand _58044_ (_06567_, _06566_, _06033_);
  and _58045_ (_06568_, _06567_, _05982_);
  and _58046_ (_06569_, _06568_, _06557_);
  or _58047_ (_06570_, _06003_, \oc8051_golden_model_1.IRAM[10] [3]);
  or _58048_ (_06571_, _06018_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _58049_ (_06572_, _06571_, _06570_);
  nand _58050_ (_06573_, _06572_, _06015_);
  or _58051_ (_06574_, _06003_, \oc8051_golden_model_1.IRAM[8] [3]);
  or _58052_ (_06575_, _06018_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand _58053_ (_06576_, _06575_, _06574_);
  nand _58054_ (_06577_, _06576_, _06016_);
  nand _58055_ (_06578_, _06577_, _06573_);
  nand _58056_ (_06579_, _06578_, _05992_);
  or _58057_ (_06580_, _06003_, \oc8051_golden_model_1.IRAM[14] [3]);
  or _58058_ (_06581_, _06018_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _58059_ (_06582_, _06581_, _06580_);
  nand _58060_ (_06583_, _06582_, _06015_);
  or _58061_ (_06584_, _06003_, \oc8051_golden_model_1.IRAM[12] [3]);
  or _58062_ (_06585_, _06018_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand _58063_ (_06586_, _06585_, _06584_);
  nand _58064_ (_06587_, _06586_, _06016_);
  nand _58065_ (_06588_, _06587_, _06583_);
  nand _58066_ (_06589_, _06588_, _06033_);
  and _58067_ (_06590_, _06589_, _06046_);
  and _58068_ (_06591_, _06590_, _06579_);
  or _58069_ (_06592_, _06591_, _06569_);
  or _58070_ (_06593_, _06003_, _04819_);
  or _58071_ (_06594_, _06018_, _04821_);
  and _58072_ (_06595_, _06594_, _06016_);
  nand _58073_ (_06596_, _06595_, _06593_);
  or _58074_ (_06597_, _06003_, _04827_);
  or _58075_ (_06598_, _06018_, _04825_);
  and _58076_ (_06599_, _06598_, _06015_);
  nand _58077_ (_06600_, _06599_, _06597_);
  nand _58078_ (_06601_, _06600_, _06596_);
  nand _58079_ (_06602_, _06601_, _05992_);
  or _58080_ (_06603_, _06003_, _04839_);
  or _58081_ (_06604_, _06018_, _04841_);
  and _58082_ (_06605_, _06604_, _06016_);
  nand _58083_ (_06606_, _06605_, _06603_);
  or _58084_ (_06607_, _06003_, _04835_);
  or _58085_ (_06608_, _06018_, _04833_);
  and _58086_ (_06609_, _06608_, _06015_);
  nand _58087_ (_06610_, _06609_, _06607_);
  nand _58088_ (_06611_, _06610_, _06606_);
  nand _58089_ (_06612_, _06611_, _06033_);
  and _58090_ (_06613_, _06612_, _05982_);
  and _58091_ (_06614_, _06613_, _06602_);
  or _58092_ (_06615_, _06003_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _58093_ (_06616_, _06018_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _58094_ (_06617_, _06616_, _06615_);
  nand _58095_ (_06618_, _06617_, _06015_);
  or _58096_ (_06619_, _06003_, \oc8051_golden_model_1.IRAM[8] [2]);
  or _58097_ (_06620_, _06018_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand _58098_ (_06621_, _06620_, _06619_);
  nand _58099_ (_06622_, _06621_, _06016_);
  nand _58100_ (_06623_, _06622_, _06618_);
  nand _58101_ (_06624_, _06623_, _05992_);
  or _58102_ (_06625_, _06003_, \oc8051_golden_model_1.IRAM[14] [2]);
  or _58103_ (_06626_, _06018_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _58104_ (_06627_, _06626_, _06625_);
  nand _58105_ (_06628_, _06627_, _06015_);
  or _58106_ (_06629_, _06003_, \oc8051_golden_model_1.IRAM[12] [2]);
  or _58107_ (_06630_, _06018_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand _58108_ (_06631_, _06630_, _06629_);
  nand _58109_ (_06632_, _06631_, _06016_);
  nand _58110_ (_06633_, _06632_, _06628_);
  nand _58111_ (_06634_, _06633_, _06033_);
  and _58112_ (_06635_, _06634_, _06046_);
  and _58113_ (_06636_, _06635_, _06624_);
  or _58114_ (_06637_, _06636_, _06614_);
  nor _58115_ (_06638_, _06637_, _06592_);
  and _58116_ (_06639_, _06638_, _06547_);
  or _58117_ (_06640_, _06003_, _05413_);
  or _58118_ (_06641_, _06018_, _05415_);
  and _58119_ (_06642_, _06641_, _06016_);
  nand _58120_ (_06643_, _06642_, _06640_);
  or _58121_ (_06644_, _06003_, _05421_);
  or _58122_ (_06645_, _06018_, _05419_);
  and _58123_ (_06646_, _06645_, _06015_);
  nand _58124_ (_06647_, _06646_, _06644_);
  nand _58125_ (_06648_, _06647_, _06643_);
  nand _58126_ (_06649_, _06648_, _05992_);
  or _58127_ (_06650_, _06003_, _05433_);
  or _58128_ (_06651_, _06018_, _05435_);
  and _58129_ (_06652_, _06651_, _06016_);
  nand _58130_ (_06653_, _06652_, _06650_);
  or _58131_ (_06654_, _06003_, _05429_);
  or _58132_ (_06655_, _06018_, _05427_);
  and _58133_ (_06656_, _06655_, _06015_);
  nand _58134_ (_06657_, _06656_, _06654_);
  nand _58135_ (_06658_, _06657_, _06653_);
  nand _58136_ (_06659_, _06658_, _06033_);
  and _58137_ (_06660_, _06659_, _05982_);
  and _58138_ (_06661_, _06660_, _06649_);
  or _58139_ (_06662_, _06003_, \oc8051_golden_model_1.IRAM[10] [5]);
  or _58140_ (_06663_, _06018_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _58141_ (_06664_, _06663_, _06662_);
  nand _58142_ (_06665_, _06664_, _06015_);
  or _58143_ (_06666_, _06003_, \oc8051_golden_model_1.IRAM[8] [5]);
  or _58144_ (_06667_, _06018_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand _58145_ (_06668_, _06667_, _06666_);
  nand _58146_ (_06669_, _06668_, _06016_);
  nand _58147_ (_06670_, _06669_, _06665_);
  nand _58148_ (_06671_, _06670_, _05992_);
  or _58149_ (_06672_, _06003_, \oc8051_golden_model_1.IRAM[14] [5]);
  or _58150_ (_06673_, _06018_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _58151_ (_06674_, _06673_, _06672_);
  nand _58152_ (_06675_, _06674_, _06015_);
  or _58153_ (_06676_, _06003_, \oc8051_golden_model_1.IRAM[12] [5]);
  or _58154_ (_06677_, _06018_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand _58155_ (_06678_, _06677_, _06676_);
  nand _58156_ (_06679_, _06678_, _06016_);
  nand _58157_ (_06680_, _06679_, _06675_);
  nand _58158_ (_06681_, _06680_, _06033_);
  and _58159_ (_06682_, _06681_, _06046_);
  and _58160_ (_06683_, _06682_, _06671_);
  or _58161_ (_06684_, _06683_, _06661_);
  or _58162_ (_06685_, _06003_, _05721_);
  or _58163_ (_06686_, _06018_, _05723_);
  and _58164_ (_06687_, _06686_, _06016_);
  nand _58165_ (_06688_, _06687_, _06685_);
  or _58166_ (_06689_, _06003_, _05729_);
  or _58167_ (_06690_, _06018_, _05727_);
  and _58168_ (_06691_, _06690_, _06015_);
  nand _58169_ (_06692_, _06691_, _06689_);
  nand _58170_ (_06693_, _06692_, _06688_);
  nand _58171_ (_06694_, _06693_, _05992_);
  or _58172_ (_06696_, _06003_, _05741_);
  or _58173_ (_06697_, _06018_, _05743_);
  and _58174_ (_06698_, _06697_, _06016_);
  nand _58175_ (_06699_, _06698_, _06696_);
  or _58176_ (_06700_, _06003_, _05737_);
  or _58177_ (_06701_, _06018_, _05735_);
  and _58178_ (_06702_, _06701_, _06015_);
  nand _58179_ (_06703_, _06702_, _06700_);
  nand _58180_ (_06704_, _06703_, _06699_);
  nand _58181_ (_06705_, _06704_, _06033_);
  and _58182_ (_06706_, _06705_, _05982_);
  and _58183_ (_06707_, _06706_, _06694_);
  or _58184_ (_06708_, _06003_, \oc8051_golden_model_1.IRAM[10] [4]);
  or _58185_ (_06709_, _06018_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _58186_ (_06710_, _06709_, _06708_);
  nand _58187_ (_06711_, _06710_, _06015_);
  or _58188_ (_06712_, _06003_, \oc8051_golden_model_1.IRAM[8] [4]);
  or _58189_ (_06713_, _06018_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand _58190_ (_06714_, _06713_, _06712_);
  nand _58191_ (_06715_, _06714_, _06016_);
  nand _58192_ (_06716_, _06715_, _06711_);
  nand _58193_ (_06717_, _06716_, _05992_);
  or _58194_ (_06718_, _06003_, \oc8051_golden_model_1.IRAM[14] [4]);
  or _58195_ (_06719_, _06018_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _58196_ (_06720_, _06719_, _06718_);
  nand _58197_ (_06721_, _06720_, _06015_);
  or _58198_ (_06722_, _06003_, \oc8051_golden_model_1.IRAM[12] [4]);
  or _58199_ (_06723_, _06018_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand _58200_ (_06724_, _06723_, _06722_);
  nand _58201_ (_06725_, _06724_, _06016_);
  nand _58202_ (_06726_, _06725_, _06721_);
  nand _58203_ (_06727_, _06726_, _06033_);
  and _58204_ (_06728_, _06727_, _06046_);
  and _58205_ (_06729_, _06728_, _06717_);
  or _58206_ (_06730_, _06729_, _06707_);
  nor _58207_ (_06731_, _06730_, _06684_);
  and _58208_ (_06732_, _06731_, _06639_);
  and _58209_ (_06733_, _06732_, _06456_);
  nor _58210_ (_06734_, _06733_, _06410_);
  and _58211_ (_06735_, _06733_, _06410_);
  or _58212_ (_06736_, _06735_, _06734_);
  or _58213_ (_06737_, _06736_, _06409_);
  and _58214_ (_06738_, _06737_, _06408_);
  and _58215_ (_06739_, _06738_, _06407_);
  and _58216_ (_06740_, _05964_, _04531_);
  or _58217_ (_06741_, _06740_, _03629_);
  or _58218_ (_06742_, _06741_, _06739_);
  and _58219_ (_06743_, _02909_, \oc8051_golden_model_1.PC [2]);
  and _58220_ (_06744_, _06743_, \oc8051_golden_model_1.PC [3]);
  and _58221_ (_06745_, _06744_, _06078_);
  and _58222_ (_06746_, _06745_, \oc8051_golden_model_1.PC [7]);
  nor _58223_ (_06747_, _06745_, \oc8051_golden_model_1.PC [7]);
  nor _58224_ (_06748_, _06747_, _06746_);
  not _58225_ (_06749_, _06748_);
  nand _58226_ (_06750_, _06749_, _03629_);
  and _58227_ (_06751_, _06750_, _06742_);
  or _58228_ (_06752_, _06751_, _03198_);
  and _58229_ (_06753_, _06143_, _03198_);
  nor _58230_ (_06754_, _06753_, _04539_);
  and _58231_ (_06755_, _06754_, _06752_);
  and _58232_ (_06756_, _05936_, _04539_);
  nor _58233_ (_06757_, _04320_, _03960_);
  not _58234_ (_06758_, _06757_);
  nor _58235_ (_06759_, _06758_, _06756_);
  not _58236_ (_06760_, _06759_);
  nor _58237_ (_06761_, _06760_, _06755_);
  not _58238_ (_06762_, _05469_);
  not _58239_ (_06763_, _05777_);
  and _58240_ (_06764_, _04405_, _04378_);
  and _58241_ (_06765_, _06764_, _04620_);
  nor _58242_ (_06766_, _04875_, _05005_);
  and _58243_ (_06767_, _06766_, _06765_);
  and _58244_ (_06768_, _06767_, _06763_);
  and _58245_ (_06769_, _06768_, _06762_);
  and _58246_ (_06770_, _05363_, _05204_);
  nor _58247_ (_06771_, _05363_, _05204_);
  nor _58248_ (_06772_, _06771_, _06770_);
  and _58249_ (_06773_, _06772_, _06769_);
  nor _58250_ (_06774_, _06769_, _05204_);
  nor _58251_ (_06775_, _06774_, _06773_);
  and _58252_ (_06776_, _06775_, _06758_);
  nor _58253_ (_06777_, _06776_, _04547_);
  not _58254_ (_06778_, _06777_);
  nor _58255_ (_06779_, _06778_, _06761_);
  not _58256_ (_06780_, _04547_);
  nor _58257_ (_06781_, _06775_, _06780_);
  nor _58258_ (_06782_, _06781_, _04552_);
  not _58259_ (_06783_, _06782_);
  nor _58260_ (_06784_, _06783_, _06779_);
  not _58261_ (_06785_, _04552_);
  and _58262_ (_06786_, _06546_, _06501_);
  and _58263_ (_06787_, _06637_, _06592_);
  and _58264_ (_06788_, _06787_, _06786_);
  and _58265_ (_06789_, _06730_, _06684_);
  and _58266_ (_06790_, _06789_, _06788_);
  and _58267_ (_06791_, _06790_, _06455_);
  nor _58268_ (_06792_, _06791_, _06410_);
  and _58269_ (_06793_, _06791_, _06410_);
  or _58270_ (_06794_, _06793_, _06792_);
  nor _58271_ (_06795_, _06794_, _06785_);
  nor _58272_ (_06796_, _06795_, _03448_);
  not _58273_ (_06797_, _06796_);
  nor _58274_ (_06798_, _06797_, _06784_);
  nor _58275_ (_06799_, _06798_, _05832_);
  nor _58276_ (_06800_, _06799_, _04797_);
  or _58277_ (_06801_, _06800_, _05143_);
  and _58278_ (_06802_, _06801_, _05142_);
  not _58279_ (_06803_, \oc8051_golden_model_1.PC [15]);
  and _58280_ (_06804_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and _58281_ (_06805_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and _58282_ (_06806_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and _58283_ (_06807_, _06806_, _06805_);
  and _58284_ (_06808_, _06807_, _06080_);
  and _58285_ (_06809_, _06808_, _06804_);
  and _58286_ (_06810_, _06809_, \oc8051_golden_model_1.PC [14]);
  and _58287_ (_06811_, _06810_, _06803_);
  nor _58288_ (_06812_, _06810_, _06803_);
  or _58289_ (_06813_, _06812_, _06811_);
  not _58290_ (_06814_, _06813_);
  nor _58291_ (_06815_, _06814_, _03629_);
  and _58292_ (_06816_, _06807_, _06746_);
  and _58293_ (_06817_, _06816_, _06804_);
  and _58294_ (_06818_, _06817_, \oc8051_golden_model_1.PC [14]);
  and _58295_ (_06819_, _06818_, _06803_);
  nor _58296_ (_06820_, _06818_, _06803_);
  or _58297_ (_06821_, _06820_, _06819_);
  and _58298_ (_06822_, _06821_, _03629_);
  or _58299_ (_06823_, _06822_, _06815_);
  and _58300_ (_06824_, _06823_, _05137_);
  and _58301_ (_06825_, _06824_, _05140_);
  or _58302_ (_40565_, _06825_, _06802_);
  not _58303_ (_06826_, \oc8051_golden_model_1.B [7]);
  nor _58304_ (_06827_, _43000_, _06826_);
  not _58305_ (_06828_, _03790_);
  nor _58306_ (_06829_, _05248_, _06826_);
  not _58307_ (_06830_, _05248_);
  nor _58308_ (_06831_, _06830_, _05204_);
  or _58309_ (_06832_, _06831_, _06829_);
  and _58310_ (_06833_, _04058_, _03168_);
  not _58311_ (_06834_, _06833_);
  and _58312_ (_06835_, _04750_, _03168_);
  not _58313_ (_06836_, _06835_);
  and _58314_ (_06837_, _06836_, _04477_);
  and _58315_ (_06838_, _06837_, _06834_);
  or _58316_ (_06839_, _06838_, _06832_);
  not _58317_ (_06840_, _03719_);
  nor _58318_ (_06841_, _05910_, _06826_);
  and _58319_ (_06842_, _05952_, _05910_);
  or _58320_ (_06843_, _06842_, _06841_);
  and _58321_ (_06844_, _06843_, _03714_);
  and _58322_ (_06845_, _05964_, _05248_);
  or _58323_ (_06846_, _06845_, _06829_);
  or _58324_ (_06847_, _06846_, _04081_);
  and _58325_ (_06848_, _05248_, \oc8051_golden_model_1.ACC [7]);
  or _58326_ (_06849_, _06848_, _06829_);
  and _58327_ (_06850_, _06849_, _04409_);
  nor _58328_ (_06851_, _04409_, _06826_);
  or _58329_ (_06852_, _06851_, _03610_);
  or _58330_ (_06853_, _06852_, _06850_);
  and _58331_ (_06854_, _06853_, _04055_);
  and _58332_ (_06855_, _06854_, _06847_);
  and _58333_ (_06856_, _06095_, _05910_);
  or _58334_ (_06857_, _06856_, _06841_);
  and _58335_ (_06858_, _06857_, _03715_);
  or _58336_ (_06859_, _06858_, _03723_);
  or _58337_ (_06860_, _06859_, _06855_);
  or _58338_ (_06861_, _06832_, _03996_);
  and _58339_ (_06862_, _06861_, _06860_);
  or _58340_ (_06863_, _06862_, _03729_);
  or _58341_ (_06864_, _06849_, _03737_);
  and _58342_ (_06865_, _06864_, _03736_);
  and _58343_ (_06866_, _06865_, _06863_);
  or _58344_ (_06867_, _06866_, _06844_);
  and _58345_ (_06868_, _06867_, _06840_);
  and _58346_ (_06869_, _03603_, _03751_);
  or _58347_ (_06870_, _06841_, _06138_);
  and _58348_ (_06871_, _06870_, _03719_);
  and _58349_ (_06872_, _06871_, _06857_);
  or _58350_ (_06873_, _06872_, _06869_);
  or _58351_ (_06874_, _06873_, _06868_);
  not _58352_ (_06875_, _06869_);
  and _58353_ (_06876_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and _58354_ (_06877_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and _58355_ (_06878_, _06877_, _06876_);
  and _58356_ (_06879_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and _58357_ (_06880_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and _58358_ (_06881_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor _58359_ (_06882_, _06881_, _06880_);
  nor _58360_ (_06883_, _06882_, _06878_);
  and _58361_ (_06884_, _06883_, _06879_);
  nor _58362_ (_06885_, _06884_, _06878_);
  and _58363_ (_06886_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and _58364_ (_06887_, _06886_, _06881_);
  and _58365_ (_06888_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor _58366_ (_06889_, _06888_, _06876_);
  nor _58367_ (_06890_, _06889_, _06887_);
  not _58368_ (_06891_, _06890_);
  nor _58369_ (_06892_, _06891_, _06885_);
  and _58370_ (_06893_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and _58371_ (_06894_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and _58372_ (_06895_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and _58373_ (_06896_, _06895_, _06894_);
  nor _58374_ (_06897_, _06895_, _06894_);
  nor _58375_ (_06898_, _06897_, _06896_);
  and _58376_ (_06899_, _06898_, _06893_);
  nor _58377_ (_06900_, _06898_, _06893_);
  nor _58378_ (_06901_, _06900_, _06899_);
  and _58379_ (_06902_, _06891_, _06885_);
  nor _58380_ (_06903_, _06902_, _06892_);
  and _58381_ (_06904_, _06903_, _06901_);
  nor _58382_ (_06905_, _06904_, _06892_);
  not _58383_ (_06906_, _06881_);
  and _58384_ (_06907_, _06886_, _06906_);
  and _58385_ (_06908_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and _58386_ (_06909_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and _58387_ (_06910_, _06909_, _06894_);
  and _58388_ (_06911_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and _58389_ (_06912_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor _58390_ (_06913_, _06912_, _06911_);
  nor _58391_ (_06914_, _06913_, _06910_);
  and _58392_ (_06915_, _06914_, _06908_);
  nor _58393_ (_06916_, _06914_, _06908_);
  nor _58394_ (_06917_, _06916_, _06915_);
  and _58395_ (_06918_, _06917_, _06907_);
  nor _58396_ (_06919_, _06917_, _06907_);
  nor _58397_ (_06920_, _06919_, _06918_);
  not _58398_ (_06921_, _06920_);
  nor _58399_ (_06922_, _06921_, _06905_);
  and _58400_ (_06923_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and _58401_ (_06924_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and _58402_ (_06925_, _06924_, _06923_);
  nor _58403_ (_06926_, _06899_, _06896_);
  and _58404_ (_06927_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and _58405_ (_06928_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and _58406_ (_06929_, _06928_, _06927_);
  nor _58407_ (_06930_, _06928_, _06927_);
  nor _58408_ (_06931_, _06930_, _06929_);
  not _58409_ (_06932_, _06931_);
  nor _58410_ (_06933_, _06932_, _06926_);
  and _58411_ (_06934_, _06932_, _06926_);
  nor _58412_ (_06935_, _06934_, _06933_);
  and _58413_ (_06936_, _06935_, _06925_);
  nor _58414_ (_06937_, _06935_, _06925_);
  nor _58415_ (_06938_, _06937_, _06936_);
  and _58416_ (_06939_, _06921_, _06905_);
  nor _58417_ (_06940_, _06939_, _06922_);
  and _58418_ (_06941_, _06940_, _06938_);
  nor _58419_ (_06942_, _06941_, _06922_);
  nor _58420_ (_06943_, _06915_, _06910_);
  and _58421_ (_06944_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and _58422_ (_06945_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and _58423_ (_06946_, _06945_, _06944_);
  nor _58424_ (_06947_, _06945_, _06944_);
  nor _58425_ (_06948_, _06947_, _06946_);
  not _58426_ (_06949_, _06948_);
  nor _58427_ (_06950_, _06949_, _06943_);
  and _58428_ (_06951_, _06949_, _06943_);
  nor _58429_ (_06952_, _06951_, _06950_);
  and _58430_ (_06953_, _06952_, _06929_);
  nor _58431_ (_06954_, _06952_, _06929_);
  nor _58432_ (_06955_, _06954_, _06953_);
  nor _58433_ (_06956_, _06918_, _06887_);
  and _58434_ (_06957_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and _58435_ (_06958_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and _58436_ (_06959_, _06958_, _06909_);
  nor _58437_ (_06960_, _06958_, _06909_);
  nor _58438_ (_06961_, _06960_, _06959_);
  and _58439_ (_06962_, _06961_, _06957_);
  nor _58440_ (_06963_, _06961_, _06957_);
  nor _58441_ (_06964_, _06963_, _06962_);
  not _58442_ (_06965_, _06964_);
  nor _58443_ (_06966_, _06965_, _06956_);
  and _58444_ (_06967_, _06965_, _06956_);
  nor _58445_ (_06968_, _06967_, _06966_);
  and _58446_ (_06969_, _06968_, _06955_);
  nor _58447_ (_06970_, _06968_, _06955_);
  nor _58448_ (_06971_, _06970_, _06969_);
  not _58449_ (_06972_, _06971_);
  nor _58450_ (_06973_, _06972_, _06942_);
  nor _58451_ (_06974_, _06936_, _06933_);
  not _58452_ (_06975_, _06974_);
  and _58453_ (_06976_, _06972_, _06942_);
  nor _58454_ (_06977_, _06976_, _06973_);
  and _58455_ (_06978_, _06977_, _06975_);
  nor _58456_ (_06979_, _06978_, _06973_);
  nor _58457_ (_06980_, _06953_, _06950_);
  not _58458_ (_06981_, _06980_);
  nor _58459_ (_06982_, _06969_, _06966_);
  not _58460_ (_06983_, _06982_);
  and _58461_ (_06984_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and _58462_ (_06985_, _06984_, _06909_);
  and _58463_ (_06986_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and _58464_ (_06987_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor _58465_ (_06988_, _06987_, _06986_);
  nor _58466_ (_06989_, _06988_, _06985_);
  nor _58467_ (_06990_, _06962_, _06959_);
  and _58468_ (_06991_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and _58469_ (_06992_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and _58470_ (_06993_, _06992_, _06991_);
  nor _58471_ (_06994_, _06992_, _06991_);
  nor _58472_ (_06995_, _06994_, _06993_);
  not _58473_ (_06996_, _06995_);
  nor _58474_ (_06997_, _06996_, _06990_);
  and _58475_ (_06998_, _06996_, _06990_);
  nor _58476_ (_06999_, _06998_, _06997_);
  and _58477_ (_07000_, _06999_, _06946_);
  nor _58478_ (_07001_, _06999_, _06946_);
  nor _58479_ (_07002_, _07001_, _07000_);
  and _58480_ (_07003_, _07002_, _06989_);
  nor _58481_ (_07004_, _07002_, _06989_);
  nor _58482_ (_07005_, _07004_, _07003_);
  and _58483_ (_07006_, _07005_, _06983_);
  nor _58484_ (_07007_, _07005_, _06983_);
  nor _58485_ (_07008_, _07007_, _07006_);
  and _58486_ (_07009_, _07008_, _06981_);
  nor _58487_ (_07010_, _07008_, _06981_);
  nor _58488_ (_07011_, _07010_, _07009_);
  not _58489_ (_07012_, _07011_);
  nor _58490_ (_07013_, _07012_, _06979_);
  nor _58491_ (_07014_, _07009_, _07006_);
  nor _58492_ (_07015_, _07000_, _06997_);
  not _58493_ (_07016_, _07015_);
  and _58494_ (_07017_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and _58495_ (_07018_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and _58496_ (_07019_, _07018_, _07017_);
  nor _58497_ (_07020_, _07018_, _07017_);
  nor _58498_ (_07021_, _07020_, _07019_);
  and _58499_ (_07022_, _07021_, _06985_);
  nor _58500_ (_07023_, _07021_, _06985_);
  nor _58501_ (_07024_, _07023_, _07022_);
  and _58502_ (_07025_, _07024_, _06993_);
  nor _58503_ (_07026_, _07024_, _06993_);
  nor _58504_ (_07027_, _07026_, _07025_);
  and _58505_ (_07028_, _07027_, _06984_);
  nor _58506_ (_07029_, _07027_, _06984_);
  nor _58507_ (_07030_, _07029_, _07028_);
  and _58508_ (_07031_, _07030_, _07003_);
  nor _58509_ (_07032_, _07030_, _07003_);
  nor _58510_ (_07033_, _07032_, _07031_);
  and _58511_ (_07034_, _07033_, _07016_);
  nor _58512_ (_07035_, _07033_, _07016_);
  nor _58513_ (_07036_, _07035_, _07034_);
  not _58514_ (_07037_, _07036_);
  nor _58515_ (_07038_, _07037_, _07014_);
  and _58516_ (_07039_, _07037_, _07014_);
  nor _58517_ (_07040_, _07039_, _07038_);
  and _58518_ (_07041_, _07040_, _07013_);
  nor _58519_ (_07042_, _07034_, _07031_);
  nor _58520_ (_07043_, _07025_, _07022_);
  not _58521_ (_07044_, _07043_);
  and _58522_ (_07045_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and _58523_ (_07046_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and _58524_ (_07047_, _07046_, _07045_);
  nor _58525_ (_07048_, _07046_, _07045_);
  nor _58526_ (_07049_, _07048_, _07047_);
  and _58527_ (_07050_, _07049_, _07019_);
  nor _58528_ (_07051_, _07049_, _07019_);
  nor _58529_ (_07052_, _07051_, _07050_);
  and _58530_ (_07053_, _07052_, _07028_);
  nor _58531_ (_07054_, _07052_, _07028_);
  nor _58532_ (_07055_, _07054_, _07053_);
  and _58533_ (_07056_, _07055_, _07044_);
  nor _58534_ (_07057_, _07055_, _07044_);
  nor _58535_ (_07058_, _07057_, _07056_);
  not _58536_ (_07059_, _07058_);
  nor _58537_ (_07060_, _07059_, _07042_);
  and _58538_ (_07061_, _07059_, _07042_);
  nor _58539_ (_07062_, _07061_, _07060_);
  and _58540_ (_07063_, _07062_, _07038_);
  nor _58541_ (_07064_, _07062_, _07038_);
  nor _58542_ (_07065_, _07064_, _07063_);
  and _58543_ (_07066_, _07065_, _07041_);
  nor _58544_ (_07067_, _07065_, _07041_);
  nor _58545_ (_07068_, _07067_, _07066_);
  and _58546_ (_07069_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and _58547_ (_07070_, _07069_, _06881_);
  and _58548_ (_07071_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and _58549_ (_07072_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor _58550_ (_07073_, _07072_, _06877_);
  nor _58551_ (_07074_, _07073_, _07070_);
  and _58552_ (_07075_, _07074_, _07071_);
  nor _58553_ (_07076_, _07075_, _07070_);
  not _58554_ (_07077_, _07076_);
  nor _58555_ (_07078_, _06883_, _06879_);
  nor _58556_ (_07079_, _07078_, _06884_);
  and _58557_ (_07080_, _07079_, _07077_);
  and _58558_ (_07081_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and _58559_ (_07082_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and _58560_ (_07083_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and _58561_ (_07084_, _07083_, _07082_);
  nor _58562_ (_07085_, _07083_, _07082_);
  nor _58563_ (_07086_, _07085_, _07084_);
  and _58564_ (_07087_, _07086_, _07081_);
  nor _58565_ (_07088_, _07086_, _07081_);
  nor _58566_ (_07089_, _07088_, _07087_);
  nor _58567_ (_07090_, _07079_, _07077_);
  nor _58568_ (_07091_, _07090_, _07080_);
  and _58569_ (_07092_, _07091_, _07089_);
  nor _58570_ (_07093_, _07092_, _07080_);
  nor _58571_ (_07094_, _06903_, _06901_);
  nor _58572_ (_07095_, _07094_, _06904_);
  not _58573_ (_07096_, _07095_);
  nor _58574_ (_07097_, _07096_, _07093_);
  and _58575_ (_07098_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and _58576_ (_07099_, _07098_, _06924_);
  nor _58577_ (_07100_, _07087_, _07084_);
  nor _58578_ (_07101_, _06924_, _06923_);
  nor _58579_ (_07102_, _07101_, _06925_);
  not _58580_ (_07103_, _07102_);
  nor _58581_ (_07104_, _07103_, _07100_);
  and _58582_ (_07105_, _07103_, _07100_);
  nor _58583_ (_07106_, _07105_, _07104_);
  and _58584_ (_07107_, _07106_, _07099_);
  nor _58585_ (_07108_, _07106_, _07099_);
  nor _58586_ (_07109_, _07108_, _07107_);
  and _58587_ (_07110_, _07096_, _07093_);
  nor _58588_ (_07111_, _07110_, _07097_);
  and _58589_ (_07112_, _07111_, _07109_);
  nor _58590_ (_07113_, _07112_, _07097_);
  nor _58591_ (_07114_, _06940_, _06938_);
  nor _58592_ (_07115_, _07114_, _06941_);
  not _58593_ (_07116_, _07115_);
  nor _58594_ (_07117_, _07116_, _07113_);
  nor _58595_ (_07118_, _07107_, _07104_);
  not _58596_ (_07119_, _07118_);
  and _58597_ (_07120_, _07116_, _07113_);
  nor _58598_ (_07121_, _07120_, _07117_);
  and _58599_ (_07122_, _07121_, _07119_);
  nor _58600_ (_07123_, _07122_, _07117_);
  nor _58601_ (_07124_, _06977_, _06975_);
  nor _58602_ (_07125_, _07124_, _06978_);
  not _58603_ (_07126_, _07125_);
  nor _58604_ (_07127_, _07126_, _07123_);
  and _58605_ (_07128_, _07012_, _06979_);
  nor _58606_ (_07129_, _07128_, _07013_);
  and _58607_ (_07130_, _07129_, _07127_);
  nor _58608_ (_07131_, _07040_, _07013_);
  nor _58609_ (_07132_, _07131_, _07041_);
  and _58610_ (_07133_, _07132_, _07130_);
  and _58611_ (_07134_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and _58612_ (_07135_, _07134_, _07069_);
  and _58613_ (_07136_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor _58614_ (_07137_, _07134_, _07069_);
  nor _58615_ (_07138_, _07137_, _07135_);
  and _58616_ (_07139_, _07138_, _07136_);
  nor _58617_ (_07140_, _07139_, _07135_);
  not _58618_ (_07141_, _07140_);
  nor _58619_ (_07142_, _07074_, _07071_);
  nor _58620_ (_07143_, _07142_, _07075_);
  and _58621_ (_07144_, _07143_, _07141_);
  and _58622_ (_07145_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and _58623_ (_07146_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and _58624_ (_07147_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and _58625_ (_07148_, _07147_, _07146_);
  nor _58626_ (_07149_, _07147_, _07146_);
  nor _58627_ (_07150_, _07149_, _07148_);
  and _58628_ (_07151_, _07150_, _07145_);
  nor _58629_ (_07152_, _07150_, _07145_);
  nor _58630_ (_07153_, _07152_, _07151_);
  nor _58631_ (_07154_, _07143_, _07141_);
  nor _58632_ (_07155_, _07154_, _07144_);
  and _58633_ (_07156_, _07155_, _07153_);
  nor _58634_ (_07157_, _07156_, _07144_);
  not _58635_ (_07158_, _07157_);
  nor _58636_ (_07159_, _07091_, _07089_);
  nor _58637_ (_07160_, _07159_, _07092_);
  and _58638_ (_07161_, _07160_, _07158_);
  nor _58639_ (_07162_, _07151_, _07148_);
  and _58640_ (_07163_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and _58641_ (_07164_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor _58642_ (_07165_, _07164_, _07163_);
  nor _58643_ (_07166_, _07165_, _07099_);
  not _58644_ (_07167_, _07166_);
  nor _58645_ (_07168_, _07167_, _07162_);
  and _58646_ (_07169_, _07167_, _07162_);
  nor _58647_ (_07170_, _07169_, _07168_);
  nor _58648_ (_07171_, _07160_, _07158_);
  nor _58649_ (_07172_, _07171_, _07161_);
  and _58650_ (_07173_, _07172_, _07170_);
  nor _58651_ (_07174_, _07173_, _07161_);
  nor _58652_ (_07175_, _07111_, _07109_);
  nor _58653_ (_07176_, _07175_, _07112_);
  not _58654_ (_07177_, _07176_);
  nor _58655_ (_07178_, _07177_, _07174_);
  and _58656_ (_07179_, _07177_, _07174_);
  nor _58657_ (_07180_, _07179_, _07178_);
  and _58658_ (_07181_, _07180_, _07168_);
  nor _58659_ (_07182_, _07181_, _07178_);
  nor _58660_ (_07183_, _07121_, _07119_);
  nor _58661_ (_07184_, _07183_, _07122_);
  not _58662_ (_07185_, _07184_);
  nor _58663_ (_07186_, _07185_, _07182_);
  and _58664_ (_07187_, _07126_, _07123_);
  nor _58665_ (_07188_, _07187_, _07127_);
  and _58666_ (_07189_, _07188_, _07186_);
  nor _58667_ (_07190_, _07129_, _07127_);
  nor _58668_ (_07191_, _07190_, _07130_);
  and _58669_ (_07192_, _07191_, _07189_);
  nor _58670_ (_07193_, _07191_, _07189_);
  nor _58671_ (_07194_, _07193_, _07192_);
  and _58672_ (_07195_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and _58673_ (_07196_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and _58674_ (_07197_, _07196_, _07195_);
  and _58675_ (_07198_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor _58676_ (_07199_, _07196_, _07195_);
  nor _58677_ (_07200_, _07199_, _07197_);
  and _58678_ (_07201_, _07200_, _07198_);
  nor _58679_ (_07202_, _07201_, _07197_);
  not _58680_ (_07203_, _07202_);
  nor _58681_ (_07204_, _07138_, _07136_);
  nor _58682_ (_07205_, _07204_, _07139_);
  and _58683_ (_07206_, _07205_, _07203_);
  and _58684_ (_07207_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and _58685_ (_07208_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and _58686_ (_07209_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and _58687_ (_07210_, _07209_, _07208_);
  nor _58688_ (_07211_, _07209_, _07208_);
  nor _58689_ (_07212_, _07211_, _07210_);
  and _58690_ (_07213_, _07212_, _07207_);
  nor _58691_ (_07214_, _07212_, _07207_);
  nor _58692_ (_07215_, _07214_, _07213_);
  nor _58693_ (_07216_, _07205_, _07203_);
  nor _58694_ (_07217_, _07216_, _07206_);
  and _58695_ (_07218_, _07217_, _07215_);
  nor _58696_ (_07219_, _07218_, _07206_);
  not _58697_ (_07220_, _07219_);
  nor _58698_ (_07221_, _07155_, _07153_);
  nor _58699_ (_07222_, _07221_, _07156_);
  and _58700_ (_07223_, _07222_, _07220_);
  not _58701_ (_07224_, _07098_);
  nor _58702_ (_07225_, _07213_, _07210_);
  nor _58703_ (_07226_, _07225_, _07224_);
  and _58704_ (_07227_, _07225_, _07224_);
  nor _58705_ (_07228_, _07227_, _07226_);
  nor _58706_ (_07229_, _07222_, _07220_);
  nor _58707_ (_07230_, _07229_, _07223_);
  and _58708_ (_07231_, _07230_, _07228_);
  nor _58709_ (_07232_, _07231_, _07223_);
  not _58710_ (_07233_, _07232_);
  nor _58711_ (_07234_, _07172_, _07170_);
  nor _58712_ (_07235_, _07234_, _07173_);
  and _58713_ (_07236_, _07235_, _07233_);
  nor _58714_ (_07237_, _07235_, _07233_);
  nor _58715_ (_07238_, _07237_, _07236_);
  and _58716_ (_07239_, _07238_, _07226_);
  nor _58717_ (_07240_, _07239_, _07236_);
  nor _58718_ (_07241_, _07180_, _07168_);
  nor _58719_ (_07242_, _07241_, _07181_);
  not _58720_ (_07243_, _07242_);
  nor _58721_ (_07244_, _07243_, _07240_);
  and _58722_ (_07245_, _07185_, _07182_);
  nor _58723_ (_07246_, _07245_, _07186_);
  and _58724_ (_07247_, _07246_, _07244_);
  nor _58725_ (_07248_, _07188_, _07186_);
  nor _58726_ (_07249_, _07248_, _07189_);
  and _58727_ (_07250_, _07249_, _07247_);
  nor _58728_ (_07251_, _07249_, _07247_);
  nor _58729_ (_07252_, _07251_, _07250_);
  and _58730_ (_07253_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and _58731_ (_07254_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and _58732_ (_07255_, _07254_, _07253_);
  and _58733_ (_07256_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor _58734_ (_07257_, _07254_, _07253_);
  nor _58735_ (_07258_, _07257_, _07255_);
  and _58736_ (_07259_, _07258_, _07256_);
  nor _58737_ (_07260_, _07259_, _07255_);
  not _58738_ (_07261_, _07260_);
  nor _58739_ (_07262_, _07200_, _07198_);
  nor _58740_ (_07263_, _07262_, _07201_);
  and _58741_ (_07264_, _07263_, _07261_);
  and _58742_ (_07265_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and _58743_ (_07266_, _07265_, _07209_);
  and _58744_ (_07267_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and _58745_ (_07268_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor _58746_ (_07269_, _07268_, _07267_);
  nor _58747_ (_07270_, _07269_, _07266_);
  nor _58748_ (_07271_, _07263_, _07261_);
  nor _58749_ (_07272_, _07271_, _07264_);
  and _58750_ (_07273_, _07272_, _07270_);
  nor _58751_ (_07274_, _07273_, _07264_);
  not _58752_ (_07275_, _07274_);
  nor _58753_ (_07276_, _07217_, _07215_);
  nor _58754_ (_07277_, _07276_, _07218_);
  and _58755_ (_07278_, _07277_, _07275_);
  nor _58756_ (_07279_, _07277_, _07275_);
  nor _58757_ (_07280_, _07279_, _07278_);
  and _58758_ (_07281_, _07280_, _07266_);
  nor _58759_ (_07282_, _07281_, _07278_);
  not _58760_ (_07283_, _07282_);
  nor _58761_ (_07284_, _07230_, _07228_);
  nor _58762_ (_07285_, _07284_, _07231_);
  and _58763_ (_07286_, _07285_, _07283_);
  nor _58764_ (_07287_, _07238_, _07226_);
  nor _58765_ (_07288_, _07287_, _07239_);
  and _58766_ (_07289_, _07288_, _07286_);
  and _58767_ (_07290_, _07243_, _07240_);
  nor _58768_ (_07291_, _07290_, _07244_);
  and _58769_ (_07292_, _07291_, _07289_);
  nor _58770_ (_07293_, _07246_, _07244_);
  nor _58771_ (_07294_, _07293_, _07247_);
  nor _58772_ (_07295_, _07294_, _07292_);
  and _58773_ (_07296_, _07294_, _07292_);
  not _58774_ (_07297_, _07296_);
  and _58775_ (_07298_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and _58776_ (_07299_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and _58777_ (_07300_, _07299_, _07298_);
  and _58778_ (_07301_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor _58779_ (_07302_, _07299_, _07298_);
  nor _58780_ (_07303_, _07302_, _07300_);
  and _58781_ (_07304_, _07303_, _07301_);
  nor _58782_ (_07305_, _07304_, _07300_);
  not _58783_ (_07306_, _07305_);
  nor _58784_ (_07307_, _07258_, _07256_);
  nor _58785_ (_07308_, _07307_, _07259_);
  and _58786_ (_07309_, _07308_, _07306_);
  nor _58787_ (_07310_, _07308_, _07306_);
  nor _58788_ (_07311_, _07310_, _07309_);
  and _58789_ (_07312_, _07311_, _07265_);
  nor _58790_ (_07313_, _07312_, _07309_);
  not _58791_ (_07314_, _07313_);
  nor _58792_ (_07315_, _07272_, _07270_);
  nor _58793_ (_07316_, _07315_, _07273_);
  and _58794_ (_07317_, _07316_, _07314_);
  nor _58795_ (_07318_, _07280_, _07266_);
  nor _58796_ (_07319_, _07318_, _07281_);
  and _58797_ (_07320_, _07319_, _07317_);
  nor _58798_ (_07321_, _07285_, _07283_);
  nor _58799_ (_07322_, _07321_, _07286_);
  and _58800_ (_07323_, _07322_, _07320_);
  nor _58801_ (_07324_, _07288_, _07286_);
  nor _58802_ (_07325_, _07324_, _07289_);
  and _58803_ (_07326_, _07325_, _07323_);
  nor _58804_ (_07327_, _07291_, _07289_);
  nor _58805_ (_07328_, _07327_, _07292_);
  and _58806_ (_07329_, _07328_, _07326_);
  and _58807_ (_07330_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and _58808_ (_07331_, _07330_, _07299_);
  nor _58809_ (_07332_, _07303_, _07301_);
  nor _58810_ (_07333_, _07332_, _07304_);
  and _58811_ (_07334_, _07333_, _07331_);
  nor _58812_ (_07335_, _07311_, _07265_);
  nor _58813_ (_07336_, _07335_, _07312_);
  and _58814_ (_07337_, _07336_, _07334_);
  nor _58815_ (_07338_, _07316_, _07314_);
  nor _58816_ (_07339_, _07338_, _07317_);
  and _58817_ (_07340_, _07339_, _07337_);
  nor _58818_ (_07341_, _07319_, _07317_);
  nor _58819_ (_07342_, _07341_, _07320_);
  and _58820_ (_07343_, _07342_, _07340_);
  nor _58821_ (_07344_, _07322_, _07320_);
  nor _58822_ (_07345_, _07344_, _07323_);
  and _58823_ (_07346_, _07345_, _07343_);
  nor _58824_ (_07347_, _07325_, _07323_);
  nor _58825_ (_07348_, _07347_, _07326_);
  and _58826_ (_07349_, _07348_, _07346_);
  nor _58827_ (_07350_, _07328_, _07326_);
  nor _58828_ (_07351_, _07350_, _07329_);
  and _58829_ (_07352_, _07351_, _07349_);
  nor _58830_ (_07353_, _07352_, _07329_);
  and _58831_ (_07354_, _07353_, _07297_);
  nor _58832_ (_07355_, _07354_, _07295_);
  and _58833_ (_07356_, _07355_, _07252_);
  nor _58834_ (_07357_, _07356_, _07250_);
  not _58835_ (_07358_, _07357_);
  and _58836_ (_07359_, _07358_, _07194_);
  nor _58837_ (_07360_, _07359_, _07192_);
  not _58838_ (_07361_, _07360_);
  nor _58839_ (_07362_, _07132_, _07130_);
  nor _58840_ (_07363_, _07362_, _07133_);
  and _58841_ (_07364_, _07363_, _07361_);
  nor _58842_ (_07365_, _07364_, _07133_);
  not _58843_ (_07366_, _07365_);
  and _58844_ (_07367_, _07366_, _07068_);
  nor _58845_ (_07368_, _07367_, _07066_);
  not _58846_ (_07369_, _07368_);
  and _58847_ (_07370_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not _58848_ (_07371_, _07370_);
  nor _58849_ (_07372_, _07371_, _07018_);
  nor _58850_ (_07373_, _07372_, _07050_);
  nor _58851_ (_07374_, _07056_, _07053_);
  nor _58852_ (_07375_, _07374_, _07373_);
  and _58853_ (_07376_, _07374_, _07373_);
  nor _58854_ (_07377_, _07376_, _07375_);
  not _58855_ (_07378_, _07377_);
  nor _58856_ (_07379_, _07063_, _07060_);
  and _58857_ (_07380_, _07379_, _07378_);
  nor _58858_ (_07381_, _07379_, _07378_);
  nor _58859_ (_07382_, _07381_, _07380_);
  and _58860_ (_07383_, _07382_, _07369_);
  or _58861_ (_07384_, _07375_, _07047_);
  or _58862_ (_07385_, _07384_, _07381_);
  or _58863_ (_07386_, _07385_, _07383_);
  or _58864_ (_07387_, _07386_, _06875_);
  and _58865_ (_07388_, _07387_, _03710_);
  and _58866_ (_07389_, _07388_, _06874_);
  not _58867_ (_07390_, _06838_);
  not _58868_ (_07391_, _05910_);
  nor _58869_ (_07392_, _05938_, _07391_);
  or _58870_ (_07393_, _07392_, _06841_);
  and _58871_ (_07394_, _07393_, _03505_);
  or _58872_ (_07395_, _07394_, _07390_);
  or _58873_ (_07396_, _07395_, _07389_);
  and _58874_ (_07397_, _07396_, _06839_);
  or _58875_ (_07398_, _07397_, _04481_);
  and _58876_ (_07399_, _06069_, _05248_);
  not _58877_ (_07400_, _04481_);
  or _58878_ (_07401_, _06829_, _07400_);
  or _58879_ (_07402_, _07401_, _07399_);
  and _58880_ (_07403_, _07402_, _03589_);
  and _58881_ (_07404_, _07403_, _07398_);
  and _58882_ (_07405_, _03603_, _03168_);
  nor _58883_ (_07406_, _06363_, _06830_);
  or _58884_ (_07407_, _07406_, _06829_);
  and _58885_ (_07408_, _07407_, _03222_);
  or _58886_ (_07409_, _07408_, _07405_);
  or _58887_ (_07410_, _07409_, _07404_);
  not _58888_ (_07411_, _07405_);
  not _58889_ (_07412_, \oc8051_golden_model_1.B [1]);
  nor _58890_ (_07413_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor _58891_ (_07414_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and _58892_ (_07415_, _07414_, _07413_);
  and _58893_ (_07416_, _07415_, _07412_);
  nor _58894_ (_07417_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not _58895_ (_07418_, \oc8051_golden_model_1.B [0]);
  and _58896_ (_07419_, _07418_, \oc8051_golden_model_1.ACC [7]);
  and _58897_ (_07420_, _07419_, _07417_);
  and _58898_ (_07421_, _07420_, _07416_);
  or _58899_ (_07422_, _07418_, \oc8051_golden_model_1.ACC [7]);
  and _58900_ (_07423_, _07422_, _07417_);
  and _58901_ (_07424_, _07423_, _07416_);
  or _58902_ (_07425_, _07424_, _06075_);
  not _58903_ (_07426_, \oc8051_golden_model_1.B [2]);
  not _58904_ (_07427_, \oc8051_golden_model_1.B [3]);
  nor _58905_ (_07428_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and _58906_ (_07429_, _07428_, _07413_);
  and _58907_ (_07430_, _07429_, _07427_);
  and _58908_ (_07431_, _07430_, _07426_);
  not _58909_ (_07432_, _07431_);
  not _58910_ (_07433_, \oc8051_golden_model_1.ACC [6]);
  and _58911_ (_07434_, \oc8051_golden_model_1.B [0], _07433_);
  nor _58912_ (_07435_, _07434_, _06075_);
  nor _58913_ (_07436_, _07435_, _07412_);
  nor _58914_ (_07437_, _07436_, _07432_);
  nor _58915_ (_07438_, _07437_, _07425_);
  nor _58916_ (_07439_, _07438_, _07421_);
  and _58917_ (_07440_, _07437_, \oc8051_golden_model_1.B [0]);
  nor _58918_ (_07441_, _07440_, _07433_);
  and _58919_ (_07442_, _07441_, _07412_);
  nor _58920_ (_07443_, _07441_, _07412_);
  nor _58921_ (_07444_, _07443_, _07442_);
  nor _58922_ (_07445_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor _58923_ (_07446_, _07445_, _07069_);
  nor _58924_ (_07447_, _07446_, \oc8051_golden_model_1.ACC [4]);
  nor _58925_ (_07448_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and _58926_ (_07449_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor _58927_ (_07450_, _07449_, _07418_);
  nor _58928_ (_07451_, _07450_, _07448_);
  nor _58929_ (_07452_, _07451_, _07447_);
  not _58930_ (_07453_, _07452_);
  and _58931_ (_07454_, _07453_, _07444_);
  nor _58932_ (_07455_, _07439_, \oc8051_golden_model_1.B [2]);
  nor _58933_ (_07456_, _07455_, _07442_);
  not _58934_ (_07457_, _07456_);
  nor _58935_ (_07458_, _07457_, _07454_);
  and _58936_ (_07459_, \oc8051_golden_model_1.B [2], _06075_);
  nor _58937_ (_07460_, _07459_, \oc8051_golden_model_1.B [7]);
  and _58938_ (_07461_, _07460_, _07415_);
  not _58939_ (_07462_, _07461_);
  nor _58940_ (_07463_, _07462_, _07458_);
  nor _58941_ (_07464_, _07463_, _07439_);
  nor _58942_ (_07465_, _07464_, _07421_);
  and _58943_ (_07466_, _07429_, \oc8051_golden_model_1.ACC [7]);
  nor _58944_ (_07467_, _07466_, _07430_);
  nor _58945_ (_07468_, _07453_, _07444_);
  nor _58946_ (_07469_, _07468_, _07454_);
  not _58947_ (_07470_, _07469_);
  and _58948_ (_07471_, _07470_, _07463_);
  nor _58949_ (_07472_, _07463_, _07441_);
  nor _58950_ (_07473_, _07472_, _07471_);
  and _58951_ (_07474_, _07473_, _07426_);
  nor _58952_ (_07475_, _07473_, _07426_);
  nor _58953_ (_07476_, _07475_, _07474_);
  not _58954_ (_07477_, _07476_);
  not _58955_ (_07478_, \oc8051_golden_model_1.ACC [5]);
  nor _58956_ (_07479_, _07463_, _07478_);
  and _58957_ (_07480_, _07463_, _07446_);
  or _58958_ (_07481_, _07480_, _07479_);
  and _58959_ (_07482_, _07481_, _07412_);
  nor _58960_ (_07483_, _07481_, _07412_);
  not _58961_ (_07484_, \oc8051_golden_model_1.ACC [4]);
  and _58962_ (_07485_, \oc8051_golden_model_1.B [0], _07484_);
  nor _58963_ (_07486_, _07485_, _07483_);
  nor _58964_ (_07487_, _07486_, _07482_);
  nor _58965_ (_07488_, _07487_, _07477_);
  nor _58966_ (_07489_, _07465_, \oc8051_golden_model_1.B [3]);
  nor _58967_ (_07490_, _07489_, _07474_);
  not _58968_ (_07491_, _07490_);
  nor _58969_ (_07492_, _07491_, _07488_);
  nor _58970_ (_07493_, _07492_, _07467_);
  nor _58971_ (_07494_, _07493_, _07465_);
  nor _58972_ (_07495_, _07494_, _07421_);
  not _58973_ (_07496_, _07493_);
  and _58974_ (_07497_, _07487_, _07477_);
  nor _58975_ (_07498_, _07497_, _07488_);
  nor _58976_ (_07499_, _07498_, _07496_);
  nor _58977_ (_07500_, _07493_, _07473_);
  nor _58978_ (_07501_, _07500_, _07499_);
  and _58979_ (_07502_, _07501_, _07427_);
  nor _58980_ (_07503_, _07501_, _07427_);
  nor _58981_ (_07504_, _07503_, _07502_);
  not _58982_ (_07505_, _07504_);
  nor _58983_ (_07506_, _07493_, _07481_);
  nor _58984_ (_07507_, _07483_, _07482_);
  and _58985_ (_07508_, _07507_, _07485_);
  nor _58986_ (_07509_, _07507_, _07485_);
  nor _58987_ (_07510_, _07509_, _07508_);
  and _58988_ (_07511_, _07510_, _07493_);
  or _58989_ (_07512_, _07511_, _07506_);
  nor _58990_ (_07513_, _07512_, \oc8051_golden_model_1.B [2]);
  and _58991_ (_07514_, _07512_, \oc8051_golden_model_1.B [2]);
  nor _58992_ (_07515_, _07493_, _07484_);
  nor _58993_ (_07516_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor _58994_ (_07517_, _07516_, _07195_);
  and _58995_ (_07518_, _07493_, _07517_);
  or _58996_ (_07519_, _07518_, _07515_);
  and _58997_ (_07520_, _07519_, _07412_);
  nor _58998_ (_07521_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor _58999_ (_07522_, _07521_, _07253_);
  nor _59000_ (_07523_, _07522_, \oc8051_golden_model_1.ACC [2]);
  nor _59001_ (_07524_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and _59002_ (_07525_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor _59003_ (_07526_, _07525_, _07418_);
  nor _59004_ (_07527_, _07526_, _07524_);
  nor _59005_ (_07528_, _07527_, _07523_);
  not _59006_ (_07529_, _07528_);
  nor _59007_ (_07530_, _07519_, _07412_);
  nor _59008_ (_07531_, _07530_, _07520_);
  and _59009_ (_07532_, _07531_, _07529_);
  nor _59010_ (_07533_, _07532_, _07520_);
  nor _59011_ (_07534_, _07533_, _07514_);
  nor _59012_ (_07535_, _07534_, _07513_);
  nor _59013_ (_07536_, _07535_, _07505_);
  nor _59014_ (_07537_, _07495_, \oc8051_golden_model_1.B [4]);
  nor _59015_ (_07538_, _07537_, _07502_);
  not _59016_ (_07539_, _07538_);
  nor _59017_ (_07540_, _07539_, _07536_);
  not _59018_ (_07541_, \oc8051_golden_model_1.B [5]);
  and _59019_ (_07542_, _07428_, _07541_);
  and _59020_ (_07543_, \oc8051_golden_model_1.B [4], _06075_);
  not _59021_ (_07544_, _07543_);
  and _59022_ (_07545_, _07544_, _07542_);
  not _59023_ (_07546_, _07545_);
  nor _59024_ (_07547_, _07546_, _07540_);
  nor _59025_ (_07548_, _07547_, _07495_);
  nor _59026_ (_07549_, _07548_, _07421_);
  not _59027_ (_07550_, \oc8051_golden_model_1.B [4]);
  and _59028_ (_07551_, _07535_, _07505_);
  nor _59029_ (_07552_, _07551_, _07536_);
  not _59030_ (_07553_, _07552_);
  and _59031_ (_07554_, _07553_, _07547_);
  nor _59032_ (_07555_, _07547_, _07501_);
  nor _59033_ (_07556_, _07555_, _07554_);
  and _59034_ (_07557_, _07556_, _07550_);
  nor _59035_ (_07558_, _07556_, _07550_);
  nor _59036_ (_07559_, _07558_, _07557_);
  not _59037_ (_07560_, _07559_);
  nor _59038_ (_07561_, _07547_, _07512_);
  nor _59039_ (_07562_, _07514_, _07513_);
  and _59040_ (_07563_, _07562_, _07533_);
  nor _59041_ (_07564_, _07562_, _07533_);
  nor _59042_ (_07565_, _07564_, _07563_);
  not _59043_ (_07566_, _07565_);
  and _59044_ (_07567_, _07566_, _07547_);
  nor _59045_ (_07568_, _07567_, _07561_);
  nor _59046_ (_07569_, _07568_, \oc8051_golden_model_1.B [3]);
  and _59047_ (_07570_, _07568_, \oc8051_golden_model_1.B [3]);
  nor _59048_ (_07571_, _07531_, _07529_);
  nor _59049_ (_07572_, _07571_, _07532_);
  not _59050_ (_07573_, _07572_);
  and _59051_ (_07574_, _07573_, _07547_);
  nor _59052_ (_07575_, _07547_, _07519_);
  nor _59053_ (_07576_, _07575_, _07574_);
  and _59054_ (_07577_, _07576_, _07426_);
  not _59055_ (_07578_, \oc8051_golden_model_1.ACC [3]);
  nor _59056_ (_07579_, _07547_, _07578_);
  and _59057_ (_07580_, _07547_, _07522_);
  or _59058_ (_07581_, _07580_, _07579_);
  and _59059_ (_07582_, _07581_, _07412_);
  nor _59060_ (_07583_, _07581_, _07412_);
  not _59061_ (_07584_, \oc8051_golden_model_1.ACC [2]);
  and _59062_ (_07585_, \oc8051_golden_model_1.B [0], _07584_);
  nor _59063_ (_07586_, _07585_, _07583_);
  nor _59064_ (_07587_, _07586_, _07582_);
  nor _59065_ (_07588_, _07576_, _07426_);
  nor _59066_ (_07589_, _07588_, _07577_);
  not _59067_ (_07590_, _07589_);
  nor _59068_ (_07591_, _07590_, _07587_);
  nor _59069_ (_07592_, _07591_, _07577_);
  nor _59070_ (_07593_, _07592_, _07570_);
  nor _59071_ (_07594_, _07593_, _07569_);
  nor _59072_ (_07595_, _07594_, _07560_);
  nor _59073_ (_07596_, _07549_, \oc8051_golden_model_1.B [5]);
  nor _59074_ (_07597_, _07596_, _07557_);
  not _59075_ (_07598_, _07597_);
  nor _59076_ (_07599_, _07598_, _07595_);
  not _59077_ (_07600_, _07599_);
  not _59078_ (_07601_, _07428_);
  and _59079_ (_07602_, \oc8051_golden_model_1.B [5], _06075_);
  nor _59080_ (_07603_, _07602_, _07601_);
  and _59081_ (_07604_, _07603_, _07600_);
  nor _59082_ (_07605_, _07604_, _07549_);
  nor _59083_ (_07606_, _07605_, _07421_);
  nor _59084_ (_07607_, _07606_, \oc8051_golden_model_1.B [6]);
  and _59085_ (_07608_, \oc8051_golden_model_1.B [6], _06075_);
  not _59086_ (_07609_, _07604_);
  and _59087_ (_07610_, _07594_, _07560_);
  nor _59088_ (_07611_, _07610_, _07595_);
  nor _59089_ (_07612_, _07611_, _07609_);
  nor _59090_ (_07613_, _07604_, _07556_);
  nor _59091_ (_07614_, _07613_, _07612_);
  and _59092_ (_07615_, _07614_, _07541_);
  nor _59093_ (_07616_, _07614_, _07541_);
  nor _59094_ (_07617_, _07616_, _07615_);
  not _59095_ (_07618_, _07617_);
  nor _59096_ (_07619_, _07570_, _07569_);
  nor _59097_ (_07620_, _07619_, _07592_);
  and _59098_ (_07621_, _07619_, _07592_);
  or _59099_ (_07622_, _07621_, _07620_);
  nor _59100_ (_07623_, _07622_, _07609_);
  and _59101_ (_07624_, _07609_, _07568_);
  nor _59102_ (_07625_, _07624_, _07623_);
  and _59103_ (_07626_, _07625_, _07550_);
  nor _59104_ (_07627_, _07625_, _07550_);
  and _59105_ (_07628_, _07590_, _07587_);
  nor _59106_ (_07629_, _07628_, _07591_);
  nor _59107_ (_07630_, _07629_, _07609_);
  nor _59108_ (_07631_, _07604_, _07576_);
  nor _59109_ (_07632_, _07631_, _07630_);
  and _59110_ (_07633_, _07632_, _07427_);
  nor _59111_ (_07634_, _07583_, _07582_);
  nor _59112_ (_07635_, _07634_, _07585_);
  and _59113_ (_07636_, _07634_, _07585_);
  or _59114_ (_07637_, _07636_, _07635_);
  nor _59115_ (_07638_, _07637_, _07609_);
  nor _59116_ (_07639_, _07604_, _07581_);
  nor _59117_ (_07640_, _07639_, _07638_);
  and _59118_ (_07641_, _07640_, _07426_);
  nor _59119_ (_07642_, _07640_, _07426_);
  nor _59120_ (_07643_, _07604_, _07584_);
  nor _59121_ (_07644_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor _59122_ (_07645_, _07644_, _07298_);
  and _59123_ (_07646_, _07604_, _07645_);
  or _59124_ (_07647_, _07646_, _07643_);
  and _59125_ (_07648_, _07647_, _07412_);
  and _59126_ (_07649_, \oc8051_golden_model_1.B [0], _03274_);
  not _59127_ (_07650_, _07649_);
  nor _59128_ (_07651_, _07647_, _07412_);
  nor _59129_ (_07652_, _07651_, _07648_);
  and _59130_ (_07653_, _07652_, _07650_);
  nor _59131_ (_07654_, _07653_, _07648_);
  nor _59132_ (_07655_, _07654_, _07642_);
  nor _59133_ (_07656_, _07655_, _07641_);
  nor _59134_ (_07657_, _07632_, _07427_);
  nor _59135_ (_07658_, _07657_, _07633_);
  not _59136_ (_07659_, _07658_);
  nor _59137_ (_07660_, _07659_, _07656_);
  nor _59138_ (_07661_, _07660_, _07633_);
  nor _59139_ (_07662_, _07661_, _07627_);
  nor _59140_ (_07663_, _07662_, _07626_);
  nor _59141_ (_07664_, _07663_, _07618_);
  nor _59142_ (_07665_, _07664_, _07615_);
  nor _59143_ (_07666_, _07665_, _07608_);
  nor _59144_ (_07667_, _07666_, _07607_);
  nor _59145_ (_07668_, _07667_, \oc8051_golden_model_1.B [7]);
  nor _59146_ (_07669_, _07668_, _07606_);
  or _59147_ (_07670_, _07669_, _07421_);
  nor _59148_ (_07671_, _07670_, \oc8051_golden_model_1.B [7]);
  nor _59149_ (_07672_, _07671_, _07370_);
  not _59150_ (_07673_, \oc8051_golden_model_1.B [6]);
  not _59151_ (_07674_, _07668_);
  and _59152_ (_07675_, _07663_, _07618_);
  nor _59153_ (_07676_, _07675_, _07664_);
  nor _59154_ (_07677_, _07676_, _07674_);
  nor _59155_ (_07678_, _07668_, _07614_);
  nor _59156_ (_07679_, _07678_, _07677_);
  nor _59157_ (_07680_, _07679_, _07673_);
  not _59158_ (_07681_, _07680_);
  nor _59159_ (_07682_, _07681_, _07672_);
  nor _59160_ (_07683_, _07642_, _07641_);
  and _59161_ (_07684_, _07683_, _07654_);
  nor _59162_ (_07685_, _07683_, _07654_);
  or _59163_ (_07686_, _07685_, _07684_);
  and _59164_ (_07687_, _07686_, _07668_);
  and _59165_ (_07688_, _07674_, _07640_);
  nor _59166_ (_07689_, _07688_, _07687_);
  nor _59167_ (_07690_, _07689_, \oc8051_golden_model_1.B [3]);
  and _59168_ (_07691_, _07689_, \oc8051_golden_model_1.B [3]);
  nor _59169_ (_07692_, _07691_, _07690_);
  nor _59170_ (_07693_, _07652_, _07650_);
  or _59171_ (_07694_, _07693_, _07653_);
  and _59172_ (_07695_, _07694_, _07668_);
  nor _59173_ (_07696_, _07668_, _07647_);
  nor _59174_ (_07697_, _07696_, _07695_);
  nor _59175_ (_07698_, _07697_, _07426_);
  and _59176_ (_07699_, _07697_, _07426_);
  nor _59177_ (_07700_, _07699_, _07698_);
  and _59178_ (_07701_, _07700_, _07692_);
  nor _59179_ (_07702_, _07668_, \oc8051_golden_model_1.ACC [1]);
  and _59180_ (_07703_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor _59181_ (_07704_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  or _59182_ (_07705_, _07704_, _07703_);
  and _59183_ (_07706_, _07668_, _07705_);
  nor _59184_ (_07707_, _07706_, _07702_);
  and _59185_ (_07708_, _07707_, _07412_);
  nor _59186_ (_07709_, _07707_, _07412_);
  and _59187_ (_07710_, _07418_, \oc8051_golden_model_1.ACC [0]);
  not _59188_ (_07711_, _07710_);
  nor _59189_ (_07712_, _07711_, _07709_);
  nor _59190_ (_07713_, _07712_, _07708_);
  and _59191_ (_07714_, _07713_, _07701_);
  not _59192_ (_07715_, _07714_);
  and _59193_ (_07716_, _07698_, _07692_);
  nor _59194_ (_07717_, _07716_, _07691_);
  and _59195_ (_07718_, _07717_, _07715_);
  and _59196_ (_07719_, _07679_, _07673_);
  nor _59197_ (_07720_, _07719_, _07680_);
  not _59198_ (_07721_, _07720_);
  nor _59199_ (_07722_, _07721_, _07672_);
  and _59200_ (_07723_, _07659_, _07656_);
  or _59201_ (_07724_, _07723_, _07660_);
  and _59202_ (_07725_, _07724_, _07668_);
  nor _59203_ (_07726_, _07668_, _07632_);
  nor _59204_ (_07727_, _07726_, _07725_);
  nor _59205_ (_07728_, _07727_, _07550_);
  and _59206_ (_07729_, _07727_, _07550_);
  nor _59207_ (_07730_, _07729_, _07728_);
  nor _59208_ (_07731_, _07627_, _07626_);
  nor _59209_ (_07732_, _07731_, _07661_);
  and _59210_ (_07733_, _07731_, _07661_);
  or _59211_ (_07734_, _07733_, _07732_);
  and _59212_ (_07735_, _07734_, _07668_);
  and _59213_ (_07736_, _07674_, _07625_);
  nor _59214_ (_07737_, _07736_, _07735_);
  and _59215_ (_07738_, _07737_, \oc8051_golden_model_1.B [5]);
  nor _59216_ (_07739_, _07737_, \oc8051_golden_model_1.B [5]);
  nor _59217_ (_07740_, _07739_, _07738_);
  and _59218_ (_07741_, _07740_, _07730_);
  and _59219_ (_07742_, _07741_, _07722_);
  not _59220_ (_07743_, _07742_);
  nor _59221_ (_07744_, _07743_, _07718_);
  and _59222_ (_07745_, _07606_, \oc8051_golden_model_1.B [7]);
  and _59223_ (_07746_, _07740_, _07728_);
  nor _59224_ (_07747_, _07746_, _07738_);
  not _59225_ (_07748_, _07747_);
  and _59226_ (_07749_, _07748_, _07722_);
  or _59227_ (_07750_, _07749_, _07745_);
  or _59228_ (_07751_, _07750_, _07744_);
  nor _59229_ (_07752_, _07751_, _07682_);
  and _59230_ (_07753_, \oc8051_golden_model_1.B [0], _03335_);
  not _59231_ (_07754_, _07753_);
  nor _59232_ (_07755_, _07709_, _07708_);
  and _59233_ (_07756_, _07755_, _07754_);
  and _59234_ (_07757_, _07756_, _07711_);
  and _59235_ (_07758_, _07757_, _07701_);
  and _59236_ (_07759_, _07758_, _07742_);
  nor _59237_ (_07760_, _07759_, _07752_);
  or _59238_ (_07761_, _07760_, _07421_);
  and _59239_ (_07762_, _07761_, _07670_);
  or _59240_ (_07763_, _07762_, _07411_);
  and _59241_ (_07764_, _07763_, _07410_);
  or _59242_ (_07765_, _07764_, _03601_);
  not _59243_ (_07766_, _03600_);
  and _59244_ (_07767_, _06171_, _05248_);
  or _59245_ (_07768_, _07767_, _06829_);
  or _59246_ (_07769_, _07768_, _05886_);
  and _59247_ (_07770_, _07769_, _07766_);
  and _59248_ (_07771_, _07770_, _07765_);
  and _59249_ (_07772_, _05884_, _05248_);
  or _59250_ (_07773_, _07772_, _06829_);
  and _59251_ (_07774_, _07773_, _03600_);
  or _59252_ (_07775_, _07774_, _03780_);
  or _59253_ (_07776_, _07775_, _07771_);
  not _59254_ (_07777_, _03622_);
  not _59255_ (_07778_, _03780_);
  and _59256_ (_07779_, _06378_, _05248_);
  or _59257_ (_07780_, _07779_, _06829_);
  or _59258_ (_07781_, _07780_, _07778_);
  and _59259_ (_07782_, _07781_, _07777_);
  and _59260_ (_07783_, _07782_, _07776_);
  or _59261_ (_07784_, _06829_, _05310_);
  and _59262_ (_07785_, _07768_, _03622_);
  and _59263_ (_07786_, _07785_, _07784_);
  or _59264_ (_07787_, _07786_, _07783_);
  and _59265_ (_07788_, _07787_, _06828_);
  and _59266_ (_07789_, _06849_, _03790_);
  and _59267_ (_07790_, _07789_, _07784_);
  or _59268_ (_07791_, _07790_, _03624_);
  or _59269_ (_07792_, _07791_, _07788_);
  not _59270_ (_07793_, _03785_);
  nor _59271_ (_07794_, _05882_, _06830_);
  not _59272_ (_07795_, _03624_);
  or _59273_ (_07796_, _06829_, _07795_);
  or _59274_ (_07797_, _07796_, _07794_);
  and _59275_ (_07798_, _07797_, _07793_);
  and _59276_ (_07799_, _07798_, _07792_);
  nor _59277_ (_07800_, _06377_, _06830_);
  or _59278_ (_07801_, _07800_, _06829_);
  and _59279_ (_07802_, _07801_, _03785_);
  or _59280_ (_07803_, _07802_, _03815_);
  or _59281_ (_07804_, _07803_, _07799_);
  or _59282_ (_07805_, _06846_, _04246_);
  and _59283_ (_07806_, _07805_, _03823_);
  and _59284_ (_07807_, _07806_, _07804_);
  and _59285_ (_07808_, _06843_, _03453_);
  or _59286_ (_07809_, _07808_, _03447_);
  or _59287_ (_07810_, _07809_, _07807_);
  and _59288_ (_07811_, _05831_, _05248_);
  or _59289_ (_07812_, _06829_, _03514_);
  or _59290_ (_07813_, _07812_, _07811_);
  and _59291_ (_07814_, _07813_, _43000_);
  and _59292_ (_07815_, _07814_, _07810_);
  or _59293_ (_07816_, _07815_, _06827_);
  and _59294_ (_40566_, _07816_, _41806_);
  nor _59295_ (_07817_, _43000_, _06075_);
  not _59296_ (_07818_, _05363_);
  and _59297_ (_07819_, _06769_, \oc8051_golden_model_1.PSW [7]);
  and _59298_ (_07820_, _07819_, _07818_);
  nor _59299_ (_07821_, _07820_, _05204_);
  and _59300_ (_07822_, _07820_, _05204_);
  nor _59301_ (_07823_, _07822_, _07821_);
  and _59302_ (_07824_, _07823_, \oc8051_golden_model_1.ACC [7]);
  nor _59303_ (_07825_, _07823_, \oc8051_golden_model_1.ACC [7]);
  nor _59304_ (_07826_, _07825_, _07824_);
  nor _59305_ (_07827_, _07819_, _07818_);
  nor _59306_ (_07828_, _07827_, _07820_);
  and _59307_ (_07829_, _07828_, \oc8051_golden_model_1.ACC [6]);
  nor _59308_ (_07830_, _07828_, _07433_);
  and _59309_ (_07831_, _07828_, _07433_);
  nor _59310_ (_07832_, _07831_, _07830_);
  and _59311_ (_07833_, _06765_, \oc8051_golden_model_1.PSW [7]);
  and _59312_ (_07834_, _07833_, _06766_);
  and _59313_ (_07835_, _07834_, _06763_);
  nor _59314_ (_07836_, _07835_, _06762_);
  nor _59315_ (_07837_, _07836_, _07819_);
  and _59316_ (_07838_, _07837_, \oc8051_golden_model_1.ACC [5]);
  nor _59317_ (_07839_, _07837_, _07478_);
  and _59318_ (_07840_, _07837_, _07478_);
  nor _59319_ (_07841_, _07840_, _07839_);
  nor _59320_ (_07842_, _07834_, _06763_);
  nor _59321_ (_07843_, _07842_, _07835_);
  and _59322_ (_07844_, _07843_, \oc8051_golden_model_1.ACC [4]);
  nor _59323_ (_07845_, _07843_, _07484_);
  and _59324_ (_07846_, _07843_, _07484_);
  nor _59325_ (_07847_, _07846_, _07845_);
  not _59326_ (_07848_, _05005_);
  not _59327_ (_07849_, _04875_);
  and _59328_ (_07850_, _06765_, _07849_);
  and _59329_ (_07851_, _07850_, \oc8051_golden_model_1.PSW [7]);
  nor _59330_ (_07852_, _07851_, _07848_);
  nor _59331_ (_07853_, _07852_, _07834_);
  and _59332_ (_07854_, _07853_, \oc8051_golden_model_1.ACC [3]);
  nor _59333_ (_07855_, _07853_, _07578_);
  and _59334_ (_07856_, _07853_, _07578_);
  nor _59335_ (_07857_, _07856_, _07855_);
  nor _59336_ (_07858_, _07833_, _07849_);
  nor _59337_ (_07859_, _07858_, _07851_);
  and _59338_ (_07860_, _07859_, \oc8051_golden_model_1.ACC [2]);
  nor _59339_ (_07861_, _07859_, _07584_);
  and _59340_ (_07862_, _07859_, _07584_);
  nor _59341_ (_07863_, _07862_, _07861_);
  and _59342_ (_07864_, _04620_, \oc8051_golden_model_1.PSW [7]);
  nor _59343_ (_07865_, _07864_, _06764_);
  nor _59344_ (_07866_, _07865_, _07833_);
  and _59345_ (_07867_, _07866_, \oc8051_golden_model_1.ACC [1]);
  and _59346_ (_07868_, _07866_, _03274_);
  nor _59347_ (_07869_, _07866_, _03274_);
  nor _59348_ (_07870_, _07869_, _07868_);
  not _59349_ (_07871_, \oc8051_golden_model_1.PSW [7]);
  and _59350_ (_07872_, _04634_, _07871_);
  nor _59351_ (_07873_, _07872_, _07864_);
  and _59352_ (_07874_, _07873_, \oc8051_golden_model_1.ACC [0]);
  not _59353_ (_07875_, _07874_);
  nor _59354_ (_07876_, _07875_, _07870_);
  nor _59355_ (_07877_, _07876_, _07867_);
  nor _59356_ (_07878_, _07877_, _07863_);
  nor _59357_ (_07879_, _07878_, _07860_);
  nor _59358_ (_07880_, _07879_, _07857_);
  nor _59359_ (_07881_, _07880_, _07854_);
  nor _59360_ (_07882_, _07881_, _07847_);
  nor _59361_ (_07883_, _07882_, _07844_);
  nor _59362_ (_07884_, _07883_, _07841_);
  nor _59363_ (_07885_, _07884_, _07838_);
  nor _59364_ (_07886_, _07885_, _07832_);
  nor _59365_ (_07887_, _07886_, _07829_);
  nor _59366_ (_07888_, _07887_, _07826_);
  and _59367_ (_07889_, _07887_, _07826_);
  nor _59368_ (_07890_, _07889_, _07888_);
  and _59369_ (_07891_, _03494_, _03187_);
  not _59370_ (_07892_, _07891_);
  and _59371_ (_07893_, _04066_, _03187_);
  and _59372_ (_07894_, _03493_, _03611_);
  nor _59373_ (_07895_, _07894_, _03489_);
  nor _59374_ (_07896_, _07895_, _04207_);
  nor _59375_ (_07897_, _07896_, _07893_);
  and _59376_ (_07898_, _07897_, _07892_);
  or _59377_ (_07899_, _07898_, _07890_);
  nor _59378_ (_07900_, _05254_, _06075_);
  and _59379_ (_07901_, _05884_, _05254_);
  nor _59380_ (_07902_, _07901_, _07900_);
  nand _59381_ (_07903_, _07902_, _03600_);
  and _59382_ (_07904_, _03603_, _03181_);
  not _59383_ (_07905_, _07904_);
  or _59384_ (_07906_, _06378_, _03779_);
  and _59385_ (_07907_, _07906_, _07905_);
  not _59386_ (_07908_, _05254_);
  nor _59387_ (_07909_, _07908_, _05204_);
  nor _59388_ (_07910_, _07909_, _07900_);
  nand _59389_ (_07911_, _07910_, _07390_);
  not _59390_ (_07912_, _03248_);
  and _59391_ (_07913_, _03603_, _03223_);
  not _59392_ (_07914_, _07913_);
  and _59393_ (_07915_, _05210_, \oc8051_golden_model_1.PSW [7]);
  and _59394_ (_07916_, _07915_, _05261_);
  and _59395_ (_07917_, _07916_, _05237_);
  and _59396_ (_07918_, _07917_, _05112_);
  nor _59397_ (_07919_, _07918_, _03446_);
  and _59398_ (_07920_, _07918_, _03446_);
  nor _59399_ (_07921_, _07920_, _07919_);
  and _59400_ (_07922_, _07921_, \oc8051_golden_model_1.ACC [7]);
  nor _59401_ (_07923_, _07921_, \oc8051_golden_model_1.ACC [7]);
  nor _59402_ (_07924_, _07923_, _07922_);
  nor _59403_ (_07925_, _07917_, _05112_);
  nor _59404_ (_07926_, _07925_, _07918_);
  nor _59405_ (_07927_, _07926_, _07433_);
  and _59406_ (_07928_, _07926_, _07433_);
  and _59407_ (_07929_, _07916_, _05218_);
  nor _59408_ (_07930_, _07929_, _05226_);
  nor _59409_ (_07931_, _07930_, _07917_);
  and _59410_ (_07932_, _07931_, _07478_);
  nor _59411_ (_07933_, _07931_, _07478_);
  nor _59412_ (_07934_, _07916_, _05218_);
  nor _59413_ (_07935_, _07934_, _07929_);
  nor _59414_ (_07936_, _07935_, _07484_);
  nor _59415_ (_07937_, _07936_, _07933_);
  nor _59416_ (_07938_, _07937_, _07932_);
  nor _59417_ (_07939_, _07933_, _07932_);
  and _59418_ (_07940_, _07935_, _07484_);
  nor _59419_ (_07941_, _07940_, _07936_);
  and _59420_ (_07942_, _07941_, _07939_);
  not _59421_ (_07943_, _07942_);
  nor _59422_ (_07944_, _05937_, _03756_);
  nor _59423_ (_07945_, _07944_, _07916_);
  nor _59424_ (_07946_, _07945_, _07578_);
  and _59425_ (_07947_, _07945_, _07578_);
  nor _59426_ (_07948_, _07947_, _07946_);
  nor _59427_ (_07949_, _07915_, _04800_);
  nor _59428_ (_07950_, _07949_, _05937_);
  nor _59429_ (_07951_, _07950_, _07584_);
  and _59430_ (_07952_, _07950_, _07584_);
  nor _59431_ (_07953_, _07952_, _07951_);
  and _59432_ (_07954_, _07953_, _07948_);
  nor _59433_ (_07955_, _04048_, _07871_);
  nor _59434_ (_07956_, _07955_, _03415_);
  nor _59435_ (_07957_, _07956_, _07915_);
  nor _59436_ (_07958_, _07957_, _03274_);
  and _59437_ (_07959_, _07957_, _03274_);
  and _59438_ (_07960_, _04048_, _07871_);
  nor _59439_ (_07961_, _07960_, _07955_);
  nor _59440_ (_07962_, _07961_, _03335_);
  not _59441_ (_07963_, _07962_);
  nor _59442_ (_07964_, _07963_, _07959_);
  nor _59443_ (_07965_, _07964_, _07958_);
  and _59444_ (_07966_, _07965_, _07954_);
  not _59445_ (_07967_, _07966_);
  and _59446_ (_07968_, _07952_, _07948_);
  nor _59447_ (_07969_, _07968_, _07947_);
  and _59448_ (_07970_, _07969_, _07967_);
  not _59449_ (_07971_, _07954_);
  nor _59450_ (_07972_, _07959_, _07958_);
  and _59451_ (_07973_, _07961_, _03335_);
  nor _59452_ (_07974_, _07962_, _07973_);
  nand _59453_ (_07975_, _07974_, _07972_);
  nor _59454_ (_07976_, _07975_, _07971_);
  nor _59455_ (_07977_, _07976_, _07970_);
  nor _59456_ (_07978_, _07977_, _07943_);
  nor _59457_ (_07979_, _07978_, _07938_);
  nor _59458_ (_07980_, _07979_, _07928_);
  or _59459_ (_07981_, _07980_, _07927_);
  or _59460_ (_07982_, _07981_, _07924_);
  nand _59461_ (_07983_, _07981_, _07924_);
  and _59462_ (_07984_, _07983_, _07982_);
  or _59463_ (_07985_, _07984_, _07914_);
  and _59464_ (_07986_, _06791_, \oc8051_golden_model_1.PSW [7]);
  nor _59465_ (_07987_, _07986_, _06410_);
  and _59466_ (_07988_, _07986_, _06410_);
  nor _59467_ (_07989_, _07988_, _07987_);
  and _59468_ (_07990_, _07989_, \oc8051_golden_model_1.ACC [7]);
  nor _59469_ (_07991_, _07989_, \oc8051_golden_model_1.ACC [7]);
  nor _59470_ (_07992_, _07991_, _07990_);
  not _59471_ (_07993_, _07992_);
  and _59472_ (_07994_, _06790_, \oc8051_golden_model_1.PSW [7]);
  nor _59473_ (_07995_, _07994_, _06455_);
  nor _59474_ (_07996_, _07995_, _07986_);
  nor _59475_ (_07997_, _07996_, _07433_);
  and _59476_ (_07998_, _07996_, _07433_);
  and _59477_ (_07999_, _06788_, _06730_);
  and _59478_ (_08000_, _07999_, \oc8051_golden_model_1.PSW [7]);
  nor _59479_ (_08001_, _08000_, _06684_);
  nor _59480_ (_08002_, _08001_, _07994_);
  and _59481_ (_08003_, _08002_, _07478_);
  nor _59482_ (_08004_, _08002_, _07478_);
  and _59483_ (_08005_, _06786_, \oc8051_golden_model_1.PSW [7]);
  and _59484_ (_08006_, _08005_, _06787_);
  nor _59485_ (_08007_, _08006_, _06730_);
  nor _59486_ (_08008_, _08007_, _08000_);
  nor _59487_ (_08009_, _08008_, _07484_);
  nor _59488_ (_08010_, _08009_, _08004_);
  nor _59489_ (_08011_, _08010_, _08003_);
  nor _59490_ (_08012_, _08004_, _08003_);
  and _59491_ (_08013_, _08008_, _07484_);
  nor _59492_ (_08014_, _08013_, _08009_);
  and _59493_ (_08015_, _08014_, _08012_);
  and _59494_ (_08016_, _06786_, _06637_);
  and _59495_ (_08017_, _08016_, \oc8051_golden_model_1.PSW [7]);
  nor _59496_ (_08018_, _08017_, _06592_);
  nor _59497_ (_08019_, _08018_, _08006_);
  nor _59498_ (_08020_, _08019_, _07578_);
  and _59499_ (_08021_, _08019_, _07578_);
  nor _59500_ (_08022_, _08021_, _08020_);
  nor _59501_ (_08023_, _08005_, _06637_);
  nor _59502_ (_08024_, _08023_, _08017_);
  nor _59503_ (_08025_, _08024_, _07584_);
  and _59504_ (_08026_, _08024_, _07584_);
  nor _59505_ (_08027_, _08026_, _08025_);
  and _59506_ (_08028_, _08027_, _08022_);
  and _59507_ (_08029_, _06546_, \oc8051_golden_model_1.PSW [7]);
  nor _59508_ (_08030_, _08029_, _06501_);
  nor _59509_ (_08031_, _08030_, _08005_);
  nor _59510_ (_08032_, _08031_, _03274_);
  and _59511_ (_08033_, _08031_, _03274_);
  nor _59512_ (_08034_, _06546_, \oc8051_golden_model_1.PSW [7]);
  nor _59513_ (_08035_, _08034_, _08029_);
  and _59514_ (_08036_, _08035_, _03335_);
  nor _59515_ (_08037_, _08036_, _08033_);
  or _59516_ (_08038_, _08037_, _08032_);
  and _59517_ (_08039_, _08038_, _08028_);
  and _59518_ (_08040_, _08025_, _08022_);
  or _59519_ (_08041_, _08040_, _08020_);
  nor _59520_ (_08042_, _08041_, _08039_);
  not _59521_ (_08043_, _08042_);
  and _59522_ (_08044_, _08043_, _08015_);
  nor _59523_ (_08045_, _08044_, _08011_);
  nor _59524_ (_08046_, _08045_, _07998_);
  or _59525_ (_08047_, _08046_, _07997_);
  and _59526_ (_08048_, _08047_, _07993_);
  nor _59527_ (_08049_, _08047_, _07993_);
  nor _59528_ (_08050_, _08049_, _08048_);
  nor _59529_ (_08051_, _03511_, _03247_);
  nand _59530_ (_08052_, _08051_, _08050_);
  and _59531_ (_08053_, _04058_, _03223_);
  not _59532_ (_08054_, _08053_);
  and _59533_ (_08055_, _04474_, _03223_);
  nor _59534_ (_08056_, _04750_, _03595_);
  nor _59535_ (_08057_, _08056_, _03247_);
  nor _59536_ (_08058_, _08057_, _08055_);
  and _59537_ (_08059_, _08058_, _08054_);
  not _59538_ (_08060_, _08059_);
  not _59539_ (_08061_, _04759_);
  nor _59540_ (_08062_, _04751_, _03985_);
  and _59541_ (_08063_, _08062_, _08061_);
  not _59542_ (_08064_, _08063_);
  nand _59543_ (_08065_, _08064_, _05204_);
  and _59544_ (_08066_, _03603_, _03725_);
  not _59545_ (_08067_, _08066_);
  or _59546_ (_08068_, _08067_, _06069_);
  and _59547_ (_08069_, _04081_, _03235_);
  nor _59548_ (_08070_, _07894_, _03595_);
  nor _59549_ (_08071_, _08070_, _03234_);
  nor _59550_ (_08072_, _08071_, _04067_);
  nor _59551_ (_08073_, _03511_, _03234_);
  nor _59552_ (_08074_, _08073_, _03726_);
  and _59553_ (_08075_, _08074_, _08072_);
  and _59554_ (_08076_, _03494_, _03725_);
  not _59555_ (_08077_, _08076_);
  and _59556_ (_08078_, _08077_, _08075_);
  not _59557_ (_08079_, _08078_);
  nand _59558_ (_08080_, _08079_, _05204_);
  nor _59559_ (_08081_, _04064_, _06075_);
  and _59560_ (_08082_, _04064_, _06075_);
  nor _59561_ (_08083_, _08082_, _08081_);
  nand _59562_ (_08084_, _08083_, _08078_);
  and _59563_ (_08085_, _08084_, _08080_);
  or _59564_ (_08086_, _08085_, _08066_);
  and _59565_ (_08087_, _08086_, _08069_);
  and _59566_ (_08088_, _08087_, _08068_);
  and _59567_ (_08089_, _03603_, _03609_);
  and _59568_ (_08090_, _05964_, _05254_);
  nor _59569_ (_08091_, _08090_, _07900_);
  nor _59570_ (_08092_, _08091_, _04081_);
  or _59571_ (_08093_, _08092_, _08089_);
  or _59572_ (_08094_, _08093_, _08088_);
  nor _59573_ (_08095_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor _59574_ (_08096_, _08095_, _07578_);
  and _59575_ (_08097_, _08096_, _07449_);
  and _59576_ (_08098_, _08097_, \oc8051_golden_model_1.ACC [6]);
  and _59577_ (_08099_, _08098_, \oc8051_golden_model_1.ACC [7]);
  nor _59578_ (_08100_, _08098_, \oc8051_golden_model_1.ACC [7]);
  nor _59579_ (_08101_, _08100_, _08099_);
  and _59580_ (_08102_, _08096_, \oc8051_golden_model_1.ACC [4]);
  nor _59581_ (_08103_, _08102_, \oc8051_golden_model_1.ACC [5]);
  nor _59582_ (_08104_, _08103_, _08097_);
  nor _59583_ (_08105_, _08097_, \oc8051_golden_model_1.ACC [6]);
  nor _59584_ (_08106_, _08105_, _08098_);
  nor _59585_ (_08107_, _08106_, _08104_);
  not _59586_ (_08108_, _08107_);
  and _59587_ (_08109_, _08108_, _08101_);
  nor _59588_ (_08110_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor _59589_ (_08111_, _08110_, _08107_);
  nor _59590_ (_08112_, _08111_, _08101_);
  nor _59591_ (_08113_, _08112_, _08109_);
  not _59592_ (_08114_, _08113_);
  nand _59593_ (_08115_, _08114_, _08089_);
  and _59594_ (_08116_, _08115_, _03730_);
  and _59595_ (_08117_, _08116_, _08094_);
  nor _59596_ (_08118_, _05903_, _06075_);
  and _59597_ (_08119_, _06095_, _05903_);
  nor _59598_ (_08120_, _08119_, _08118_);
  nor _59599_ (_08121_, _08120_, _04055_);
  nor _59600_ (_08122_, _07910_, _03996_);
  or _59601_ (_08123_, _08122_, _08064_);
  or _59602_ (_08124_, _08123_, _08121_);
  or _59603_ (_08125_, _08124_, _08117_);
  and _59604_ (_08126_, _08125_, _08065_);
  or _59605_ (_08127_, _08126_, _04443_);
  not _59606_ (_08128_, _04443_);
  or _59607_ (_08129_, _06069_, _08128_);
  and _59608_ (_08130_, _08129_, _03737_);
  and _59609_ (_08131_, _08130_, _08127_);
  and _59610_ (_08132_, _03603_, _03507_);
  nor _59611_ (_08133_, _06133_, _03737_);
  or _59612_ (_08134_, _08133_, _08132_);
  or _59613_ (_08135_, _08134_, _08131_);
  nand _59614_ (_08136_, _08132_, _07578_);
  and _59615_ (_08137_, _08136_, _08135_);
  or _59616_ (_08138_, _08137_, _03714_);
  and _59617_ (_08139_, _05952_, _05903_);
  nor _59618_ (_08140_, _08139_, _08118_);
  nand _59619_ (_08141_, _08140_, _03714_);
  and _59620_ (_08142_, _08141_, _06840_);
  and _59621_ (_08143_, _08142_, _08138_);
  and _59622_ (_08144_, _08119_, _06138_);
  nor _59623_ (_08145_, _08144_, _08118_);
  nor _59624_ (_08146_, _08145_, _06840_);
  or _59625_ (_08147_, _08146_, _06869_);
  or _59626_ (_08148_, _08147_, _08143_);
  nor _59627_ (_08149_, _07348_, _07346_);
  nor _59628_ (_08150_, _08149_, _07349_);
  or _59629_ (_08151_, _08150_, _06875_);
  and _59630_ (_08152_, _08151_, _08148_);
  or _59631_ (_08153_, _08152_, _08060_);
  not _59632_ (_08154_, _07826_);
  nor _59633_ (_08155_, _07845_, _07839_);
  nor _59634_ (_08156_, _08155_, _07840_);
  and _59635_ (_08157_, _07847_, _07841_);
  not _59636_ (_08158_, _08157_);
  and _59637_ (_08159_, _07863_, _07857_);
  nor _59638_ (_08160_, _07873_, _03335_);
  not _59639_ (_08161_, _08160_);
  nor _59640_ (_08162_, _08161_, _07868_);
  nor _59641_ (_08163_, _08162_, _07869_);
  and _59642_ (_08164_, _08163_, _08159_);
  not _59643_ (_08165_, _08164_);
  and _59644_ (_08166_, _07862_, _07857_);
  nor _59645_ (_08167_, _08166_, _07856_);
  and _59646_ (_08168_, _08167_, _08165_);
  and _59647_ (_08169_, _07873_, _03335_);
  nor _59648_ (_08170_, _08160_, _08169_);
  and _59649_ (_08171_, _08170_, _07870_);
  and _59650_ (_08172_, _08171_, _08159_);
  nor _59651_ (_08173_, _08172_, _08168_);
  nor _59652_ (_08174_, _08173_, _08158_);
  nor _59653_ (_08175_, _08174_, _08156_);
  nor _59654_ (_08176_, _08175_, _07831_);
  or _59655_ (_08177_, _08176_, _07830_);
  and _59656_ (_08178_, _08177_, _08154_);
  nor _59657_ (_08179_, _08177_, _08154_);
  or _59658_ (_08180_, _08179_, _08178_);
  or _59659_ (_08181_, _08180_, _08059_);
  and _59660_ (_08182_, _08181_, _08153_);
  or _59661_ (_08183_, _08182_, _08051_);
  and _59662_ (_08184_, _08183_, _03766_);
  and _59663_ (_08185_, _08184_, _08052_);
  nor _59664_ (_08186_, _07913_, _03761_);
  not _59665_ (_08187_, _08186_);
  and _59666_ (_08188_, _06133_, _06075_);
  nor _59667_ (_08189_, _06133_, _06075_);
  nor _59668_ (_08190_, _08189_, _08188_);
  not _59669_ (_08191_, _08190_);
  and _59670_ (_08192_, _05293_, \oc8051_golden_model_1.P0INREG [6]);
  and _59671_ (_08193_, _05266_, \oc8051_golden_model_1.P1INREG [6]);
  not _59672_ (_08194_, _08193_);
  and _59673_ (_08195_, _05235_, \oc8051_golden_model_1.P2INREG [6]);
  and _59674_ (_08196_, _05239_, \oc8051_golden_model_1.P3INREG [6]);
  nor _59675_ (_08197_, _08196_, _08195_);
  and _59676_ (_08198_, _08197_, _08194_);
  nand _59677_ (_08199_, _08198_, _05398_);
  nor _59678_ (_08200_, _08199_, _08192_);
  and _59679_ (_08201_, _08200_, _05391_);
  and _59680_ (_08202_, _08201_, _05381_);
  and _59681_ (_08203_, _08202_, _05364_);
  and _59682_ (_08204_, _08203_, \oc8051_golden_model_1.ACC [6]);
  nor _59683_ (_08205_, _08203_, \oc8051_golden_model_1.ACC [6]);
  nor _59684_ (_08206_, _08205_, _08204_);
  and _59685_ (_08207_, _05293_, \oc8051_golden_model_1.P0INREG [5]);
  and _59686_ (_08208_, _05266_, \oc8051_golden_model_1.P1INREG [5]);
  not _59687_ (_08209_, _08208_);
  and _59688_ (_08210_, _05235_, \oc8051_golden_model_1.P2INREG [5]);
  and _59689_ (_08211_, _05239_, \oc8051_golden_model_1.P3INREG [5]);
  nor _59690_ (_08212_, _08211_, _08210_);
  and _59691_ (_08213_, _08212_, _08209_);
  nand _59692_ (_08214_, _08213_, _05506_);
  nor _59693_ (_08215_, _08214_, _08207_);
  and _59694_ (_08216_, _08215_, _05497_);
  and _59695_ (_08217_, _08216_, _05491_);
  and _59696_ (_08218_, _08217_, _05470_);
  and _59697_ (_08219_, _08218_, \oc8051_golden_model_1.ACC [5]);
  nor _59698_ (_08220_, _08218_, \oc8051_golden_model_1.ACC [5]);
  and _59699_ (_08221_, _05266_, \oc8051_golden_model_1.P1INREG [4]);
  not _59700_ (_08222_, _08221_);
  not _59701_ (_08223_, _05799_);
  and _59702_ (_08224_, _05235_, \oc8051_golden_model_1.P2INREG [4]);
  and _59703_ (_08225_, _05239_, \oc8051_golden_model_1.P3INREG [4]);
  nor _59704_ (_08226_, _08225_, _08224_);
  and _59705_ (_08227_, _08226_, _08223_);
  and _59706_ (_08228_, _08227_, _08222_);
  and _59707_ (_08229_, _05293_, \oc8051_golden_model_1.P0INREG [4]);
  not _59708_ (_08230_, _08229_);
  and _59709_ (_08231_, _08230_, _05819_);
  and _59710_ (_08232_, _08231_, _05814_);
  and _59711_ (_08233_, _08232_, _08228_);
  and _59712_ (_08234_, _08233_, _05796_);
  and _59713_ (_08235_, _08234_, _05778_);
  and _59714_ (_08236_, _08235_, \oc8051_golden_model_1.ACC [4]);
  and _59715_ (_08237_, _05293_, \oc8051_golden_model_1.P0INREG [3]);
  and _59716_ (_08238_, _05266_, \oc8051_golden_model_1.P1INREG [3]);
  not _59717_ (_08239_, _08238_);
  and _59718_ (_08240_, _05235_, \oc8051_golden_model_1.P2INREG [3]);
  and _59719_ (_08241_, _05239_, \oc8051_golden_model_1.P3INREG [3]);
  nor _59720_ (_08242_, _08241_, _08240_);
  and _59721_ (_08243_, _08242_, _08239_);
  nand _59722_ (_08244_, _08243_, _05555_);
  nor _59723_ (_08245_, _08244_, _08237_);
  and _59724_ (_08246_, _08245_, _05546_);
  and _59725_ (_08247_, _08246_, _05540_);
  and _59726_ (_08248_, _08247_, _05519_);
  and _59727_ (_08249_, _08248_, \oc8051_golden_model_1.ACC [3]);
  nor _59728_ (_08250_, _08248_, \oc8051_golden_model_1.ACC [3]);
  and _59729_ (_08251_, _05235_, \oc8051_golden_model_1.P2INREG [2]);
  and _59730_ (_08252_, _05239_, \oc8051_golden_model_1.P3INREG [2]);
  nor _59731_ (_08253_, _08252_, _08251_);
  and _59732_ (_08254_, _05293_, \oc8051_golden_model_1.P0INREG [2]);
  and _59733_ (_08255_, _05266_, \oc8051_golden_model_1.P1INREG [2]);
  nor _59734_ (_08256_, _08255_, _08254_);
  and _59735_ (_08257_, _08256_, _08253_);
  and _59736_ (_08258_, _08257_, _05674_);
  and _59737_ (_08259_, _08258_, _05715_);
  and _59738_ (_08260_, _08259_, _05668_);
  and _59739_ (_08261_, _08260_, \oc8051_golden_model_1.ACC [2]);
  and _59740_ (_08262_, _05235_, \oc8051_golden_model_1.P2INREG [1]);
  and _59741_ (_08263_, _05239_, \oc8051_golden_model_1.P3INREG [1]);
  nor _59742_ (_08264_, _08263_, _08262_);
  and _59743_ (_08265_, _05293_, \oc8051_golden_model_1.P0INREG [1]);
  and _59744_ (_08266_, _05266_, \oc8051_golden_model_1.P1INREG [1]);
  nor _59745_ (_08267_, _08266_, _08265_);
  and _59746_ (_08268_, _08267_, _08264_);
  and _59747_ (_08269_, _08268_, _05574_);
  and _59748_ (_08270_, _08269_, _05615_);
  and _59749_ (_08271_, _08270_, _05568_);
  and _59750_ (_08272_, _08271_, \oc8051_golden_model_1.ACC [1]);
  nor _59751_ (_08273_, _08271_, \oc8051_golden_model_1.ACC [1]);
  and _59752_ (_08274_, _05293_, \oc8051_golden_model_1.P0INREG [0]);
  and _59753_ (_08275_, _05266_, \oc8051_golden_model_1.P1INREG [0]);
  not _59754_ (_08276_, _08275_);
  and _59755_ (_08277_, _05235_, \oc8051_golden_model_1.P2INREG [0]);
  and _59756_ (_08278_, _05239_, \oc8051_golden_model_1.P3INREG [0]);
  nor _59757_ (_08279_, _08278_, _08277_);
  and _59758_ (_08280_, _08279_, _08276_);
  nand _59759_ (_08281_, _08280_, _05655_);
  nor _59760_ (_08282_, _08281_, _08274_);
  and _59761_ (_08283_, _08282_, _05646_);
  and _59762_ (_08284_, _08283_, _05640_);
  and _59763_ (_08285_, _08284_, _05619_);
  nor _59764_ (_08286_, _08285_, \oc8051_golden_model_1.ACC [0]);
  nor _59765_ (_08287_, _08286_, _08273_);
  or _59766_ (_08288_, _08287_, _08272_);
  nor _59767_ (_08289_, _08260_, \oc8051_golden_model_1.ACC [2]);
  nor _59768_ (_08290_, _08289_, _08261_);
  and _59769_ (_08291_, _08290_, _08288_);
  nor _59770_ (_08292_, _08291_, _08261_);
  nor _59771_ (_08293_, _08292_, _08250_);
  or _59772_ (_08294_, _08293_, _08249_);
  nor _59773_ (_08295_, _08235_, \oc8051_golden_model_1.ACC [4]);
  nor _59774_ (_08296_, _08295_, _08236_);
  and _59775_ (_08297_, _08296_, _08294_);
  nor _59776_ (_08298_, _08297_, _08236_);
  nor _59777_ (_08299_, _08298_, _08220_);
  or _59778_ (_08300_, _08299_, _08219_);
  and _59779_ (_08301_, _08300_, _08206_);
  nor _59780_ (_08302_, _08301_, _08204_);
  and _59781_ (_08303_, _08302_, _08191_);
  nor _59782_ (_08304_, _08302_, _08191_);
  nor _59783_ (_08305_, _08304_, _08303_);
  nor _59784_ (_08306_, _08300_, _08206_);
  nor _59785_ (_08307_, _08306_, _08301_);
  nor _59786_ (_08308_, _08219_, _08220_);
  nor _59787_ (_08309_, _08308_, _08298_);
  and _59788_ (_08310_, _08308_, _08298_);
  or _59789_ (_08311_, _08310_, _08309_);
  nor _59790_ (_08312_, _08296_, _08294_);
  nor _59791_ (_08313_, _08312_, _08297_);
  nor _59792_ (_08314_, _08249_, _08250_);
  and _59793_ (_08315_, _08314_, _08290_);
  nor _59794_ (_08316_, _08272_, _08273_);
  and _59795_ (_08317_, _08285_, \oc8051_golden_model_1.ACC [0]);
  nor _59796_ (_08318_, _08317_, _08286_);
  and _59797_ (_08319_, _08318_, _08316_);
  and _59798_ (_08320_, _08319_, _08315_);
  and _59799_ (_08321_, _08320_, \oc8051_golden_model_1.PSW [7]);
  not _59800_ (_08322_, _08321_);
  nor _59801_ (_08323_, _08322_, _08313_);
  not _59802_ (_08324_, _08323_);
  nor _59803_ (_08325_, _08324_, _08311_);
  not _59804_ (_08326_, _08325_);
  nor _59805_ (_08327_, _08326_, _08307_);
  nor _59806_ (_08328_, _08327_, _08305_);
  and _59807_ (_08329_, _08327_, _08305_);
  nor _59808_ (_08330_, _08329_, _08328_);
  nand _59809_ (_08331_, _08330_, _07914_);
  and _59810_ (_08332_, _08331_, _08187_);
  or _59811_ (_08333_, _08332_, _08185_);
  and _59812_ (_08334_, _08333_, _07985_);
  or _59813_ (_08335_, _08334_, _07912_);
  nand _59814_ (_08336_, _03446_, _07912_);
  and _59815_ (_08337_, _08336_, _03710_);
  and _59816_ (_08338_, _08337_, _08335_);
  not _59817_ (_08339_, _05903_);
  nor _59818_ (_08340_, _05938_, _08339_);
  nor _59819_ (_08341_, _08340_, _08118_);
  nor _59820_ (_08342_, _08341_, _03710_);
  or _59821_ (_08343_, _08342_, _07390_);
  or _59822_ (_08344_, _08343_, _08338_);
  and _59823_ (_08345_, _08344_, _07911_);
  or _59824_ (_08346_, _08345_, _04481_);
  and _59825_ (_08347_, _06069_, _05254_);
  nor _59826_ (_08348_, _08347_, _07900_);
  nand _59827_ (_08349_, _08348_, _04481_);
  and _59828_ (_08350_, _08349_, _03589_);
  and _59829_ (_08351_, _08350_, _08346_);
  nor _59830_ (_08352_, _06363_, _07908_);
  nor _59831_ (_08353_, _08352_, _07900_);
  nor _59832_ (_08354_, _08353_, _03589_);
  or _59833_ (_08355_, _08354_, _07405_);
  or _59834_ (_08356_, _08355_, _08351_);
  or _59835_ (_08357_, _07424_, _07411_);
  and _59836_ (_08358_, _08357_, _08356_);
  or _59837_ (_08359_, _08358_, _03216_);
  nand _59838_ (_08360_, _03446_, _03216_);
  and _59839_ (_08361_, _08360_, _08359_);
  or _59840_ (_08362_, _08361_, _03601_);
  and _59841_ (_08363_, _03603_, _03176_);
  not _59842_ (_08364_, _08363_);
  and _59843_ (_08365_, _06171_, _05254_);
  nor _59844_ (_08366_, _08365_, _07900_);
  nand _59845_ (_08367_, _08366_, _03601_);
  and _59846_ (_08368_, _08367_, _08364_);
  and _59847_ (_08369_, _08368_, _08362_);
  nor _59848_ (_08370_, _08364_, _03446_);
  and _59849_ (_08371_, _04474_, _03181_);
  or _59850_ (_08372_, _08371_, _08370_);
  or _59851_ (_08373_, _08372_, _08369_);
  and _59852_ (_08374_, _05204_, _06075_);
  nor _59853_ (_08375_, _05204_, _06075_);
  nor _59854_ (_08376_, _08375_, _08374_);
  not _59855_ (_08377_, _08371_);
  or _59856_ (_08378_, _08377_, _08376_);
  not _59857_ (_08379_, _04181_);
  and _59858_ (_08380_, _03595_, _03181_);
  and _59859_ (_08381_, _07894_, _03181_);
  nor _59860_ (_08382_, _08381_, _08380_);
  and _59861_ (_08383_, _08382_, _08379_);
  and _59862_ (_08384_, _08383_, _08378_);
  and _59863_ (_08385_, _08384_, _08373_);
  and _59864_ (_08386_, _03494_, _03181_);
  nor _59865_ (_08387_, _08386_, _04181_);
  nand _59866_ (_08388_, _08387_, _08382_);
  or _59867_ (_08389_, _08386_, _08376_);
  and _59868_ (_08390_, _08389_, _08388_);
  or _59869_ (_08391_, _08390_, _08385_);
  nor _59870_ (_08392_, _03511_, _04175_);
  not _59871_ (_08393_, _08392_);
  not _59872_ (_08394_, _08386_);
  or _59873_ (_08395_, _08394_, _08376_);
  and _59874_ (_08396_, _08395_, _08393_);
  and _59875_ (_08397_, _08396_, _08391_);
  nor _59876_ (_08398_, _06069_, \oc8051_golden_model_1.ACC [7]);
  and _59877_ (_08399_, _06069_, \oc8051_golden_model_1.ACC [7]);
  nor _59878_ (_08400_, _08399_, _08398_);
  and _59879_ (_08401_, _08392_, _08400_);
  or _59880_ (_08402_, _08401_, _03778_);
  or _59881_ (_08403_, _08402_, _08397_);
  and _59882_ (_08404_, _08403_, _07907_);
  nor _59883_ (_08405_, _03446_, _06075_);
  and _59884_ (_08406_, _03446_, _06075_);
  nor _59885_ (_08407_, _08406_, _08405_);
  and _59886_ (_08408_, _08407_, _07904_);
  or _59887_ (_08409_, _08408_, _03600_);
  or _59888_ (_08410_, _08409_, _08404_);
  and _59889_ (_08411_, _08410_, _07903_);
  or _59890_ (_08412_, _08411_, _03780_);
  or _59891_ (_08413_, _07900_, _07778_);
  not _59892_ (_08414_, _04198_);
  and _59893_ (_08415_, _03489_, _03191_);
  nor _59894_ (_08416_, _08415_, _04315_);
  and _59895_ (_08417_, _08416_, _08414_);
  and _59896_ (_08418_, _08417_, _08413_);
  and _59897_ (_08419_, _08418_, _08412_);
  nor _59898_ (_08420_, _03511_, _04193_);
  not _59899_ (_08421_, _08417_);
  and _59900_ (_08422_, _08421_, _08375_);
  or _59901_ (_08423_, _08422_, _08420_);
  or _59902_ (_08424_, _08423_, _08419_);
  not _59903_ (_08425_, _08420_);
  or _59904_ (_08426_, _08425_, _08399_);
  and _59905_ (_08427_, _08426_, _03789_);
  and _59906_ (_08428_, _08427_, _08424_);
  and _59907_ (_08429_, _03603_, _03191_);
  nor _59908_ (_08430_, _08429_, _03788_);
  not _59909_ (_08431_, _08430_);
  or _59910_ (_08432_, _08429_, _06376_);
  and _59911_ (_08433_, _08432_, _08431_);
  or _59912_ (_08434_, _08433_, _08428_);
  not _59913_ (_08435_, _08429_);
  or _59914_ (_08436_, _08435_, _08405_);
  and _59915_ (_08437_, _08436_, _07777_);
  and _59916_ (_08438_, _08437_, _08434_);
  or _59917_ (_08439_, _08366_, _06377_);
  nor _59918_ (_08440_, _08439_, _07777_);
  and _59919_ (_08441_, _03489_, _03200_);
  or _59920_ (_08442_, _08441_, _08440_);
  or _59921_ (_08443_, _08442_, _08438_);
  and _59922_ (_08444_, _03493_, _03200_);
  nor _59923_ (_08445_, _08444_, _08374_);
  and _59924_ (_08446_, _03200_, _02962_);
  not _59925_ (_08447_, _08446_);
  or _59926_ (_08448_, _08447_, _08445_);
  and _59927_ (_08449_, _08448_, _08443_);
  nor _59928_ (_08450_, _03511_, _04190_);
  not _59929_ (_08451_, _08374_);
  and _59930_ (_08452_, _08444_, _08451_);
  or _59931_ (_08453_, _08452_, _08450_);
  or _59932_ (_08454_, _08453_, _08449_);
  nand _59933_ (_08455_, _08450_, _08398_);
  and _59934_ (_08456_, _08455_, _03784_);
  and _59935_ (_08457_, _08456_, _08454_);
  and _59936_ (_08458_, _03603_, _03200_);
  nor _59937_ (_08459_, _08458_, _03783_);
  not _59938_ (_08460_, _08459_);
  not _59939_ (_08461_, _08458_);
  nand _59940_ (_08462_, _08461_, _06377_);
  and _59941_ (_08463_, _08462_, _08460_);
  or _59942_ (_08464_, _08463_, _08457_);
  nand _59943_ (_08465_, _08458_, _08406_);
  and _59944_ (_08466_, _08465_, _07795_);
  and _59945_ (_08467_, _08466_, _08464_);
  not _59946_ (_08468_, _07898_);
  nor _59947_ (_08469_, _05882_, _07908_);
  nor _59948_ (_08470_, _08469_, _07900_);
  nor _59949_ (_08471_, _08470_, _07795_);
  or _59950_ (_08472_, _08471_, _08468_);
  or _59951_ (_08473_, _08472_, _08467_);
  and _59952_ (_08474_, _08473_, _07899_);
  nor _59953_ (_08475_, _03511_, _04207_);
  or _59954_ (_08476_, _08475_, _08474_);
  not _59955_ (_08477_, _08475_);
  and _59956_ (_08478_, _07996_, \oc8051_golden_model_1.ACC [6]);
  nor _59957_ (_08479_, _07997_, _07998_);
  and _59958_ (_08480_, _08002_, \oc8051_golden_model_1.ACC [5]);
  and _59959_ (_08481_, _08008_, \oc8051_golden_model_1.ACC [4]);
  and _59960_ (_08482_, _08019_, \oc8051_golden_model_1.ACC [3]);
  and _59961_ (_08483_, _08024_, \oc8051_golden_model_1.ACC [2]);
  and _59962_ (_08484_, _08031_, \oc8051_golden_model_1.ACC [1]);
  nor _59963_ (_08485_, _08032_, _08033_);
  and _59964_ (_08486_, _08035_, \oc8051_golden_model_1.ACC [0]);
  not _59965_ (_08487_, _08486_);
  nor _59966_ (_08488_, _08487_, _08485_);
  nor _59967_ (_08489_, _08488_, _08484_);
  nor _59968_ (_08490_, _08489_, _08027_);
  nor _59969_ (_08491_, _08490_, _08483_);
  nor _59970_ (_08492_, _08491_, _08022_);
  nor _59971_ (_08493_, _08492_, _08482_);
  nor _59972_ (_08494_, _08493_, _08014_);
  nor _59973_ (_08495_, _08494_, _08481_);
  nor _59974_ (_08496_, _08495_, _08012_);
  nor _59975_ (_08497_, _08496_, _08480_);
  nor _59976_ (_08498_, _08497_, _08479_);
  nor _59977_ (_08499_, _08498_, _08478_);
  nor _59978_ (_08500_, _08499_, _07992_);
  and _59979_ (_08501_, _08499_, _07992_);
  nor _59980_ (_08502_, _08501_, _08500_);
  or _59981_ (_08503_, _08502_, _08477_);
  and _59982_ (_08504_, _08503_, _03777_);
  and _59983_ (_08505_, _08504_, _08476_);
  and _59984_ (_08506_, _03603_, _03187_);
  nor _59985_ (_08507_, _08506_, _03776_);
  not _59986_ (_08508_, _08507_);
  not _59987_ (_08509_, _08203_);
  not _59988_ (_08510_, _08248_);
  not _59989_ (_08511_, _08260_);
  not _59990_ (_08512_, _08271_);
  nor _59991_ (_08513_, _08285_, _07871_);
  and _59992_ (_08514_, _08513_, _08512_);
  and _59993_ (_08515_, _08514_, _08511_);
  and _59994_ (_08516_, _08515_, _08510_);
  nor _59995_ (_08517_, _08235_, _08218_);
  and _59996_ (_08518_, _08517_, _08516_);
  and _59997_ (_08519_, _08518_, _08509_);
  nor _59998_ (_08520_, _08519_, _06133_);
  and _59999_ (_08521_, _08519_, _06133_);
  nor _60000_ (_08522_, _08521_, _08520_);
  and _60001_ (_08523_, _08522_, \oc8051_golden_model_1.ACC [7]);
  nor _60002_ (_08524_, _08522_, \oc8051_golden_model_1.ACC [7]);
  nor _60003_ (_08525_, _08524_, _08523_);
  nor _60004_ (_08526_, _08518_, _08509_);
  nor _60005_ (_08527_, _08526_, _08519_);
  and _60006_ (_08528_, _08527_, \oc8051_golden_model_1.ACC [6]);
  and _60007_ (_08529_, _08527_, _07433_);
  nor _60008_ (_08530_, _08527_, _07433_);
  nor _60009_ (_08531_, _08530_, _08529_);
  not _60010_ (_08532_, _08218_);
  not _60011_ (_08533_, _08235_);
  and _60012_ (_08534_, _08516_, _08533_);
  nor _60013_ (_08535_, _08534_, _08532_);
  nor _60014_ (_08536_, _08535_, _08518_);
  and _60015_ (_08537_, _08536_, \oc8051_golden_model_1.ACC [5]);
  and _60016_ (_08538_, _08536_, _07478_);
  nor _60017_ (_08539_, _08536_, _07478_);
  nor _60018_ (_08540_, _08539_, _08538_);
  nor _60019_ (_08541_, _08516_, _08533_);
  nor _60020_ (_08542_, _08541_, _08534_);
  and _60021_ (_08543_, _08542_, \oc8051_golden_model_1.ACC [4]);
  nor _60022_ (_08544_, _08542_, _07484_);
  and _60023_ (_08545_, _08542_, _07484_);
  nor _60024_ (_08546_, _08545_, _08544_);
  nor _60025_ (_08547_, _08515_, _08510_);
  nor _60026_ (_08548_, _08547_, _08516_);
  and _60027_ (_08549_, _08548_, \oc8051_golden_model_1.ACC [3]);
  nor _60028_ (_08550_, _08548_, _07578_);
  and _60029_ (_08551_, _08548_, _07578_);
  nor _60030_ (_08552_, _08551_, _08550_);
  nor _60031_ (_08553_, _08514_, _08511_);
  nor _60032_ (_08554_, _08553_, _08515_);
  and _60033_ (_08555_, _08554_, \oc8051_golden_model_1.ACC [2]);
  nor _60034_ (_08556_, _08554_, _07584_);
  and _60035_ (_08557_, _08554_, _07584_);
  nor _60036_ (_08558_, _08557_, _08556_);
  nor _60037_ (_08559_, _08513_, _08512_);
  nor _60038_ (_08560_, _08559_, _08514_);
  and _60039_ (_08561_, _08560_, \oc8051_golden_model_1.ACC [1]);
  and _60040_ (_08562_, _08560_, _03274_);
  nor _60041_ (_08563_, _08560_, _03274_);
  nor _60042_ (_08564_, _08563_, _08562_);
  and _60043_ (_08565_, _08285_, _07871_);
  nor _60044_ (_08566_, _08565_, _08513_);
  and _60045_ (_08567_, _08566_, \oc8051_golden_model_1.ACC [0]);
  not _60046_ (_08568_, _08567_);
  nor _60047_ (_08569_, _08568_, _08564_);
  nor _60048_ (_08570_, _08569_, _08561_);
  nor _60049_ (_08571_, _08570_, _08558_);
  nor _60050_ (_08572_, _08571_, _08555_);
  nor _60051_ (_08573_, _08572_, _08552_);
  nor _60052_ (_08574_, _08573_, _08549_);
  nor _60053_ (_08575_, _08574_, _08546_);
  nor _60054_ (_08576_, _08575_, _08543_);
  nor _60055_ (_08577_, _08576_, _08540_);
  nor _60056_ (_08578_, _08577_, _08537_);
  nor _60057_ (_08579_, _08578_, _08531_);
  nor _60058_ (_08580_, _08579_, _08528_);
  nor _60059_ (_08581_, _08580_, _08525_);
  and _60060_ (_08582_, _08580_, _08525_);
  nor _60061_ (_08583_, _08582_, _08581_);
  or _60062_ (_08584_, _08583_, _08506_);
  and _60063_ (_08585_, _08584_, _08508_);
  or _60064_ (_08586_, _08585_, _08505_);
  and _60065_ (_08587_, _03599_, _03187_);
  not _60066_ (_08588_, _08587_);
  not _60067_ (_08589_, _08506_);
  and _60068_ (_08590_, _07926_, \oc8051_golden_model_1.ACC [6]);
  nor _60069_ (_08591_, _07927_, _07928_);
  and _60070_ (_08592_, _07931_, \oc8051_golden_model_1.ACC [5]);
  and _60071_ (_08593_, _07935_, \oc8051_golden_model_1.ACC [4]);
  and _60072_ (_08594_, _07945_, \oc8051_golden_model_1.ACC [3]);
  and _60073_ (_08595_, _07950_, \oc8051_golden_model_1.ACC [2]);
  and _60074_ (_08596_, _07957_, \oc8051_golden_model_1.ACC [1]);
  and _60075_ (_08597_, _07961_, \oc8051_golden_model_1.ACC [0]);
  not _60076_ (_08598_, _08597_);
  nor _60077_ (_08599_, _08598_, _07972_);
  nor _60078_ (_08600_, _08599_, _08596_);
  nor _60079_ (_08601_, _08600_, _07953_);
  nor _60080_ (_08602_, _08601_, _08595_);
  nor _60081_ (_08603_, _08602_, _07948_);
  nor _60082_ (_08604_, _08603_, _08594_);
  nor _60083_ (_08605_, _08604_, _07941_);
  nor _60084_ (_08606_, _08605_, _08593_);
  nor _60085_ (_08607_, _08606_, _07939_);
  nor _60086_ (_08608_, _08607_, _08592_);
  nor _60087_ (_08609_, _08608_, _08591_);
  nor _60088_ (_08610_, _08609_, _08590_);
  nor _60089_ (_08611_, _08610_, _07924_);
  and _60090_ (_08612_, _08610_, _07924_);
  nor _60091_ (_08613_, _08612_, _08611_);
  or _60092_ (_08614_, _08613_, _08589_);
  and _60093_ (_08615_, _08614_, _08588_);
  and _60094_ (_08616_, _08615_, _08586_);
  nand _60095_ (_08617_, _03202_, _02962_);
  not _60096_ (_08618_, _08617_);
  and _60097_ (_08619_, _08587_, \oc8051_golden_model_1.ACC [6]);
  nor _60098_ (_08620_, _03511_, _03949_);
  or _60099_ (_08621_, _08620_, _08619_);
  or _60100_ (_08622_, _08621_, _08618_);
  or _60101_ (_08623_, _08622_, _08616_);
  not _60102_ (_08624_, _08620_);
  and _60103_ (_08625_, _06455_, \oc8051_golden_model_1.ACC [6]);
  nor _60104_ (_08626_, _06455_, \oc8051_golden_model_1.ACC [6]);
  nor _60105_ (_08627_, _08626_, _08625_);
  and _60106_ (_08628_, _06684_, \oc8051_golden_model_1.ACC [5]);
  nor _60107_ (_08629_, _06684_, \oc8051_golden_model_1.ACC [5]);
  nor _60108_ (_08630_, _08629_, _08628_);
  not _60109_ (_08631_, _08630_);
  and _60110_ (_08632_, _06730_, \oc8051_golden_model_1.ACC [4]);
  nor _60111_ (_08633_, _06730_, \oc8051_golden_model_1.ACC [4]);
  nor _60112_ (_08634_, _08633_, _08632_);
  and _60113_ (_08635_, _06592_, \oc8051_golden_model_1.ACC [3]);
  nor _60114_ (_08636_, _06591_, _06569_);
  and _60115_ (_08637_, _08636_, _07578_);
  and _60116_ (_08638_, _06637_, \oc8051_golden_model_1.ACC [2]);
  nor _60117_ (_08639_, _06637_, \oc8051_golden_model_1.ACC [2]);
  nor _60118_ (_08640_, _08639_, _08638_);
  not _60119_ (_08641_, _08640_);
  and _60120_ (_08642_, _06501_, \oc8051_golden_model_1.ACC [1]);
  nor _60121_ (_08643_, _06501_, \oc8051_golden_model_1.ACC [1]);
  nor _60122_ (_08644_, _08643_, _08642_);
  and _60123_ (_08645_, _06546_, \oc8051_golden_model_1.ACC [0]);
  and _60124_ (_08646_, _08645_, _08644_);
  nor _60125_ (_08647_, _08646_, _08642_);
  nor _60126_ (_08648_, _08647_, _08641_);
  nor _60127_ (_08649_, _08648_, _08638_);
  nor _60128_ (_08650_, _08649_, _08637_);
  or _60129_ (_08651_, _08650_, _08635_);
  and _60130_ (_08652_, _08651_, _08634_);
  nor _60131_ (_08653_, _08652_, _08632_);
  nor _60132_ (_08654_, _08653_, _08631_);
  or _60133_ (_08655_, _08654_, _08628_);
  and _60134_ (_08656_, _08655_, _08627_);
  nor _60135_ (_08657_, _08656_, _08625_);
  nor _60136_ (_08658_, _08657_, _08400_);
  and _60137_ (_08659_, _08657_, _08400_);
  or _60138_ (_08660_, _08659_, _08658_);
  or _60139_ (_08661_, _08660_, _08624_);
  nor _60140_ (_08662_, _05363_, _07433_);
  and _60141_ (_08663_, _05363_, _07433_);
  nor _60142_ (_08664_, _08663_, _08662_);
  nor _60143_ (_08665_, _05469_, _07478_);
  and _60144_ (_08666_, _05469_, _07478_);
  nor _60145_ (_08667_, _05777_, _07484_);
  and _60146_ (_08668_, _05777_, _07484_);
  nor _60147_ (_08669_, _08668_, _08667_);
  not _60148_ (_08670_, _08669_);
  nor _60149_ (_08671_, _05005_, _07578_);
  not _60150_ (_08672_, _08671_);
  and _60151_ (_08673_, _05005_, _07578_);
  nor _60152_ (_08674_, _04875_, _07584_);
  and _60153_ (_08675_, _04875_, _07584_);
  nor _60154_ (_08676_, _08675_, _08674_);
  not _60155_ (_08677_, _08676_);
  and _60156_ (_08678_, _06764_, \oc8051_golden_model_1.ACC [1]);
  and _60157_ (_08679_, _04406_, _03274_);
  nor _60158_ (_08680_, _08679_, _08678_);
  and _60159_ (_08681_, _04620_, \oc8051_golden_model_1.ACC [0]);
  and _60160_ (_08682_, _08681_, _08680_);
  nor _60161_ (_08683_, _08682_, _08678_);
  nor _60162_ (_08684_, _08683_, _08677_);
  nor _60163_ (_08685_, _08684_, _08674_);
  or _60164_ (_08686_, _08685_, _08673_);
  and _60165_ (_08687_, _08686_, _08672_);
  nor _60166_ (_08688_, _08687_, _08670_);
  nor _60167_ (_08689_, _08688_, _08667_);
  nor _60168_ (_08690_, _08689_, _08666_);
  or _60169_ (_08691_, _08690_, _08665_);
  and _60170_ (_08692_, _08691_, _08664_);
  nor _60171_ (_08693_, _08692_, _08662_);
  nor _60172_ (_08694_, _08693_, _08376_);
  and _60173_ (_08695_, _08693_, _08376_);
  or _60174_ (_08696_, _08695_, _08694_);
  or _60175_ (_08697_, _08696_, _08617_);
  and _60176_ (_08698_, _08697_, _03518_);
  and _60177_ (_08699_, _08698_, _08661_);
  and _60178_ (_08700_, _08699_, _08623_);
  and _60179_ (_08701_, _03603_, _03202_);
  nor _60180_ (_08702_, _08701_, _03517_);
  not _60181_ (_08703_, _08702_);
  nor _60182_ (_08704_, _08203_, _07433_);
  nor _60183_ (_08705_, _08218_, _07478_);
  nor _60184_ (_08706_, _08235_, _07484_);
  not _60185_ (_08707_, _08296_);
  nor _60186_ (_08708_, _08260_, _07584_);
  nor _60187_ (_08709_, _08271_, _03274_);
  nor _60188_ (_08710_, _08285_, _03335_);
  not _60189_ (_08711_, _08710_);
  nor _60190_ (_08712_, _08711_, _08316_);
  nor _60191_ (_08713_, _08712_, _08709_);
  nor _60192_ (_08714_, _08713_, _08290_);
  nor _60193_ (_08715_, _08714_, _08708_);
  nor _60194_ (_08716_, _08715_, _08248_);
  or _60195_ (_08717_, _08716_, \oc8051_golden_model_1.ACC [3]);
  nand _60196_ (_08718_, _08715_, _08248_);
  and _60197_ (_08719_, _08718_, _08717_);
  and _60198_ (_08720_, _08719_, _08707_);
  nor _60199_ (_08721_, _08720_, _08706_);
  nor _60200_ (_08722_, _08721_, _08308_);
  nor _60201_ (_08723_, _08722_, _08705_);
  nor _60202_ (_08724_, _08723_, _08206_);
  nor _60203_ (_08725_, _08724_, _08704_);
  nor _60204_ (_08726_, _08725_, _08190_);
  and _60205_ (_08727_, _08725_, _08190_);
  or _60206_ (_08728_, _08727_, _08726_);
  or _60207_ (_08729_, _08728_, _08701_);
  and _60208_ (_08730_, _08729_, _08703_);
  or _60209_ (_08731_, _08730_, _08700_);
  and _60210_ (_08732_, _03599_, _03202_);
  not _60211_ (_08733_, _08732_);
  not _60212_ (_08734_, _08701_);
  nor _60213_ (_08735_, _03549_, _07433_);
  and _60214_ (_08736_, _03549_, _07433_);
  or _60215_ (_08737_, _08736_, _08735_);
  not _60216_ (_08738_, _08737_);
  nor _60217_ (_08739_, _03860_, _07478_);
  and _60218_ (_08740_, _03860_, _07478_);
  nor _60219_ (_08741_, _03486_, _07484_);
  and _60220_ (_08742_, _03486_, _07484_);
  nor _60221_ (_08743_, _08742_, _08741_);
  nor _60222_ (_08744_, _03581_, _07578_);
  and _60223_ (_08745_, _03581_, _07578_);
  nor _60224_ (_08746_, _03904_, _07584_);
  and _60225_ (_08747_, _03904_, _07584_);
  nor _60226_ (_08748_, _08747_, _08746_);
  not _60227_ (_08749_, _08748_);
  nor _60228_ (_08750_, _03414_, _03274_);
  nor _60229_ (_08751_, _04048_, _03335_);
  and _60230_ (_08752_, _03414_, _03274_);
  nor _60231_ (_08753_, _08752_, _08750_);
  and _60232_ (_08754_, _08753_, _08751_);
  nor _60233_ (_08755_, _08754_, _08750_);
  nor _60234_ (_08756_, _08755_, _08749_);
  nor _60235_ (_08757_, _08756_, _08746_);
  nor _60236_ (_08758_, _08757_, _08745_);
  or _60237_ (_08759_, _08758_, _08744_);
  and _60238_ (_08760_, _08759_, _08743_);
  nor _60239_ (_08761_, _08760_, _08741_);
  nor _60240_ (_08762_, _08761_, _08740_);
  or _60241_ (_08763_, _08762_, _08739_);
  and _60242_ (_08764_, _08763_, _08738_);
  nor _60243_ (_08765_, _08764_, _08735_);
  nor _60244_ (_08766_, _08765_, _08407_);
  and _60245_ (_08767_, _08765_, _08407_);
  or _60246_ (_08768_, _08767_, _08766_);
  or _60247_ (_08769_, _08768_, _08734_);
  and _60248_ (_08770_, _08769_, _08733_);
  and _60249_ (_08771_, _08770_, _08731_);
  and _60250_ (_08772_, _08732_, \oc8051_golden_model_1.ACC [6]);
  or _60251_ (_08773_, _08772_, _03815_);
  or _60252_ (_08774_, _08773_, _08771_);
  and _60253_ (_08775_, _03603_, _03197_);
  not _60254_ (_08776_, _08775_);
  nand _60255_ (_08777_, _08091_, _03815_);
  and _60256_ (_08778_, _08777_, _08776_);
  and _60257_ (_08779_, _08778_, _08774_);
  and _60258_ (_08780_, _03599_, _03197_);
  nor _60259_ (_08781_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and _60260_ (_08782_, _08781_, _07524_);
  and _60261_ (_08783_, _08782_, _07448_);
  and _60262_ (_08784_, _08783_, _07433_);
  nor _60263_ (_08785_, _08784_, _06075_);
  and _60264_ (_08786_, _08784_, _06075_);
  nor _60265_ (_08787_, _08786_, _08785_);
  not _60266_ (_08788_, _08787_);
  and _60267_ (_08789_, _08788_, _08775_);
  or _60268_ (_08790_, _08789_, _08780_);
  or _60269_ (_08791_, _08790_, _08779_);
  nand _60270_ (_08792_, _08780_, _07871_);
  and _60271_ (_08793_, _08792_, _03823_);
  and _60272_ (_08794_, _08793_, _08791_);
  nor _60273_ (_08795_, _08140_, _03823_);
  or _60274_ (_08796_, _08795_, _03447_);
  or _60275_ (_08797_, _08796_, _08794_);
  and _60276_ (_08798_, _03603_, _03195_);
  not _60277_ (_08799_, _08798_);
  and _60278_ (_08800_, _05831_, _05254_);
  nor _60279_ (_08801_, _08800_, _07900_);
  nand _60280_ (_08802_, _08801_, _03447_);
  and _60281_ (_08803_, _08802_, _08799_);
  and _60282_ (_08804_, _08803_, _08797_);
  and _60283_ (_08805_, _03599_, _03195_);
  and _60284_ (_08806_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand _60285_ (_08807_, _08806_, _07525_);
  nor _60286_ (_08808_, _08807_, _07484_);
  and _60287_ (_08809_, _08808_, \oc8051_golden_model_1.ACC [5]);
  and _60288_ (_08810_, _08809_, \oc8051_golden_model_1.ACC [6]);
  nor _60289_ (_08811_, _08810_, \oc8051_golden_model_1.ACC [7]);
  and _60290_ (_08812_, _08810_, \oc8051_golden_model_1.ACC [7]);
  nor _60291_ (_08813_, _08812_, _08811_);
  and _60292_ (_08814_, _08813_, _08798_);
  or _60293_ (_08815_, _08814_, _08805_);
  or _60294_ (_08816_, _08815_, _08804_);
  nand _60295_ (_08817_, _08805_, _03335_);
  and _60296_ (_08818_, _08817_, _43000_);
  and _60297_ (_08819_, _08818_, _08816_);
  or _60298_ (_08820_, _08819_, _07817_);
  and _60299_ (_40567_, _08820_, _41806_);
  not _60300_ (_08821_, \oc8051_golden_model_1.DPL [7]);
  nor _60301_ (_08822_, _43000_, _08821_);
  nor _60302_ (_08823_, _05303_, _08821_);
  not _60303_ (_08824_, _05303_);
  nor _60304_ (_08825_, _06377_, _08824_);
  or _60305_ (_08826_, _08825_, _08823_);
  and _60306_ (_08827_, _08826_, _03785_);
  not _60307_ (_08828_, _03602_);
  nor _60308_ (_08829_, _08824_, _05204_);
  or _60309_ (_08830_, _08829_, _08823_);
  or _60310_ (_08831_, _08830_, _06838_);
  not _60311_ (_08832_, _03625_);
  and _60312_ (_08833_, _05964_, _05303_);
  or _60313_ (_08834_, _08833_, _08823_);
  or _60314_ (_08835_, _08834_, _04081_);
  and _60315_ (_08836_, _05303_, \oc8051_golden_model_1.ACC [7]);
  or _60316_ (_08837_, _08836_, _08823_);
  and _60317_ (_08838_, _08837_, _04409_);
  nor _60318_ (_08839_, _04409_, _08821_);
  or _60319_ (_08840_, _08839_, _03610_);
  or _60320_ (_08841_, _08840_, _08838_);
  and _60321_ (_08842_, _08841_, _03996_);
  and _60322_ (_08843_, _08842_, _08835_);
  and _60323_ (_08844_, _08830_, _03723_);
  or _60324_ (_08845_, _08844_, _03729_);
  or _60325_ (_08846_, _08845_, _08843_);
  nor _60326_ (_08847_, _03237_, _03215_);
  not _60327_ (_08848_, _08847_);
  or _60328_ (_08849_, _08837_, _03737_);
  and _60329_ (_08850_, _08849_, _08848_);
  and _60330_ (_08851_, _08850_, _08846_);
  and _60331_ (_08852_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and _60332_ (_08853_, _08852_, \oc8051_golden_model_1.DPL [2]);
  and _60333_ (_08854_, _08853_, \oc8051_golden_model_1.DPL [3]);
  and _60334_ (_08855_, _08854_, \oc8051_golden_model_1.DPL [4]);
  and _60335_ (_08856_, _08855_, \oc8051_golden_model_1.DPL [5]);
  and _60336_ (_08857_, _08856_, \oc8051_golden_model_1.DPL [6]);
  nor _60337_ (_08858_, _08857_, \oc8051_golden_model_1.DPL [7]);
  and _60338_ (_08859_, _08857_, \oc8051_golden_model_1.DPL [7]);
  nor _60339_ (_08860_, _08859_, _08858_);
  and _60340_ (_08861_, _08860_, _08847_);
  or _60341_ (_08862_, _08861_, _08851_);
  and _60342_ (_08863_, _08862_, _08832_);
  nor _60343_ (_08864_, _05881_, _08832_);
  or _60344_ (_08865_, _08864_, _07390_);
  or _60345_ (_08866_, _08865_, _08863_);
  and _60346_ (_08867_, _08866_, _08831_);
  or _60347_ (_08868_, _08867_, _04481_);
  and _60348_ (_08869_, _06069_, _05303_);
  or _60349_ (_08870_, _08823_, _07400_);
  or _60350_ (_08871_, _08870_, _08869_);
  and _60351_ (_08872_, _08871_, _03589_);
  and _60352_ (_08873_, _08872_, _08868_);
  nor _60353_ (_08874_, _06363_, _08824_);
  or _60354_ (_08875_, _08874_, _08823_);
  and _60355_ (_08876_, _08875_, _03222_);
  or _60356_ (_08877_, _08876_, _08873_);
  or _60357_ (_08878_, _08877_, _08828_);
  and _60358_ (_08879_, _05884_, _05303_);
  or _60359_ (_08880_, _08823_, _07766_);
  or _60360_ (_08881_, _08880_, _08879_);
  and _60361_ (_08882_, _06171_, _05303_);
  or _60362_ (_08883_, _08882_, _08823_);
  or _60363_ (_08884_, _08883_, _05886_);
  and _60364_ (_08885_, _08884_, _07778_);
  and _60365_ (_08886_, _08885_, _08881_);
  and _60366_ (_08887_, _08886_, _08878_);
  and _60367_ (_08888_, _06378_, _05303_);
  or _60368_ (_08889_, _08888_, _08823_);
  and _60369_ (_08890_, _08889_, _03780_);
  or _60370_ (_08891_, _08890_, _08887_);
  and _60371_ (_08892_, _08891_, _07777_);
  or _60372_ (_08893_, _08823_, _05310_);
  and _60373_ (_08894_, _08883_, _03622_);
  and _60374_ (_08895_, _08894_, _08893_);
  or _60375_ (_08896_, _08895_, _08892_);
  and _60376_ (_08897_, _08896_, _06828_);
  and _60377_ (_08898_, _08837_, _03790_);
  and _60378_ (_08899_, _08898_, _08893_);
  or _60379_ (_08900_, _08899_, _03624_);
  or _60380_ (_08901_, _08900_, _08897_);
  nor _60381_ (_08902_, _05882_, _08824_);
  or _60382_ (_08903_, _08823_, _07795_);
  or _60383_ (_08904_, _08903_, _08902_);
  and _60384_ (_08905_, _08904_, _07793_);
  and _60385_ (_08906_, _08905_, _08901_);
  or _60386_ (_08907_, _08906_, _08827_);
  and _60387_ (_08908_, _08907_, _04246_);
  and _60388_ (_08909_, _08834_, _03815_);
  or _60389_ (_08910_, _08909_, _03447_);
  or _60390_ (_08911_, _08910_, _08908_);
  and _60391_ (_08912_, _05831_, _05303_);
  or _60392_ (_08913_, _08823_, _03514_);
  or _60393_ (_08914_, _08913_, _08912_);
  and _60394_ (_08915_, _08914_, _43000_);
  and _60395_ (_08916_, _08915_, _08911_);
  or _60396_ (_08917_, _08916_, _08822_);
  and _60397_ (_40568_, _08917_, _41806_);
  not _60398_ (_08918_, \oc8051_golden_model_1.DPH [7]);
  nor _60399_ (_08919_, _43000_, _08918_);
  nor _60400_ (_08920_, _05297_, _08918_);
  not _60401_ (_08921_, _05297_);
  nor _60402_ (_08922_, _06377_, _08921_);
  or _60403_ (_08923_, _08922_, _08920_);
  and _60404_ (_08924_, _08923_, _03785_);
  nor _60405_ (_08925_, _08921_, _05204_);
  or _60406_ (_08926_, _08925_, _08920_);
  or _60407_ (_08927_, _08926_, _06838_);
  and _60408_ (_08928_, _05964_, _05297_);
  or _60409_ (_08929_, _08928_, _08920_);
  or _60410_ (_08930_, _08929_, _04081_);
  and _60411_ (_08931_, _05297_, \oc8051_golden_model_1.ACC [7]);
  or _60412_ (_08933_, _08931_, _08920_);
  and _60413_ (_08934_, _08933_, _04409_);
  nor _60414_ (_08935_, _04409_, _08918_);
  or _60415_ (_08936_, _08935_, _03610_);
  or _60416_ (_08937_, _08936_, _08934_);
  and _60417_ (_08938_, _08937_, _03996_);
  and _60418_ (_08939_, _08938_, _08930_);
  and _60419_ (_08940_, _08926_, _03723_);
  or _60420_ (_08941_, _08940_, _03729_);
  or _60421_ (_08942_, _08941_, _08939_);
  or _60422_ (_08944_, _08933_, _03737_);
  and _60423_ (_08945_, _08944_, _08848_);
  and _60424_ (_08946_, _08945_, _08942_);
  and _60425_ (_08947_, _08859_, \oc8051_golden_model_1.DPH [0]);
  and _60426_ (_08948_, _08947_, \oc8051_golden_model_1.DPH [1]);
  and _60427_ (_08949_, _08948_, \oc8051_golden_model_1.DPH [2]);
  and _60428_ (_08950_, _08949_, \oc8051_golden_model_1.DPH [3]);
  and _60429_ (_08951_, _08950_, \oc8051_golden_model_1.DPH [4]);
  and _60430_ (_08952_, _08951_, \oc8051_golden_model_1.DPH [5]);
  and _60431_ (_08953_, _08952_, \oc8051_golden_model_1.DPH [6]);
  nor _60432_ (_08955_, _08953_, _08918_);
  and _60433_ (_08956_, _08953_, _08918_);
  or _60434_ (_08957_, _08956_, _08955_);
  and _60435_ (_08958_, _08957_, _08847_);
  or _60436_ (_08959_, _08958_, _08946_);
  and _60437_ (_08960_, _08959_, _08832_);
  nor _60438_ (_08961_, _08832_, _03446_);
  or _60439_ (_08962_, _08961_, _07390_);
  or _60440_ (_08963_, _08962_, _08960_);
  and _60441_ (_08964_, _08963_, _08927_);
  or _60442_ (_08966_, _08964_, _04481_);
  and _60443_ (_08967_, _06069_, _05297_);
  or _60444_ (_08968_, _08920_, _07400_);
  or _60445_ (_08969_, _08968_, _08967_);
  and _60446_ (_08970_, _08969_, _03589_);
  and _60447_ (_08971_, _08970_, _08966_);
  nor _60448_ (_08972_, _06363_, _08921_);
  or _60449_ (_08973_, _08972_, _08920_);
  and _60450_ (_08974_, _08973_, _03222_);
  or _60451_ (_08975_, _08974_, _08971_);
  or _60452_ (_08977_, _08975_, _08828_);
  and _60453_ (_08978_, _05884_, _05297_);
  or _60454_ (_08979_, _08920_, _07766_);
  or _60455_ (_08980_, _08979_, _08978_);
  and _60456_ (_08981_, _06171_, _05297_);
  or _60457_ (_08982_, _08981_, _08920_);
  or _60458_ (_08983_, _08982_, _05886_);
  and _60459_ (_08984_, _08983_, _07778_);
  and _60460_ (_08985_, _08984_, _08980_);
  and _60461_ (_08986_, _08985_, _08977_);
  and _60462_ (_08988_, _06378_, _05297_);
  or _60463_ (_08989_, _08988_, _08920_);
  and _60464_ (_08990_, _08989_, _03780_);
  or _60465_ (_08991_, _08990_, _08986_);
  and _60466_ (_08992_, _08991_, _07777_);
  or _60467_ (_08993_, _08920_, _05310_);
  and _60468_ (_08994_, _08982_, _03622_);
  and _60469_ (_08995_, _08994_, _08993_);
  or _60470_ (_08996_, _08995_, _08992_);
  and _60471_ (_08997_, _08996_, _06828_);
  and _60472_ (_08999_, _08933_, _03790_);
  and _60473_ (_09000_, _08999_, _08993_);
  or _60474_ (_09001_, _09000_, _03624_);
  or _60475_ (_09002_, _09001_, _08997_);
  nor _60476_ (_09003_, _05882_, _08921_);
  or _60477_ (_09004_, _08920_, _07795_);
  or _60478_ (_09005_, _09004_, _09003_);
  and _60479_ (_09006_, _09005_, _07793_);
  and _60480_ (_09007_, _09006_, _09002_);
  or _60481_ (_09008_, _09007_, _08924_);
  and _60482_ (_09009_, _09008_, _04246_);
  and _60483_ (_09010_, _08929_, _03815_);
  or _60484_ (_09011_, _09010_, _03447_);
  or _60485_ (_09012_, _09011_, _09009_);
  and _60486_ (_09013_, _05831_, _05297_);
  or _60487_ (_09014_, _08920_, _03514_);
  or _60488_ (_09015_, _09014_, _09013_);
  and _60489_ (_09016_, _09015_, _43000_);
  and _60490_ (_09017_, _09016_, _09012_);
  or _60491_ (_09018_, _09017_, _08919_);
  and _60492_ (_40569_, _09018_, _41806_);
  not _60493_ (_09019_, \oc8051_golden_model_1.IE [7]);
  nor _60494_ (_09020_, _05229_, _09019_);
  not _60495_ (_09021_, _05229_);
  nor _60496_ (_09022_, _09021_, _05204_);
  nor _60497_ (_09023_, _09022_, _09020_);
  and _60498_ (_09024_, _09023_, _07390_);
  nor _60499_ (_09025_, _05924_, _09019_);
  and _60500_ (_09026_, _05952_, _05924_);
  nor _60501_ (_09027_, _09026_, _09025_);
  nor _60502_ (_09028_, _09027_, _03736_);
  not _60503_ (_09029_, _04409_);
  and _60504_ (_09030_, _05229_, \oc8051_golden_model_1.ACC [7]);
  nor _60505_ (_09031_, _09030_, _09020_);
  nor _60506_ (_09032_, _09031_, _09029_);
  nor _60507_ (_09033_, _04409_, _09019_);
  or _60508_ (_09034_, _09033_, _09032_);
  and _60509_ (_09035_, _09034_, _04081_);
  and _60510_ (_09036_, _05964_, _05229_);
  nor _60511_ (_09037_, _09036_, _09020_);
  nor _60512_ (_09038_, _09037_, _04081_);
  or _60513_ (_09039_, _09038_, _09035_);
  and _60514_ (_09040_, _09039_, _04055_);
  and _60515_ (_09041_, _06095_, _05924_);
  nor _60516_ (_09042_, _09041_, _09025_);
  nor _60517_ (_09043_, _09042_, _04055_);
  or _60518_ (_09044_, _09043_, _03723_);
  or _60519_ (_09045_, _09044_, _09040_);
  nand _60520_ (_09046_, _09023_, _03723_);
  and _60521_ (_09047_, _09046_, _09045_);
  and _60522_ (_09048_, _09047_, _03737_);
  nor _60523_ (_09049_, _09031_, _03737_);
  or _60524_ (_09050_, _09049_, _09048_);
  and _60525_ (_09051_, _09050_, _03736_);
  nor _60526_ (_09052_, _09051_, _09028_);
  nor _60527_ (_09053_, _09052_, _03719_);
  nor _60528_ (_09054_, _09025_, _06138_);
  or _60529_ (_09055_, _09042_, _06840_);
  nor _60530_ (_09056_, _09055_, _09054_);
  nor _60531_ (_09057_, _09056_, _09053_);
  nor _60532_ (_09058_, _09057_, _03505_);
  not _60533_ (_09059_, _05924_);
  nor _60534_ (_09060_, _05938_, _09059_);
  nor _60535_ (_09061_, _09060_, _09025_);
  nor _60536_ (_09062_, _09061_, _03710_);
  nor _60537_ (_09063_, _09062_, _07390_);
  not _60538_ (_09064_, _09063_);
  nor _60539_ (_09065_, _09064_, _09058_);
  nor _60540_ (_09066_, _09065_, _09024_);
  nor _60541_ (_09067_, _09066_, _04481_);
  and _60542_ (_09068_, _06069_, _05229_);
  nor _60543_ (_09069_, _09020_, _07400_);
  not _60544_ (_09070_, _09069_);
  nor _60545_ (_09071_, _09070_, _09068_);
  nor _60546_ (_09072_, _09071_, _03222_);
  not _60547_ (_09073_, _09072_);
  nor _60548_ (_09074_, _09073_, _09067_);
  nor _60549_ (_09075_, _06363_, _09021_);
  nor _60550_ (_09076_, _09075_, _09020_);
  nor _60551_ (_09077_, _09076_, _03589_);
  or _60552_ (_09078_, _09077_, _08828_);
  or _60553_ (_09079_, _09078_, _09074_);
  and _60554_ (_09080_, _05884_, _05229_);
  or _60555_ (_09081_, _09020_, _07766_);
  or _60556_ (_09082_, _09081_, _09080_);
  and _60557_ (_09083_, _06171_, _05229_);
  nor _60558_ (_09084_, _09083_, _09020_);
  and _60559_ (_09085_, _09084_, _03601_);
  nor _60560_ (_09086_, _09085_, _03780_);
  and _60561_ (_09087_, _09086_, _09082_);
  and _60562_ (_09088_, _09087_, _09079_);
  and _60563_ (_09089_, _06378_, _05229_);
  nor _60564_ (_09090_, _09089_, _09020_);
  nor _60565_ (_09091_, _09090_, _07778_);
  nor _60566_ (_09092_, _09091_, _09088_);
  nor _60567_ (_09093_, _09092_, _03622_);
  nor _60568_ (_09094_, _09020_, _05310_);
  not _60569_ (_09095_, _09094_);
  nor _60570_ (_09096_, _09084_, _07777_);
  and _60571_ (_09097_, _09096_, _09095_);
  nor _60572_ (_09098_, _09097_, _09093_);
  nor _60573_ (_09099_, _09098_, _03790_);
  nor _60574_ (_09100_, _09031_, _06828_);
  and _60575_ (_09101_, _09100_, _09095_);
  or _60576_ (_09102_, _09101_, _09099_);
  and _60577_ (_09103_, _09102_, _07795_);
  nor _60578_ (_09104_, _05882_, _09021_);
  nor _60579_ (_09105_, _09104_, _09020_);
  nor _60580_ (_09106_, _09105_, _07795_);
  or _60581_ (_09107_, _09106_, _09103_);
  and _60582_ (_09108_, _09107_, _07793_);
  nor _60583_ (_09109_, _06377_, _09021_);
  nor _60584_ (_09110_, _09109_, _09020_);
  nor _60585_ (_09111_, _09110_, _07793_);
  or _60586_ (_09112_, _09111_, _09108_);
  and _60587_ (_09113_, _09112_, _04246_);
  nor _60588_ (_09114_, _09037_, _04246_);
  or _60589_ (_09115_, _09114_, _09113_);
  and _60590_ (_09116_, _09115_, _03823_);
  nor _60591_ (_09117_, _09027_, _03823_);
  or _60592_ (_09118_, _09117_, _09116_);
  and _60593_ (_09119_, _09118_, _03514_);
  and _60594_ (_09120_, _05831_, _05229_);
  nor _60595_ (_09121_, _09120_, _09020_);
  nor _60596_ (_09122_, _09121_, _03514_);
  or _60597_ (_09123_, _09122_, _09119_);
  or _60598_ (_09124_, _09123_, _43004_);
  or _60599_ (_09125_, _43000_, \oc8051_golden_model_1.IE [7]);
  and _60600_ (_09126_, _09125_, _41806_);
  and _60601_ (_40571_, _09126_, _09124_);
  not _60602_ (_09127_, \oc8051_golden_model_1.IP [7]);
  nor _60603_ (_09128_, _05251_, _09127_);
  not _60604_ (_09129_, _05251_);
  nor _60605_ (_09130_, _09129_, _05204_);
  nor _60606_ (_09131_, _09130_, _09128_);
  and _60607_ (_09132_, _09131_, _07390_);
  nor _60608_ (_09133_, _05908_, _09127_);
  and _60609_ (_09134_, _05952_, _05908_);
  nor _60610_ (_09135_, _09134_, _09133_);
  nor _60611_ (_09136_, _09135_, _03736_);
  and _60612_ (_09137_, _05251_, \oc8051_golden_model_1.ACC [7]);
  nor _60613_ (_09138_, _09137_, _09128_);
  nor _60614_ (_09139_, _09138_, _09029_);
  nor _60615_ (_09140_, _04409_, _09127_);
  or _60616_ (_09141_, _09140_, _09139_);
  and _60617_ (_09142_, _09141_, _04081_);
  and _60618_ (_09143_, _05964_, _05251_);
  nor _60619_ (_09144_, _09143_, _09128_);
  nor _60620_ (_09145_, _09144_, _04081_);
  or _60621_ (_09146_, _09145_, _09142_);
  and _60622_ (_09147_, _09146_, _04055_);
  and _60623_ (_09148_, _06095_, _05908_);
  nor _60624_ (_09149_, _09148_, _09133_);
  nor _60625_ (_09150_, _09149_, _04055_);
  or _60626_ (_09151_, _09150_, _03723_);
  or _60627_ (_09152_, _09151_, _09147_);
  nand _60628_ (_09153_, _09131_, _03723_);
  and _60629_ (_09154_, _09153_, _09152_);
  and _60630_ (_09155_, _09154_, _03737_);
  nor _60631_ (_09156_, _09138_, _03737_);
  or _60632_ (_09157_, _09156_, _09155_);
  and _60633_ (_09158_, _09157_, _03736_);
  nor _60634_ (_09159_, _09158_, _09136_);
  nor _60635_ (_09160_, _09159_, _03719_);
  nor _60636_ (_09161_, _09133_, _06138_);
  or _60637_ (_09162_, _09149_, _06840_);
  nor _60638_ (_09163_, _09162_, _09161_);
  nor _60639_ (_09164_, _09163_, _09160_);
  nor _60640_ (_09165_, _09164_, _03505_);
  not _60641_ (_09166_, _05908_);
  nor _60642_ (_09167_, _05938_, _09166_);
  nor _60643_ (_09168_, _09167_, _09133_);
  nor _60644_ (_09169_, _09168_, _03710_);
  nor _60645_ (_09170_, _09169_, _07390_);
  not _60646_ (_09171_, _09170_);
  nor _60647_ (_09172_, _09171_, _09165_);
  nor _60648_ (_09173_, _09172_, _09132_);
  nor _60649_ (_09174_, _09173_, _04481_);
  and _60650_ (_09175_, _06069_, _05251_);
  nor _60651_ (_09176_, _09128_, _07400_);
  not _60652_ (_09177_, _09176_);
  nor _60653_ (_09178_, _09177_, _09175_);
  nor _60654_ (_09179_, _09178_, _03222_);
  not _60655_ (_09180_, _09179_);
  nor _60656_ (_09181_, _09180_, _09174_);
  nor _60657_ (_09182_, _06363_, _09129_);
  nor _60658_ (_09183_, _09182_, _09128_);
  nor _60659_ (_09184_, _09183_, _03589_);
  or _60660_ (_09185_, _09184_, _08828_);
  or _60661_ (_09186_, _09185_, _09181_);
  and _60662_ (_09187_, _05884_, _05251_);
  or _60663_ (_09188_, _09128_, _07766_);
  or _60664_ (_09189_, _09188_, _09187_);
  and _60665_ (_09190_, _06171_, _05251_);
  nor _60666_ (_09191_, _09190_, _09128_);
  and _60667_ (_09192_, _09191_, _03601_);
  nor _60668_ (_09193_, _09192_, _03780_);
  and _60669_ (_09194_, _09193_, _09189_);
  and _60670_ (_09195_, _09194_, _09186_);
  and _60671_ (_09196_, _06378_, _05251_);
  nor _60672_ (_09197_, _09196_, _09128_);
  nor _60673_ (_09198_, _09197_, _07778_);
  nor _60674_ (_09199_, _09198_, _09195_);
  nor _60675_ (_09200_, _09199_, _03622_);
  nor _60676_ (_09201_, _09128_, _05310_);
  not _60677_ (_09202_, _09201_);
  nor _60678_ (_09203_, _09191_, _07777_);
  and _60679_ (_09204_, _09203_, _09202_);
  nor _60680_ (_09205_, _09204_, _09200_);
  nor _60681_ (_09206_, _09205_, _03790_);
  nor _60682_ (_09207_, _09138_, _06828_);
  and _60683_ (_09208_, _09207_, _09202_);
  or _60684_ (_09209_, _09208_, _09206_);
  and _60685_ (_09210_, _09209_, _07795_);
  nor _60686_ (_09211_, _05882_, _09129_);
  nor _60687_ (_09212_, _09211_, _09128_);
  nor _60688_ (_09213_, _09212_, _07795_);
  or _60689_ (_09214_, _09213_, _09210_);
  and _60690_ (_09215_, _09214_, _07793_);
  nor _60691_ (_09216_, _06377_, _09129_);
  nor _60692_ (_09217_, _09216_, _09128_);
  nor _60693_ (_09218_, _09217_, _07793_);
  or _60694_ (_09219_, _09218_, _09215_);
  and _60695_ (_09220_, _09219_, _04246_);
  nor _60696_ (_09221_, _09144_, _04246_);
  or _60697_ (_09222_, _09221_, _09220_);
  and _60698_ (_09223_, _09222_, _03823_);
  nor _60699_ (_09224_, _09135_, _03823_);
  or _60700_ (_09225_, _09224_, _09223_);
  and _60701_ (_09226_, _09225_, _03514_);
  and _60702_ (_09227_, _05831_, _05251_);
  nor _60703_ (_09228_, _09227_, _09128_);
  nor _60704_ (_09229_, _09228_, _03514_);
  or _60705_ (_09230_, _09229_, _09226_);
  or _60706_ (_09231_, _09230_, _43004_);
  or _60707_ (_09232_, _43000_, \oc8051_golden_model_1.IP [7]);
  and _60708_ (_09233_, _09232_, _41806_);
  and _60709_ (_40572_, _09233_, _09231_);
  not _60710_ (_09234_, \oc8051_golden_model_1.P0 [7]);
  nor _60711_ (_09235_, _05293_, _09234_);
  not _60712_ (_09236_, _05293_);
  nor _60713_ (_09237_, _09236_, _05204_);
  or _60714_ (_09238_, _09237_, _09235_);
  or _60715_ (_09239_, _09238_, _06838_);
  nor _60716_ (_09240_, _05209_, _09234_);
  and _60717_ (_09241_, _05952_, _05209_);
  or _60718_ (_09242_, _09241_, _09240_);
  and _60719_ (_09243_, _09242_, _03714_);
  and _60720_ (_09244_, _05964_, _05293_);
  or _60721_ (_09245_, _09244_, _09235_);
  or _60722_ (_09246_, _09245_, _04081_);
  and _60723_ (_09247_, _05293_, \oc8051_golden_model_1.ACC [7]);
  or _60724_ (_09248_, _09247_, _09235_);
  and _60725_ (_09249_, _09248_, _04409_);
  nor _60726_ (_09250_, _04409_, _09234_);
  or _60727_ (_09251_, _09250_, _03610_);
  or _60728_ (_09252_, _09251_, _09249_);
  and _60729_ (_09253_, _09252_, _04055_);
  and _60730_ (_09254_, _09253_, _09246_);
  and _60731_ (_09255_, _06095_, _05209_);
  or _60732_ (_09256_, _09255_, _09240_);
  and _60733_ (_09257_, _09256_, _03715_);
  or _60734_ (_09258_, _09257_, _03723_);
  or _60735_ (_09259_, _09258_, _09254_);
  or _60736_ (_09260_, _09238_, _03996_);
  and _60737_ (_09261_, _09260_, _09259_);
  or _60738_ (_09262_, _09261_, _03729_);
  or _60739_ (_09263_, _09248_, _03737_);
  and _60740_ (_09264_, _09263_, _03736_);
  and _60741_ (_09265_, _09264_, _09262_);
  or _60742_ (_09266_, _09265_, _09243_);
  and _60743_ (_09267_, _09266_, _06840_);
  or _60744_ (_09268_, _09240_, _06138_);
  and _60745_ (_09269_, _09268_, _03719_);
  and _60746_ (_09270_, _09269_, _09256_);
  or _60747_ (_09271_, _09270_, _09267_);
  and _60748_ (_09272_, _09271_, _03710_);
  or _60749_ (_09273_, _05952_, _05937_);
  and _60750_ (_09274_, _09273_, _05209_);
  or _60751_ (_09275_, _09274_, _09240_);
  and _60752_ (_09276_, _09275_, _03505_);
  or _60753_ (_09277_, _09276_, _07390_);
  or _60754_ (_09278_, _09277_, _09272_);
  and _60755_ (_09279_, _09278_, _09239_);
  or _60756_ (_09280_, _09279_, _04481_);
  and _60757_ (_09281_, _06069_, _05293_);
  or _60758_ (_09282_, _09235_, _07400_);
  or _60759_ (_09283_, _09282_, _09281_);
  and _60760_ (_09284_, _09283_, _03589_);
  and _60761_ (_09285_, _09284_, _09280_);
  and _60762_ (_09286_, _06340_, \oc8051_golden_model_1.P1 [7]);
  and _60763_ (_09287_, _06343_, \oc8051_golden_model_1.P0 [7]);
  and _60764_ (_09288_, _06346_, \oc8051_golden_model_1.P2 [7]);
  and _60765_ (_09289_, _06348_, \oc8051_golden_model_1.P3 [7]);
  or _60766_ (_09290_, _09289_, _09288_);
  or _60767_ (_09291_, _09290_, _09287_);
  nor _60768_ (_09292_, _09291_, _09286_);
  and _60769_ (_09293_, _09292_, _06358_);
  and _60770_ (_09294_, _09293_, _06339_);
  nand _60771_ (_09295_, _09294_, _06326_);
  or _60772_ (_09296_, _09295_, _06172_);
  and _60773_ (_09297_, _09296_, _05293_);
  or _60774_ (_09298_, _09297_, _09235_);
  and _60775_ (_09299_, _09298_, _03222_);
  or _60776_ (_09300_, _09299_, _08828_);
  or _60777_ (_09301_, _09300_, _09285_);
  and _60778_ (_09302_, _05884_, _05293_);
  or _60779_ (_09303_, _09235_, _07766_);
  or _60780_ (_09304_, _09303_, _09302_);
  and _60781_ (_09305_, _06171_, _05293_);
  or _60782_ (_09306_, _09305_, _09235_);
  or _60783_ (_09307_, _09306_, _05886_);
  and _60784_ (_09308_, _09307_, _07778_);
  and _60785_ (_09309_, _09308_, _09304_);
  and _60786_ (_09310_, _09309_, _09301_);
  and _60787_ (_09311_, _06378_, _05293_);
  or _60788_ (_09312_, _09311_, _09235_);
  and _60789_ (_09313_, _09312_, _03780_);
  or _60790_ (_09314_, _09313_, _09310_);
  and _60791_ (_09315_, _09314_, _07777_);
  or _60792_ (_09316_, _09235_, _05310_);
  and _60793_ (_09317_, _09306_, _03622_);
  and _60794_ (_09318_, _09317_, _09316_);
  or _60795_ (_09319_, _09318_, _09315_);
  and _60796_ (_09320_, _09319_, _06828_);
  and _60797_ (_09321_, _09248_, _03790_);
  and _60798_ (_09322_, _09321_, _09316_);
  or _60799_ (_09323_, _09322_, _03624_);
  or _60800_ (_09324_, _09323_, _09320_);
  nor _60801_ (_09325_, _05882_, _09236_);
  or _60802_ (_09326_, _09235_, _07795_);
  or _60803_ (_09327_, _09326_, _09325_);
  and _60804_ (_09328_, _09327_, _07793_);
  and _60805_ (_09329_, _09328_, _09324_);
  nor _60806_ (_09330_, _06377_, _09236_);
  or _60807_ (_09331_, _09330_, _09235_);
  and _60808_ (_09332_, _09331_, _03785_);
  or _60809_ (_09333_, _09332_, _03815_);
  or _60810_ (_09334_, _09333_, _09329_);
  or _60811_ (_09335_, _09245_, _04246_);
  and _60812_ (_09336_, _09335_, _03823_);
  and _60813_ (_09337_, _09336_, _09334_);
  and _60814_ (_09338_, _09242_, _03453_);
  or _60815_ (_09339_, _09338_, _03447_);
  or _60816_ (_09340_, _09339_, _09337_);
  and _60817_ (_09341_, _05831_, _05293_);
  or _60818_ (_09342_, _09235_, _03514_);
  or _60819_ (_09343_, _09342_, _09341_);
  and _60820_ (_09344_, _09343_, _43000_);
  and _60821_ (_09345_, _09344_, _09340_);
  nor _60822_ (_09346_, _43000_, _09234_);
  or _60823_ (_09347_, _09346_, rst);
  or _60824_ (_40573_, _09347_, _09345_);
  not _60825_ (_09348_, \oc8051_golden_model_1.P1 [7]);
  nor _60826_ (_09349_, _43000_, _09348_);
  or _60827_ (_09350_, _09349_, rst);
  nor _60828_ (_09351_, _05266_, _09348_);
  not _60829_ (_09352_, _05266_);
  nor _60830_ (_09353_, _09352_, _05204_);
  or _60831_ (_09354_, _09353_, _09351_);
  or _60832_ (_09355_, _09354_, _06838_);
  nor _60833_ (_09356_, _05916_, _09348_);
  and _60834_ (_09357_, _05952_, _05916_);
  or _60835_ (_09358_, _09357_, _09356_);
  and _60836_ (_09359_, _09358_, _03714_);
  and _60837_ (_09360_, _05964_, _05266_);
  or _60838_ (_09361_, _09360_, _09351_);
  or _60839_ (_09362_, _09361_, _04081_);
  and _60840_ (_09363_, _05266_, \oc8051_golden_model_1.ACC [7]);
  or _60841_ (_09364_, _09363_, _09351_);
  and _60842_ (_09365_, _09364_, _04409_);
  nor _60843_ (_09366_, _04409_, _09348_);
  or _60844_ (_09367_, _09366_, _03610_);
  or _60845_ (_09368_, _09367_, _09365_);
  and _60846_ (_09369_, _09368_, _04055_);
  and _60847_ (_09370_, _09369_, _09362_);
  and _60848_ (_09371_, _06095_, _05916_);
  or _60849_ (_09372_, _09371_, _09356_);
  and _60850_ (_09373_, _09372_, _03715_);
  or _60851_ (_09374_, _09373_, _03723_);
  or _60852_ (_09375_, _09374_, _09370_);
  or _60853_ (_09376_, _09354_, _03996_);
  and _60854_ (_09377_, _09376_, _09375_);
  or _60855_ (_09378_, _09377_, _03729_);
  or _60856_ (_09379_, _09364_, _03737_);
  and _60857_ (_09380_, _09379_, _03736_);
  and _60858_ (_09381_, _09380_, _09378_);
  or _60859_ (_09382_, _09381_, _09359_);
  and _60860_ (_09383_, _09382_, _06840_);
  and _60861_ (_09384_, _06139_, _05916_);
  or _60862_ (_09385_, _09384_, _09356_);
  and _60863_ (_09386_, _09385_, _03719_);
  or _60864_ (_09387_, _09386_, _09383_);
  and _60865_ (_09388_, _09387_, _03710_);
  and _60866_ (_09389_, _09273_, _05916_);
  or _60867_ (_09390_, _09389_, _09356_);
  and _60868_ (_09391_, _09390_, _03505_);
  or _60869_ (_09392_, _09391_, _07390_);
  or _60870_ (_09393_, _09392_, _09388_);
  and _60871_ (_09394_, _09393_, _09355_);
  or _60872_ (_09395_, _09394_, _04481_);
  and _60873_ (_09396_, _06069_, _05266_);
  or _60874_ (_09397_, _09351_, _07400_);
  or _60875_ (_09398_, _09397_, _09396_);
  and _60876_ (_09399_, _09398_, _03589_);
  and _60877_ (_09400_, _09399_, _09395_);
  and _60878_ (_09401_, _09296_, _05266_);
  or _60879_ (_09402_, _09401_, _09351_);
  and _60880_ (_09403_, _09402_, _03222_);
  or _60881_ (_09404_, _09403_, _08828_);
  or _60882_ (_09405_, _09404_, _09400_);
  and _60883_ (_09406_, _05884_, _05266_);
  or _60884_ (_09407_, _09351_, _07766_);
  or _60885_ (_09408_, _09407_, _09406_);
  and _60886_ (_09409_, _06171_, _05266_);
  or _60887_ (_09410_, _09409_, _09351_);
  or _60888_ (_09411_, _09410_, _05886_);
  and _60889_ (_09412_, _09411_, _07778_);
  and _60890_ (_09413_, _09412_, _09408_);
  and _60891_ (_09414_, _09413_, _09405_);
  and _60892_ (_09415_, _06378_, _05266_);
  or _60893_ (_09416_, _09415_, _09351_);
  and _60894_ (_09417_, _09416_, _03780_);
  or _60895_ (_09418_, _09417_, _09414_);
  and _60896_ (_09419_, _09418_, _07777_);
  or _60897_ (_09420_, _09351_, _05310_);
  and _60898_ (_09421_, _09410_, _03622_);
  and _60899_ (_09422_, _09421_, _09420_);
  or _60900_ (_09423_, _09422_, _09419_);
  and _60901_ (_09424_, _09423_, _06828_);
  and _60902_ (_09425_, _09364_, _03790_);
  and _60903_ (_09426_, _09425_, _09420_);
  or _60904_ (_09427_, _09426_, _03624_);
  or _60905_ (_09428_, _09427_, _09424_);
  nor _60906_ (_09429_, _05882_, _09352_);
  or _60907_ (_09430_, _09351_, _07795_);
  or _60908_ (_09431_, _09430_, _09429_);
  and _60909_ (_09432_, _09431_, _07793_);
  and _60910_ (_09433_, _09432_, _09428_);
  nor _60911_ (_09434_, _06377_, _09352_);
  or _60912_ (_09435_, _09434_, _09351_);
  and _60913_ (_09436_, _09435_, _03785_);
  or _60914_ (_09437_, _09436_, _03815_);
  or _60915_ (_09438_, _09437_, _09433_);
  or _60916_ (_09439_, _09361_, _04246_);
  and _60917_ (_09440_, _09439_, _03823_);
  and _60918_ (_09441_, _09440_, _09438_);
  and _60919_ (_09442_, _09358_, _03453_);
  or _60920_ (_09443_, _09442_, _03447_);
  or _60921_ (_09444_, _09443_, _09441_);
  and _60922_ (_09445_, _05831_, _05266_);
  or _60923_ (_09446_, _09351_, _03514_);
  or _60924_ (_09447_, _09446_, _09445_);
  and _60925_ (_09448_, _09447_, _43000_);
  and _60926_ (_09449_, _09448_, _09444_);
  or _60927_ (_40574_, _09449_, _09350_);
  not _60928_ (_09450_, \oc8051_golden_model_1.P2 [7]);
  nor _60929_ (_09451_, _43000_, _09450_);
  or _60930_ (_09452_, _09451_, rst);
  nor _60931_ (_09453_, _05235_, _09450_);
  not _60932_ (_09454_, _05235_);
  nor _60933_ (_09455_, _09454_, _05204_);
  or _60934_ (_09456_, _09455_, _09453_);
  or _60935_ (_09457_, _09456_, _06838_);
  nor _60936_ (_09458_, _05918_, _09450_);
  and _60937_ (_09459_, _05952_, _05918_);
  or _60938_ (_09460_, _09459_, _09458_);
  and _60939_ (_09461_, _09460_, _03714_);
  and _60940_ (_09462_, _05964_, _05235_);
  or _60941_ (_09463_, _09462_, _09453_);
  or _60942_ (_09464_, _09463_, _04081_);
  and _60943_ (_09465_, _05235_, \oc8051_golden_model_1.ACC [7]);
  or _60944_ (_09466_, _09465_, _09453_);
  and _60945_ (_09467_, _09466_, _04409_);
  nor _60946_ (_09468_, _04409_, _09450_);
  or _60947_ (_09469_, _09468_, _03610_);
  or _60948_ (_09470_, _09469_, _09467_);
  and _60949_ (_09471_, _09470_, _04055_);
  and _60950_ (_09472_, _09471_, _09464_);
  and _60951_ (_09473_, _06095_, _05918_);
  or _60952_ (_09474_, _09473_, _09458_);
  and _60953_ (_09475_, _09474_, _03715_);
  or _60954_ (_09476_, _09475_, _03723_);
  or _60955_ (_09477_, _09476_, _09472_);
  or _60956_ (_09478_, _09456_, _03996_);
  and _60957_ (_09479_, _09478_, _09477_);
  or _60958_ (_09480_, _09479_, _03729_);
  or _60959_ (_09481_, _09466_, _03737_);
  and _60960_ (_09482_, _09481_, _03736_);
  and _60961_ (_09483_, _09482_, _09480_);
  or _60962_ (_09484_, _09483_, _09461_);
  and _60963_ (_09485_, _09484_, _06840_);
  and _60964_ (_09486_, _06139_, _05918_);
  or _60965_ (_09487_, _09486_, _09458_);
  and _60966_ (_09488_, _09487_, _03719_);
  or _60967_ (_09489_, _09488_, _09485_);
  and _60968_ (_09490_, _09489_, _03710_);
  and _60969_ (_09491_, _09273_, _05918_);
  or _60970_ (_09492_, _09491_, _09458_);
  and _60971_ (_09493_, _09492_, _03505_);
  or _60972_ (_09494_, _09493_, _07390_);
  or _60973_ (_09495_, _09494_, _09490_);
  and _60974_ (_09496_, _09495_, _09457_);
  or _60975_ (_09497_, _09496_, _04481_);
  and _60976_ (_09498_, _06069_, _05235_);
  or _60977_ (_09499_, _09453_, _07400_);
  or _60978_ (_09500_, _09499_, _09498_);
  and _60979_ (_09501_, _09500_, _03589_);
  and _60980_ (_09502_, _09501_, _09497_);
  and _60981_ (_09503_, _09296_, _05235_);
  or _60982_ (_09504_, _09503_, _09453_);
  and _60983_ (_09505_, _09504_, _03222_);
  or _60984_ (_09506_, _09505_, _08828_);
  or _60985_ (_09507_, _09506_, _09502_);
  and _60986_ (_09508_, _05884_, _05235_);
  or _60987_ (_09509_, _09453_, _07766_);
  or _60988_ (_09510_, _09509_, _09508_);
  and _60989_ (_09511_, _06171_, _05235_);
  or _60990_ (_09512_, _09511_, _09453_);
  or _60991_ (_09513_, _09512_, _05886_);
  and _60992_ (_09514_, _09513_, _07778_);
  and _60993_ (_09515_, _09514_, _09510_);
  and _60994_ (_09516_, _09515_, _09507_);
  and _60995_ (_09517_, _06378_, _05235_);
  or _60996_ (_09518_, _09517_, _09453_);
  and _60997_ (_09519_, _09518_, _03780_);
  or _60998_ (_09520_, _09519_, _09516_);
  and _60999_ (_09521_, _09520_, _07777_);
  or _61000_ (_09522_, _09453_, _05310_);
  and _61001_ (_09523_, _09512_, _03622_);
  and _61002_ (_09524_, _09523_, _09522_);
  or _61003_ (_09525_, _09524_, _09521_);
  and _61004_ (_09526_, _09525_, _06828_);
  and _61005_ (_09527_, _09466_, _03790_);
  and _61006_ (_09528_, _09527_, _09522_);
  or _61007_ (_09529_, _09528_, _03624_);
  or _61008_ (_09530_, _09529_, _09526_);
  nor _61009_ (_09531_, _05882_, _09454_);
  or _61010_ (_09532_, _09453_, _07795_);
  or _61011_ (_09533_, _09532_, _09531_);
  and _61012_ (_09534_, _09533_, _07793_);
  and _61013_ (_09535_, _09534_, _09530_);
  nor _61014_ (_09536_, _06377_, _09454_);
  or _61015_ (_09537_, _09536_, _09453_);
  and _61016_ (_09538_, _09537_, _03785_);
  or _61017_ (_09539_, _09538_, _03815_);
  or _61018_ (_09540_, _09539_, _09535_);
  or _61019_ (_09541_, _09463_, _04246_);
  and _61020_ (_09542_, _09541_, _03823_);
  and _61021_ (_09543_, _09542_, _09540_);
  and _61022_ (_09545_, _09460_, _03453_);
  or _61023_ (_09546_, _09545_, _03447_);
  or _61024_ (_09547_, _09546_, _09543_);
  and _61025_ (_09548_, _05831_, _05235_);
  or _61026_ (_09549_, _09453_, _03514_);
  or _61027_ (_09550_, _09549_, _09548_);
  and _61028_ (_09551_, _09550_, _43000_);
  and _61029_ (_09552_, _09551_, _09547_);
  or _61030_ (_40575_, _09552_, _09452_);
  not _61031_ (_09553_, \oc8051_golden_model_1.P3 [7]);
  nor _61032_ (_09554_, _43000_, _09553_);
  or _61033_ (_09555_, _09554_, rst);
  nor _61034_ (_09556_, _05239_, _09553_);
  not _61035_ (_09557_, _05239_);
  nor _61036_ (_09558_, _09557_, _05204_);
  or _61037_ (_09559_, _09558_, _09556_);
  or _61038_ (_09560_, _09559_, _06838_);
  nor _61039_ (_09561_, _05929_, _09553_);
  and _61040_ (_09562_, _05952_, _05929_);
  or _61041_ (_09563_, _09562_, _09561_);
  and _61042_ (_09565_, _09563_, _03714_);
  and _61043_ (_09566_, _05964_, _05239_);
  or _61044_ (_09567_, _09566_, _09556_);
  or _61045_ (_09568_, _09567_, _04081_);
  and _61046_ (_09569_, _05239_, \oc8051_golden_model_1.ACC [7]);
  or _61047_ (_09570_, _09569_, _09556_);
  and _61048_ (_09571_, _09570_, _04409_);
  nor _61049_ (_09572_, _04409_, _09553_);
  or _61050_ (_09573_, _09572_, _03610_);
  or _61051_ (_09574_, _09573_, _09571_);
  and _61052_ (_09575_, _09574_, _04055_);
  and _61053_ (_09576_, _09575_, _09568_);
  and _61054_ (_09577_, _06095_, _05929_);
  or _61055_ (_09578_, _09577_, _09561_);
  and _61056_ (_09579_, _09578_, _03715_);
  or _61057_ (_09580_, _09579_, _03723_);
  or _61058_ (_09581_, _09580_, _09576_);
  or _61059_ (_09582_, _09559_, _03996_);
  and _61060_ (_09583_, _09582_, _09581_);
  or _61061_ (_09584_, _09583_, _03729_);
  or _61062_ (_09585_, _09570_, _03737_);
  and _61063_ (_09586_, _09585_, _03736_);
  and _61064_ (_09587_, _09586_, _09584_);
  or _61065_ (_09588_, _09587_, _09565_);
  and _61066_ (_09589_, _09588_, _06840_);
  and _61067_ (_09590_, _06139_, _05929_);
  or _61068_ (_09591_, _09590_, _09561_);
  and _61069_ (_09592_, _09591_, _03719_);
  or _61070_ (_09593_, _09592_, _09589_);
  and _61071_ (_09594_, _09593_, _03710_);
  and _61072_ (_09595_, _09273_, _05929_);
  or _61073_ (_09596_, _09595_, _09561_);
  and _61074_ (_09597_, _09596_, _03505_);
  or _61075_ (_09598_, _09597_, _07390_);
  or _61076_ (_09599_, _09598_, _09594_);
  and _61077_ (_09600_, _09599_, _09560_);
  or _61078_ (_09601_, _09600_, _04481_);
  and _61079_ (_09602_, _06069_, _05239_);
  or _61080_ (_09603_, _09556_, _07400_);
  or _61081_ (_09604_, _09603_, _09602_);
  and _61082_ (_09605_, _09604_, _03589_);
  and _61083_ (_09606_, _09605_, _09601_);
  and _61084_ (_09607_, _09296_, _05239_);
  or _61085_ (_09608_, _09607_, _09556_);
  and _61086_ (_09609_, _09608_, _03222_);
  or _61087_ (_09610_, _09609_, _08828_);
  or _61088_ (_09611_, _09610_, _09606_);
  and _61089_ (_09612_, _05884_, _05239_);
  or _61090_ (_09613_, _09556_, _07766_);
  or _61091_ (_09614_, _09613_, _09612_);
  and _61092_ (_09615_, _06171_, _05239_);
  or _61093_ (_09616_, _09615_, _09556_);
  or _61094_ (_09617_, _09616_, _05886_);
  and _61095_ (_09618_, _09617_, _07778_);
  and _61096_ (_09619_, _09618_, _09614_);
  and _61097_ (_09620_, _09619_, _09611_);
  and _61098_ (_09621_, _06378_, _05239_);
  or _61099_ (_09622_, _09621_, _09556_);
  and _61100_ (_09623_, _09622_, _03780_);
  or _61101_ (_09624_, _09623_, _09620_);
  and _61102_ (_09625_, _09624_, _07777_);
  or _61103_ (_09626_, _09556_, _05310_);
  and _61104_ (_09627_, _09616_, _03622_);
  and _61105_ (_09628_, _09627_, _09626_);
  or _61106_ (_09629_, _09628_, _09625_);
  and _61107_ (_09630_, _09629_, _06828_);
  and _61108_ (_09631_, _09570_, _03790_);
  and _61109_ (_09632_, _09631_, _09626_);
  or _61110_ (_09633_, _09632_, _03624_);
  or _61111_ (_09634_, _09633_, _09630_);
  nor _61112_ (_09635_, _05882_, _09557_);
  or _61113_ (_09636_, _09556_, _07795_);
  or _61114_ (_09637_, _09636_, _09635_);
  and _61115_ (_09638_, _09637_, _07793_);
  and _61116_ (_09639_, _09638_, _09634_);
  nor _61117_ (_09640_, _06377_, _09557_);
  or _61118_ (_09641_, _09640_, _09556_);
  and _61119_ (_09642_, _09641_, _03785_);
  or _61120_ (_09643_, _09642_, _03815_);
  or _61121_ (_09644_, _09643_, _09639_);
  or _61122_ (_09645_, _09567_, _04246_);
  and _61123_ (_09646_, _09645_, _03823_);
  and _61124_ (_09647_, _09646_, _09644_);
  and _61125_ (_09648_, _09563_, _03453_);
  or _61126_ (_09649_, _09648_, _03447_);
  or _61127_ (_09650_, _09649_, _09647_);
  and _61128_ (_09651_, _05831_, _05239_);
  or _61129_ (_09652_, _09556_, _03514_);
  or _61130_ (_09653_, _09652_, _09651_);
  and _61131_ (_09654_, _09653_, _43000_);
  and _61132_ (_09655_, _09654_, _09650_);
  or _61133_ (_40577_, _09655_, _09555_);
  and _61134_ (_09656_, _08780_, \oc8051_golden_model_1.ACC [0]);
  nor _61135_ (_09657_, _05245_, _07871_);
  and _61136_ (_09658_, _06378_, _05245_);
  or _61137_ (_09659_, _09658_, _09657_);
  and _61138_ (_09660_, _09659_, _03780_);
  not _61139_ (_09661_, _05245_);
  nor _61140_ (_09662_, _06363_, _09661_);
  or _61141_ (_09663_, _09662_, _09657_);
  and _61142_ (_09664_, _09663_, _03222_);
  nor _61143_ (_09665_, _09661_, _05204_);
  or _61144_ (_09666_, _09665_, _09657_);
  or _61145_ (_09667_, _09666_, _06838_);
  not _61146_ (_09668_, _03752_);
  not _61147_ (_09669_, _03753_);
  not _61148_ (_09670_, _05302_);
  and _61149_ (_09671_, _05927_, \oc8051_golden_model_1.TCON [2]);
  and _61150_ (_09672_, _05910_, \oc8051_golden_model_1.B [2]);
  nor _61151_ (_09673_, _09672_, _09671_);
  and _61152_ (_09674_, _05908_, \oc8051_golden_model_1.IP [2]);
  not _61153_ (_09675_, _09674_);
  and _61154_ (_09676_, _05901_, \oc8051_golden_model_1.PSW [2]);
  and _61155_ (_09677_, _05903_, \oc8051_golden_model_1.ACC [2]);
  nor _61156_ (_09678_, _09677_, _09676_);
  and _61157_ (_09679_, _09678_, _09675_);
  and _61158_ (_09680_, _09679_, _09673_);
  and _61159_ (_09681_, _05922_, \oc8051_golden_model_1.SCON [2]);
  and _61160_ (_09682_, _05924_, \oc8051_golden_model_1.IE [2]);
  nor _61161_ (_09683_, _09682_, _09681_);
  and _61162_ (_09684_, _05209_, \oc8051_golden_model_1.P0INREG [2]);
  and _61163_ (_09685_, _05918_, \oc8051_golden_model_1.P2INREG [2]);
  nor _61164_ (_09686_, _09685_, _09684_);
  and _61165_ (_09687_, _05916_, \oc8051_golden_model_1.P1INREG [2]);
  and _61166_ (_09688_, _05929_, \oc8051_golden_model_1.P3INREG [2]);
  nor _61167_ (_09689_, _09688_, _09687_);
  and _61168_ (_09690_, _09689_, _09686_);
  and _61169_ (_09691_, _09690_, _09683_);
  and _61170_ (_09692_, _09691_, _09680_);
  and _61171_ (_09693_, _09692_, _05668_);
  nor _61172_ (_09694_, _09693_, _09670_);
  not _61173_ (_09695_, _05216_);
  and _61174_ (_09696_, _05901_, \oc8051_golden_model_1.PSW [1]);
  and _61175_ (_09697_, _05910_, \oc8051_golden_model_1.B [1]);
  nor _61176_ (_09698_, _09697_, _09696_);
  and _61177_ (_09699_, _05908_, \oc8051_golden_model_1.IP [1]);
  and _61178_ (_09700_, _05903_, \oc8051_golden_model_1.ACC [1]);
  nor _61179_ (_09701_, _09700_, _09699_);
  and _61180_ (_09702_, _09701_, _09698_);
  and _61181_ (_09703_, _05929_, \oc8051_golden_model_1.P3INREG [1]);
  not _61182_ (_09704_, _09703_);
  and _61183_ (_09705_, _05209_, \oc8051_golden_model_1.P0INREG [1]);
  and _61184_ (_09706_, _05918_, \oc8051_golden_model_1.P2INREG [1]);
  nor _61185_ (_09707_, _09706_, _09705_);
  and _61186_ (_09708_, _09707_, _09704_);
  and _61187_ (_09709_, _05922_, \oc8051_golden_model_1.SCON [1]);
  and _61188_ (_09710_, _05924_, \oc8051_golden_model_1.IE [1]);
  nor _61189_ (_09711_, _09710_, _09709_);
  and _61190_ (_09712_, _05927_, \oc8051_golden_model_1.TCON [1]);
  and _61191_ (_09713_, _05916_, \oc8051_golden_model_1.P1INREG [1]);
  nor _61192_ (_09714_, _09713_, _09712_);
  and _61193_ (_09715_, _09714_, _09711_);
  and _61194_ (_09716_, _09715_, _09708_);
  and _61195_ (_09717_, _09716_, _09702_);
  and _61196_ (_09718_, _09717_, _05568_);
  nor _61197_ (_09719_, _09718_, _09695_);
  nor _61198_ (_09720_, _09719_, _09694_);
  and _61199_ (_09721_, _05223_, _04800_);
  not _61200_ (_09722_, _09721_);
  and _61201_ (_09723_, _05901_, \oc8051_golden_model_1.PSW [4]);
  and _61202_ (_09724_, _05910_, \oc8051_golden_model_1.B [4]);
  nor _61203_ (_09725_, _09724_, _09723_);
  and _61204_ (_09726_, _05908_, \oc8051_golden_model_1.IP [4]);
  and _61205_ (_09727_, _05903_, \oc8051_golden_model_1.ACC [4]);
  nor _61206_ (_09728_, _09727_, _09726_);
  and _61207_ (_09729_, _09728_, _09725_);
  and _61208_ (_09730_, _05922_, \oc8051_golden_model_1.SCON [4]);
  and _61209_ (_09731_, _05924_, \oc8051_golden_model_1.IE [4]);
  nor _61210_ (_09732_, _09731_, _09730_);
  and _61211_ (_09733_, _05927_, \oc8051_golden_model_1.TCON [4]);
  and _61212_ (_09734_, _05929_, \oc8051_golden_model_1.P3INREG [4]);
  nor _61213_ (_09735_, _09734_, _09733_);
  and _61214_ (_09736_, _09735_, _09732_);
  and _61215_ (_09737_, _05916_, \oc8051_golden_model_1.P1INREG [4]);
  not _61216_ (_09738_, _09737_);
  and _61217_ (_09739_, _05209_, \oc8051_golden_model_1.P0INREG [4]);
  and _61218_ (_09740_, _05918_, \oc8051_golden_model_1.P2INREG [4]);
  nor _61219_ (_09741_, _09740_, _09739_);
  and _61220_ (_09742_, _09741_, _09738_);
  and _61221_ (_09743_, _09742_, _09736_);
  and _61222_ (_09744_, _09743_, _09729_);
  and _61223_ (_09745_, _09744_, _05778_);
  nor _61224_ (_09746_, _09745_, _09722_);
  nor _61225_ (_09747_, _05935_, _06094_);
  nor _61226_ (_09748_, _09747_, _09746_);
  and _61227_ (_09749_, _09748_, _09720_);
  not _61228_ (_09750_, _05224_);
  and _61229_ (_09751_, _05927_, \oc8051_golden_model_1.TCON [0]);
  and _61230_ (_09752_, _05910_, \oc8051_golden_model_1.B [0]);
  nor _61231_ (_09753_, _09752_, _09751_);
  and _61232_ (_09754_, _05901_, \oc8051_golden_model_1.PSW [0]);
  not _61233_ (_09755_, _09754_);
  and _61234_ (_09756_, _05908_, \oc8051_golden_model_1.IP [0]);
  and _61235_ (_09757_, _05903_, \oc8051_golden_model_1.ACC [0]);
  nor _61236_ (_09758_, _09757_, _09756_);
  and _61237_ (_09759_, _09758_, _09755_);
  and _61238_ (_09760_, _09759_, _09753_);
  and _61239_ (_09761_, _05922_, \oc8051_golden_model_1.SCON [0]);
  and _61240_ (_09762_, _05924_, \oc8051_golden_model_1.IE [0]);
  nor _61241_ (_09763_, _09762_, _09761_);
  and _61242_ (_09764_, _05916_, \oc8051_golden_model_1.P1INREG [0]);
  and _61243_ (_09765_, _05929_, \oc8051_golden_model_1.P3INREG [0]);
  nor _61244_ (_09766_, _09765_, _09764_);
  and _61245_ (_09767_, _05209_, \oc8051_golden_model_1.P0INREG [0]);
  and _61246_ (_09768_, _05918_, \oc8051_golden_model_1.P2INREG [0]);
  nor _61247_ (_09769_, _09768_, _09767_);
  and _61248_ (_09770_, _09769_, _09766_);
  and _61249_ (_09771_, _09770_, _09763_);
  and _61250_ (_09772_, _09771_, _09760_);
  and _61251_ (_09773_, _09772_, _05619_);
  nor _61252_ (_09774_, _09773_, _09750_);
  and _61253_ (_09775_, _05281_, _04800_);
  not _61254_ (_09776_, _09775_);
  and _61255_ (_09777_, _05927_, \oc8051_golden_model_1.TCON [6]);
  and _61256_ (_09778_, _05910_, \oc8051_golden_model_1.B [6]);
  nor _61257_ (_09779_, _09778_, _09777_);
  and _61258_ (_09780_, _05901_, \oc8051_golden_model_1.PSW [6]);
  not _61259_ (_09781_, _09780_);
  and _61260_ (_09782_, _05908_, \oc8051_golden_model_1.IP [6]);
  and _61261_ (_09783_, _05903_, \oc8051_golden_model_1.ACC [6]);
  nor _61262_ (_09784_, _09783_, _09782_);
  and _61263_ (_09785_, _09784_, _09781_);
  and _61264_ (_09786_, _09785_, _09779_);
  and _61265_ (_09787_, _05922_, \oc8051_golden_model_1.SCON [6]);
  and _61266_ (_09788_, _05924_, \oc8051_golden_model_1.IE [6]);
  nor _61267_ (_09789_, _09788_, _09787_);
  and _61268_ (_09790_, _05209_, \oc8051_golden_model_1.P0INREG [6]);
  and _61269_ (_09791_, _05918_, \oc8051_golden_model_1.P2INREG [6]);
  nor _61270_ (_09792_, _09791_, _09790_);
  and _61271_ (_09793_, _05916_, \oc8051_golden_model_1.P1INREG [6]);
  and _61272_ (_09794_, _05929_, \oc8051_golden_model_1.P3INREG [6]);
  nor _61273_ (_09795_, _09794_, _09793_);
  and _61274_ (_09796_, _09795_, _09792_);
  and _61275_ (_09797_, _09796_, _09789_);
  and _61276_ (_09798_, _09797_, _09786_);
  and _61277_ (_09799_, _09798_, _05364_);
  nor _61278_ (_09800_, _09799_, _09776_);
  nor _61279_ (_09801_, _09800_, _09774_);
  not _61280_ (_09802_, _05296_);
  and _61281_ (_09803_, _05901_, \oc8051_golden_model_1.PSW [3]);
  and _61282_ (_09804_, _05910_, \oc8051_golden_model_1.B [3]);
  nor _61283_ (_09805_, _09804_, _09803_);
  and _61284_ (_09806_, _05908_, \oc8051_golden_model_1.IP [3]);
  and _61285_ (_09807_, _05903_, \oc8051_golden_model_1.ACC [3]);
  nor _61286_ (_09808_, _09807_, _09806_);
  and _61287_ (_09809_, _09808_, _09805_);
  and _61288_ (_09810_, _05929_, \oc8051_golden_model_1.P3INREG [3]);
  not _61289_ (_09811_, _09810_);
  and _61290_ (_09812_, _05916_, \oc8051_golden_model_1.P1INREG [3]);
  and _61291_ (_09813_, _05918_, \oc8051_golden_model_1.P2INREG [3]);
  nor _61292_ (_09814_, _09813_, _09812_);
  and _61293_ (_09815_, _09814_, _09811_);
  and _61294_ (_09816_, _05922_, \oc8051_golden_model_1.SCON [3]);
  and _61295_ (_09817_, _05924_, \oc8051_golden_model_1.IE [3]);
  nor _61296_ (_09818_, _09817_, _09816_);
  and _61297_ (_09819_, _05927_, \oc8051_golden_model_1.TCON [3]);
  and _61298_ (_09820_, _05209_, \oc8051_golden_model_1.P0INREG [3]);
  nor _61299_ (_09821_, _09820_, _09819_);
  and _61300_ (_09822_, _09821_, _09818_);
  and _61301_ (_09823_, _09822_, _09815_);
  and _61302_ (_09824_, _09823_, _09809_);
  and _61303_ (_09825_, _09824_, _05519_);
  nor _61304_ (_09826_, _09825_, _09802_);
  and _61305_ (_09827_, _05215_, _04800_);
  not _61306_ (_09828_, _09827_);
  and _61307_ (_09829_, _05922_, \oc8051_golden_model_1.SCON [5]);
  and _61308_ (_09830_, _05924_, \oc8051_golden_model_1.IE [5]);
  nor _61309_ (_09831_, _09830_, _09829_);
  and _61310_ (_09832_, _05927_, \oc8051_golden_model_1.TCON [5]);
  and _61311_ (_09833_, _05929_, \oc8051_golden_model_1.P3INREG [5]);
  nor _61312_ (_09834_, _09833_, _09832_);
  and _61313_ (_09835_, _09834_, _09831_);
  and _61314_ (_09836_, _05908_, \oc8051_golden_model_1.IP [5]);
  and _61315_ (_09837_, _05903_, \oc8051_golden_model_1.ACC [5]);
  nor _61316_ (_09838_, _09837_, _09836_);
  and _61317_ (_09839_, _05901_, \oc8051_golden_model_1.PSW [5]);
  and _61318_ (_09840_, _05910_, \oc8051_golden_model_1.B [5]);
  nor _61319_ (_09841_, _09840_, _09839_);
  and _61320_ (_09842_, _09841_, _09838_);
  and _61321_ (_09843_, _05916_, \oc8051_golden_model_1.P1INREG [5]);
  and _61322_ (_09844_, _05918_, \oc8051_golden_model_1.P2INREG [5]);
  and _61323_ (_09845_, _05209_, \oc8051_golden_model_1.P0INREG [5]);
  or _61324_ (_09846_, _09845_, _09844_);
  nor _61325_ (_09847_, _09846_, _09843_);
  and _61326_ (_09848_, _09847_, _09842_);
  and _61327_ (_09849_, _09848_, _09835_);
  and _61328_ (_09850_, _09849_, _05470_);
  nor _61329_ (_09851_, _09850_, _09828_);
  nor _61330_ (_09852_, _09851_, _09826_);
  and _61331_ (_09853_, _09852_, _09801_);
  and _61332_ (_09854_, _09853_, _09749_);
  nor _61333_ (_09855_, _09854_, _09669_);
  not _61334_ (_09856_, _03604_);
  not _61335_ (_09857_, _08316_);
  nor _61336_ (_09858_, _08317_, _09857_);
  or _61337_ (_09859_, _09858_, _08273_);
  and _61338_ (_09860_, _09859_, _08315_);
  and _61339_ (_09861_, _08314_, _08289_);
  or _61340_ (_09862_, _09861_, _08250_);
  or _61341_ (_09863_, _09862_, _09860_);
  and _61342_ (_09864_, _08308_, _08296_);
  and _61343_ (_09865_, _08206_, _08191_);
  and _61344_ (_09866_, _09865_, _09864_);
  and _61345_ (_09867_, _09866_, _09863_);
  nor _61346_ (_09868_, _08295_, _08220_);
  nor _61347_ (_09869_, _09868_, _08219_);
  and _61348_ (_09870_, _09869_, _09865_);
  nor _61349_ (_09871_, _06133_, \oc8051_golden_model_1.ACC [7]);
  and _61350_ (_09872_, _08205_, _08191_);
  or _61351_ (_09873_, _09872_, _09871_);
  or _61352_ (_09874_, _09873_, _09870_);
  or _61353_ (_09875_, _09874_, _09867_);
  and _61354_ (_09876_, _09866_, _08320_);
  nor _61355_ (_09877_, _09876_, _04107_);
  and _61356_ (_09878_, _09877_, _09875_);
  and _61357_ (_09879_, _05964_, _05245_);
  or _61358_ (_09880_, _09879_, _09657_);
  or _61359_ (_09881_, _09880_, _04081_);
  not _61360_ (_09882_, _08089_);
  and _61361_ (_09883_, _05245_, \oc8051_golden_model_1.ACC [7]);
  or _61362_ (_09884_, _09883_, _09657_);
  and _61363_ (_09885_, _09884_, _04409_);
  nor _61364_ (_09886_, _04409_, _07871_);
  or _61365_ (_09887_, _09886_, _03610_);
  or _61366_ (_09888_, _09887_, _09885_);
  and _61367_ (_09889_, _09888_, _09882_);
  and _61368_ (_09890_, _09889_, _09881_);
  nor _61369_ (_09891_, _08099_, \oc8051_golden_model_1.PSW [7]);
  not _61370_ (_09892_, _09891_);
  nor _61371_ (_09893_, _09892_, _08109_);
  nor _61372_ (_09894_, _09893_, _09882_);
  nor _61373_ (_09895_, _03229_, _03215_);
  not _61374_ (_09896_, _09895_);
  nand _61375_ (_09897_, _09896_, _03730_);
  or _61376_ (_09898_, _09897_, _09894_);
  or _61377_ (_09899_, _09898_, _09890_);
  nor _61378_ (_09900_, _05901_, _07871_);
  and _61379_ (_09901_, _06095_, _05901_);
  or _61380_ (_09902_, _09901_, _09900_);
  or _61381_ (_09903_, _09902_, _04055_);
  or _61382_ (_09904_, _09666_, _03996_);
  and _61383_ (_09905_, _09904_, _09903_);
  and _61384_ (_09906_, _09905_, _09899_);
  or _61385_ (_09907_, _09906_, _03729_);
  or _61386_ (_09908_, _09884_, _03737_);
  nor _61387_ (_09909_, _03232_, _03215_);
  nor _61388_ (_09910_, _09909_, _03714_);
  and _61389_ (_09911_, _09910_, _09908_);
  and _61390_ (_09912_, _09911_, _09907_);
  and _61391_ (_09913_, _05952_, _05901_);
  or _61392_ (_09914_, _09913_, _09900_);
  and _61393_ (_09915_, _09914_, _03714_);
  or _61394_ (_09916_, _09915_, _09912_);
  nor _61395_ (_09917_, _03226_, _03219_);
  or _61396_ (_09918_, _09917_, _09916_);
  nor _61397_ (_09919_, _03511_, _03226_);
  not _61398_ (_09920_, _09919_);
  not _61399_ (_09921_, _09917_);
  nor _61400_ (_09922_, _05005_, _03756_);
  and _61401_ (_09923_, _04875_, _04800_);
  nor _61402_ (_09924_, _09923_, _09922_);
  and _61403_ (_09925_, _05005_, _03756_);
  nor _61404_ (_09926_, _04875_, _04800_);
  nor _61405_ (_09927_, _09926_, _09925_);
  and _61406_ (_09928_, _09927_, _09924_);
  and _61407_ (_09929_, _04406_, _03415_);
  and _61408_ (_09930_, _06764_, _03414_);
  and _61409_ (_09931_, _04620_, _04048_);
  or _61410_ (_09932_, _09931_, _09929_);
  nor _61411_ (_09933_, _09932_, _09930_);
  or _61412_ (_09934_, _09933_, _09929_);
  and _61413_ (_09935_, _09934_, _09928_);
  not _61414_ (_09936_, _09923_);
  nor _61415_ (_09937_, _09936_, _09922_);
  or _61416_ (_09938_, _09937_, _09925_);
  or _61417_ (_09939_, _09938_, _09935_);
  and _61418_ (_09940_, _05204_, _03454_);
  not _61419_ (_09941_, _09940_);
  and _61420_ (_09942_, _09941_, _05205_);
  and _61421_ (_09943_, _05363_, _03549_);
  nor _61422_ (_09944_, _05363_, _03549_);
  or _61423_ (_09945_, _09944_, _09943_);
  and _61424_ (_09946_, _09945_, _09942_);
  and _61425_ (_09947_, _05469_, _05226_);
  nor _61426_ (_09948_, _05469_, _05226_);
  nor _61427_ (_09949_, _09948_, _09947_);
  and _61428_ (_09950_, _05777_, _03486_);
  nor _61429_ (_09951_, _05777_, _03486_);
  or _61430_ (_09952_, _09951_, _09950_);
  and _61431_ (_09953_, _09952_, _09949_);
  and _61432_ (_09954_, _09953_, _09946_);
  and _61433_ (_09955_, _09954_, _09939_);
  and _61434_ (_09956_, _05777_, _05218_);
  and _61435_ (_09957_, _09949_, _09956_);
  or _61436_ (_09958_, _09957_, _09947_);
  and _61437_ (_09959_, _09958_, _09946_);
  and _61438_ (_09960_, _05363_, _05112_);
  and _61439_ (_09961_, _09942_, _09960_);
  or _61440_ (_09962_, _09961_, _09940_);
  or _61441_ (_09963_, _09962_, _09959_);
  nor _61442_ (_09964_, _09963_, _09955_);
  and _61443_ (_09965_, _04634_, _04188_);
  not _61444_ (_09966_, _09965_);
  and _61445_ (_09967_, _09933_, _09928_);
  and _61446_ (_09968_, _09967_, _09966_);
  and _61447_ (_09969_, _09968_, _09954_);
  nor _61448_ (_09970_, _09969_, _09964_);
  or _61449_ (_09971_, _09970_, _09921_);
  and _61450_ (_09972_, _09971_, _09920_);
  and _61451_ (_09973_, _09972_, _09918_);
  or _61452_ (_09974_, _06592_, _03581_);
  or _61453_ (_09975_, _06637_, _03904_);
  or _61454_ (_09976_, _08636_, _03756_);
  and _61455_ (_09977_, _09976_, _09974_);
  not _61456_ (_09978_, _09977_);
  or _61457_ (_09979_, _09978_, _09975_);
  nand _61458_ (_09980_, _09979_, _09974_);
  nor _61459_ (_09981_, _06501_, _03414_);
  nand _61460_ (_09982_, _06501_, _03414_);
  and _61461_ (_09983_, _06546_, _04048_);
  nor _61462_ (_09984_, _09983_, _09981_);
  and _61463_ (_09985_, _09984_, _09982_);
  or _61464_ (_09986_, _09985_, _09981_);
  nand _61465_ (_09987_, _06637_, _03904_);
  and _61466_ (_09988_, _09987_, _09977_);
  and _61467_ (_09989_, _09988_, _09975_);
  and _61468_ (_09990_, _09989_, _09986_);
  or _61469_ (_09991_, _09990_, _09980_);
  nand _61470_ (_09992_, _06455_, _03549_);
  or _61471_ (_09993_, _06455_, _03549_);
  nor _61472_ (_09994_, _06069_, _03446_);
  nor _61473_ (_09995_, _09994_, _06150_);
  and _61474_ (_09996_, _09995_, _09993_);
  and _61475_ (_09997_, _09996_, _09992_);
  nor _61476_ (_09998_, _06730_, _03486_);
  not _61477_ (_09999_, _09998_);
  nand _61478_ (_10000_, _06684_, _03860_);
  and _61479_ (_10001_, _10000_, _09999_);
  nor _61480_ (_10002_, _06684_, _03860_);
  and _61481_ (_10003_, _06730_, _03486_);
  nor _61482_ (_10004_, _10003_, _10002_);
  and _61483_ (_10005_, _10004_, _10001_);
  and _61484_ (_10006_, _10005_, _09997_);
  and _61485_ (_10007_, _10006_, _09991_);
  or _61486_ (_10008_, _09998_, _10002_);
  and _61487_ (_10009_, _09997_, _10008_);
  and _61488_ (_10010_, _10009_, _10000_);
  nor _61489_ (_10011_, _09993_, _06150_);
  or _61490_ (_10012_, _10011_, _09994_);
  or _61491_ (_10013_, _10012_, _10010_);
  or _61492_ (_10014_, _10013_, _10007_);
  or _61493_ (_10015_, _06546_, _04048_);
  and _61494_ (_10016_, _09989_, _09985_);
  and _61495_ (_10017_, _10016_, _10015_);
  nand _61496_ (_10018_, _10017_, _10006_);
  and _61497_ (_10019_, _10018_, _09919_);
  and _61498_ (_10020_, _10019_, _10014_);
  or _61499_ (_10021_, _10020_, _09973_);
  and _61500_ (_10022_, _10021_, _04107_);
  or _61501_ (_10023_, _10022_, _09878_);
  and _61502_ (_10024_, _10023_, _09856_);
  nor _61503_ (_10025_, _03226_, _03215_);
  nor _61504_ (_10026_, _08740_, _08739_);
  nor _61505_ (_10027_, _10026_, _08743_);
  nor _61506_ (_10028_, _08738_, _08407_);
  and _61507_ (_10029_, _10028_, _10027_);
  nor _61508_ (_10030_, _08744_, _08745_);
  nor _61509_ (_10031_, _10030_, _08748_);
  nor _61510_ (_10032_, _03414_, \oc8051_golden_model_1.ACC [1]);
  and _61511_ (_10033_, _03414_, \oc8051_golden_model_1.ACC [1]);
  and _61512_ (_10034_, _04048_, \oc8051_golden_model_1.ACC [0]);
  nor _61513_ (_10035_, _10034_, _10033_);
  or _61514_ (_10036_, _10035_, _10032_);
  and _61515_ (_10037_, _10036_, _10031_);
  nand _61516_ (_10038_, _03581_, \oc8051_golden_model_1.ACC [3]);
  nor _61517_ (_10039_, _03581_, \oc8051_golden_model_1.ACC [3]);
  nor _61518_ (_10040_, _03904_, \oc8051_golden_model_1.ACC [2]);
  or _61519_ (_10041_, _10040_, _10039_);
  and _61520_ (_10042_, _10041_, _10038_);
  or _61521_ (_10043_, _10042_, _10037_);
  and _61522_ (_10044_, _10043_, _10029_);
  nand _61523_ (_10045_, _03860_, \oc8051_golden_model_1.ACC [5]);
  nor _61524_ (_10046_, _03860_, \oc8051_golden_model_1.ACC [5]);
  nor _61525_ (_10047_, _03486_, \oc8051_golden_model_1.ACC [4]);
  or _61526_ (_10048_, _10047_, _10046_);
  and _61527_ (_10049_, _10048_, _10045_);
  and _61528_ (_10050_, _10049_, _10028_);
  nor _61529_ (_10051_, _03446_, \oc8051_golden_model_1.ACC [7]);
  or _61530_ (_10052_, _03549_, \oc8051_golden_model_1.ACC [6]);
  nor _61531_ (_10053_, _10052_, _08407_);
  or _61532_ (_10054_, _10053_, _10051_);
  or _61533_ (_10055_, _10054_, _10050_);
  or _61534_ (_10056_, _10055_, _10044_);
  and _61535_ (_10057_, _04048_, _03335_);
  nor _61536_ (_10058_, _10057_, _08751_);
  nor _61537_ (_10059_, _08753_, _10058_);
  and _61538_ (_10060_, _10059_, _10031_);
  and _61539_ (_10061_, _10060_, _10029_);
  nor _61540_ (_10062_, _10061_, _09856_);
  and _61541_ (_10063_, _10062_, _10056_);
  or _61542_ (_10064_, _10063_, _10025_);
  or _61543_ (_10065_, _10064_, _10024_);
  nand _61544_ (_10066_, _10025_, \oc8051_golden_model_1.PSW [7]);
  and _61545_ (_10067_, _10066_, _06840_);
  and _61546_ (_10068_, _10067_, _10065_);
  or _61547_ (_10069_, _09900_, _06138_);
  and _61548_ (_10070_, _09902_, _03719_);
  and _61549_ (_10071_, _10070_, _10069_);
  nor _61550_ (_10072_, _10071_, _10068_);
  nor _61551_ (_10073_, _10072_, _03718_);
  and _61552_ (_10074_, _05918_, \oc8051_golden_model_1.P2 [2]);
  and _61553_ (_10075_, _05929_, \oc8051_golden_model_1.P3 [2]);
  nor _61554_ (_10076_, _10075_, _10074_);
  and _61555_ (_10077_, _05209_, \oc8051_golden_model_1.P0 [2]);
  and _61556_ (_10078_, _05916_, \oc8051_golden_model_1.P1 [2]);
  nor _61557_ (_10079_, _10078_, _10077_);
  and _61558_ (_10080_, _10079_, _10076_);
  and _61559_ (_10081_, _10080_, _09683_);
  and _61560_ (_10082_, _10081_, _09680_);
  and _61561_ (_10083_, _10082_, _05668_);
  nor _61562_ (_10084_, _10083_, _09670_);
  and _61563_ (_10085_, _05209_, \oc8051_golden_model_1.P0 [1]);
  and _61564_ (_10086_, _05916_, \oc8051_golden_model_1.P1 [1]);
  nor _61565_ (_10087_, _10086_, _10085_);
  and _61566_ (_10088_, _05929_, \oc8051_golden_model_1.P3 [1]);
  and _61567_ (_10089_, _05918_, \oc8051_golden_model_1.P2 [1]);
  or _61568_ (_10090_, _10089_, _10088_);
  nor _61569_ (_10091_, _10090_, _09712_);
  and _61570_ (_10092_, _10091_, _09702_);
  and _61571_ (_10093_, _10092_, _09711_);
  and _61572_ (_10094_, _10093_, _10087_);
  and _61573_ (_10095_, _10094_, _05568_);
  nor _61574_ (_10096_, _10095_, _09695_);
  nor _61575_ (_10097_, _10096_, _10084_);
  and _61576_ (_10098_, _05929_, \oc8051_golden_model_1.P3 [4]);
  not _61577_ (_10099_, _10098_);
  and _61578_ (_10100_, _05918_, \oc8051_golden_model_1.P2 [4]);
  nor _61579_ (_10101_, _10100_, _09733_);
  and _61580_ (_10102_, _10101_, _10099_);
  and _61581_ (_10103_, _05209_, \oc8051_golden_model_1.P0 [4]);
  and _61582_ (_10104_, _05916_, \oc8051_golden_model_1.P1 [4]);
  nor _61583_ (_10105_, _10104_, _10103_);
  and _61584_ (_10106_, _10105_, _09732_);
  and _61585_ (_10107_, _10106_, _10102_);
  and _61586_ (_10108_, _10107_, _09729_);
  and _61587_ (_10109_, _10108_, _05778_);
  nor _61588_ (_10110_, _09722_, _10109_);
  nor _61589_ (_10111_, _10110_, _06137_);
  and _61590_ (_10112_, _10111_, _10097_);
  and _61591_ (_10113_, _05918_, \oc8051_golden_model_1.P2 [0]);
  and _61592_ (_10114_, _05929_, \oc8051_golden_model_1.P3 [0]);
  nor _61593_ (_10115_, _10114_, _10113_);
  and _61594_ (_10116_, _05209_, \oc8051_golden_model_1.P0 [0]);
  and _61595_ (_10117_, _05916_, \oc8051_golden_model_1.P1 [0]);
  nor _61596_ (_10118_, _10117_, _10116_);
  and _61597_ (_10119_, _10118_, _10115_);
  and _61598_ (_10120_, _10119_, _09763_);
  and _61599_ (_10121_, _10120_, _09760_);
  and _61600_ (_10122_, _10121_, _05619_);
  nor _61601_ (_10123_, _10122_, _09750_);
  and _61602_ (_10124_, _05918_, \oc8051_golden_model_1.P2 [6]);
  and _61603_ (_10125_, _05929_, \oc8051_golden_model_1.P3 [6]);
  nor _61604_ (_10126_, _10125_, _10124_);
  and _61605_ (_10127_, _05209_, \oc8051_golden_model_1.P0 [6]);
  and _61606_ (_10128_, _05916_, \oc8051_golden_model_1.P1 [6]);
  nor _61607_ (_10129_, _10128_, _10127_);
  and _61608_ (_10130_, _10129_, _10126_);
  and _61609_ (_10131_, _10130_, _09789_);
  and _61610_ (_10132_, _10131_, _09786_);
  and _61611_ (_10133_, _10132_, _05364_);
  nor _61612_ (_10134_, _09776_, _10133_);
  nor _61613_ (_10135_, _10134_, _10123_);
  and _61614_ (_10136_, _05209_, \oc8051_golden_model_1.P0 [3]);
  and _61615_ (_10137_, _05916_, \oc8051_golden_model_1.P1 [3]);
  nor _61616_ (_10138_, _10137_, _10136_);
  and _61617_ (_10139_, _05929_, \oc8051_golden_model_1.P3 [3]);
  and _61618_ (_10140_, _05918_, \oc8051_golden_model_1.P2 [3]);
  or _61619_ (_10141_, _10140_, _10139_);
  nor _61620_ (_10142_, _10141_, _09819_);
  and _61621_ (_10143_, _10142_, _09809_);
  and _61622_ (_10144_, _10143_, _09818_);
  and _61623_ (_10145_, _10144_, _10138_);
  and _61624_ (_10146_, _10145_, _05519_);
  nor _61625_ (_10147_, _10146_, _09802_);
  and _61626_ (_10148_, _05209_, \oc8051_golden_model_1.P0 [5]);
  and _61627_ (_10149_, _05916_, \oc8051_golden_model_1.P1 [5]);
  nor _61628_ (_10150_, _10149_, _10148_);
  and _61629_ (_10151_, _05929_, \oc8051_golden_model_1.P3 [5]);
  and _61630_ (_10152_, _05918_, \oc8051_golden_model_1.P2 [5]);
  or _61631_ (_10153_, _10152_, _10151_);
  nor _61632_ (_10154_, _10153_, _09832_);
  and _61633_ (_10155_, _10154_, _09842_);
  and _61634_ (_10156_, _10155_, _09831_);
  and _61635_ (_10157_, _10156_, _10150_);
  and _61636_ (_10158_, _10157_, _05470_);
  nor _61637_ (_10159_, _09828_, _10158_);
  nor _61638_ (_10160_, _10159_, _10147_);
  and _61639_ (_10161_, _10160_, _10135_);
  and _61640_ (_10162_, _10161_, _10112_);
  and _61641_ (_10163_, _03718_, \oc8051_golden_model_1.PSW [7]);
  and _61642_ (_10164_, _10163_, _10162_);
  or _61643_ (_10165_, _10164_, _10073_);
  nor _61644_ (_10166_, _06869_, _03753_);
  and _61645_ (_10167_, _10166_, _10165_);
  or _61646_ (_10168_, _10167_, _09855_);
  and _61647_ (_10169_, _10168_, _09668_);
  not _61648_ (_10170_, _08058_);
  or _61649_ (_10171_, _10162_, \oc8051_golden_model_1.PSW [7]);
  and _61650_ (_10172_, _10171_, _03752_);
  or _61651_ (_10173_, _10172_, _10170_);
  or _61652_ (_10174_, _10173_, _10169_);
  and _61653_ (_10175_, _07835_, _06762_);
  and _61654_ (_10176_, _10175_, _06771_);
  and _61655_ (_10177_, _07830_, _07826_);
  nor _61656_ (_10178_, _10177_, _07824_);
  not _61657_ (_10179_, _10178_);
  and _61658_ (_10180_, _07832_, _07826_);
  not _61659_ (_10181_, _10180_);
  nor _61660_ (_10182_, _10181_, _08175_);
  nor _61661_ (_10183_, _10182_, _10179_);
  or _61662_ (_10184_, _10183_, _10176_);
  and _61663_ (_10185_, _10184_, _08054_);
  or _61664_ (_10186_, _10185_, _08059_);
  and _61665_ (_10187_, _10186_, _10174_);
  and _61666_ (_10188_, _10184_, _08053_);
  or _61667_ (_10189_, _10188_, _08051_);
  or _61668_ (_10190_, _10189_, _10187_);
  and _61669_ (_10191_, _07997_, _07992_);
  nor _61670_ (_10192_, _10191_, _07990_);
  not _61671_ (_10193_, _10192_);
  and _61672_ (_10194_, _08479_, _07992_);
  not _61673_ (_10195_, _10194_);
  nor _61674_ (_10196_, _10195_, _08045_);
  nor _61675_ (_10197_, _10196_, _10193_);
  and _61676_ (_10198_, _08000_, _06684_);
  and _61677_ (_10199_, _10198_, _06455_);
  and _61678_ (_10200_, _10199_, _06069_);
  not _61679_ (_10201_, _08051_);
  or _61680_ (_10202_, _10201_, _10200_);
  or _61681_ (_10203_, _10202_, _10197_);
  and _61682_ (_10204_, _10203_, _10190_);
  or _61683_ (_10205_, _10204_, _03761_);
  and _61684_ (_10206_, _08534_, _08532_);
  nand _61685_ (_10207_, _10206_, _08509_);
  nor _61686_ (_10208_, _10207_, _06133_);
  and _61687_ (_10209_, _08530_, _08525_);
  nor _61688_ (_10210_, _10209_, _08523_);
  nor _61689_ (_10211_, _08544_, _08539_);
  nor _61690_ (_10212_, _10211_, _08538_);
  and _61691_ (_10213_, _08531_, _08525_);
  nand _61692_ (_10214_, _10213_, _10212_);
  and _61693_ (_10215_, _10214_, _10210_);
  and _61694_ (_10216_, _08558_, _08552_);
  and _61695_ (_10217_, _08566_, _03335_);
  nor _61696_ (_10218_, _10217_, _08562_);
  or _61697_ (_10219_, _10218_, _08563_);
  and _61698_ (_10220_, _10219_, _10216_);
  and _61699_ (_10221_, _08556_, _08552_);
  or _61700_ (_10222_, _10221_, _08550_);
  nor _61701_ (_10223_, _10222_, _10220_);
  and _61702_ (_10224_, _08546_, _08540_);
  nand _61703_ (_10225_, _10213_, _10224_);
  or _61704_ (_10226_, _10225_, _10223_);
  and _61705_ (_10227_, _10226_, _10215_);
  or _61706_ (_10228_, _10227_, _10208_);
  or _61707_ (_10229_, _10228_, _03766_);
  and _61708_ (_10230_, _10229_, _07914_);
  and _61709_ (_10231_, _10230_, _10205_);
  and _61710_ (_10232_, _07916_, _05247_);
  and _61711_ (_10233_, _07927_, _07924_);
  nor _61712_ (_10234_, _10233_, _07922_);
  not _61713_ (_10235_, _10234_);
  and _61714_ (_10236_, _08591_, _07924_);
  not _61715_ (_10237_, _10236_);
  nor _61716_ (_10238_, _10237_, _07979_);
  nor _61717_ (_10239_, _10238_, _10235_);
  or _61718_ (_10240_, _10239_, _10232_);
  and _61719_ (_10241_, _10240_, _07913_);
  or _61720_ (_10242_, _10241_, _07390_);
  or _61721_ (_10243_, _10242_, _10231_);
  and _61722_ (_10244_, _10243_, _09667_);
  or _61723_ (_10245_, _10244_, _04481_);
  and _61724_ (_10246_, _06069_, _05245_);
  or _61725_ (_10247_, _09657_, _07400_);
  or _61726_ (_10248_, _10247_, _10246_);
  and _61727_ (_10249_, _10248_, _03589_);
  and _61728_ (_10250_, _10249_, _10245_);
  or _61729_ (_10251_, _10250_, _09664_);
  nor _61730_ (_10252_, _07405_, _03585_);
  and _61731_ (_10253_, _10252_, _10251_);
  nor _61732_ (_10254_, _10162_, _07871_);
  and _61733_ (_10255_, _10254_, _03585_);
  or _61734_ (_10256_, _10255_, _03601_);
  or _61735_ (_10257_, _10256_, _10253_);
  and _61736_ (_10258_, _06171_, _05245_);
  or _61737_ (_10259_, _10258_, _09657_);
  or _61738_ (_10260_, _10259_, _05886_);
  and _61739_ (_10261_, _10260_, _10257_);
  or _61740_ (_10262_, _10261_, _03584_);
  not _61741_ (_10263_, _03584_);
  nand _61742_ (_10264_, _10162_, _07871_);
  or _61743_ (_10265_, _10264_, _10263_);
  and _61744_ (_10266_, _10265_, _10262_);
  or _61745_ (_10267_, _10266_, _03600_);
  and _61746_ (_10268_, _05884_, _05245_);
  or _61747_ (_10269_, _10268_, _09657_);
  or _61748_ (_10270_, _10269_, _07766_);
  and _61749_ (_10271_, _10270_, _07778_);
  and _61750_ (_10272_, _10271_, _10267_);
  or _61751_ (_10273_, _10272_, _09660_);
  and _61752_ (_10274_, _10273_, _07777_);
  or _61753_ (_10275_, _09657_, _05310_);
  and _61754_ (_10276_, _10259_, _03622_);
  and _61755_ (_10277_, _10276_, _10275_);
  or _61756_ (_10278_, _10277_, _10274_);
  and _61757_ (_10279_, _10278_, _06828_);
  and _61758_ (_10280_, _09884_, _03790_);
  and _61759_ (_10281_, _10280_, _10275_);
  or _61760_ (_10282_, _10281_, _03624_);
  or _61761_ (_10283_, _10282_, _10279_);
  nor _61762_ (_10284_, _05882_, _09661_);
  or _61763_ (_10285_, _09657_, _07795_);
  or _61764_ (_10286_, _10285_, _10284_);
  and _61765_ (_10287_, _10286_, _07793_);
  and _61766_ (_10288_, _10287_, _10283_);
  nor _61767_ (_10289_, _06377_, _09661_);
  or _61768_ (_10290_, _10289_, _09657_);
  and _61769_ (_10291_, _10290_, _03785_);
  or _61770_ (_10292_, _10291_, _08468_);
  or _61771_ (_10293_, _10292_, _10288_);
  nor _61772_ (_10294_, _07823_, _06075_);
  or _61773_ (_10295_, _10294_, _07888_);
  or _61774_ (_10296_, _10295_, _10176_);
  or _61775_ (_10297_, _10296_, _07898_);
  and _61776_ (_10298_, _10297_, _10293_);
  or _61777_ (_10299_, _10298_, _08475_);
  nor _61778_ (_10300_, _07989_, _06075_);
  or _61779_ (_10301_, _10300_, _08500_);
  or _61780_ (_10302_, _08477_, _10200_);
  or _61781_ (_10303_, _10302_, _10301_);
  and _61782_ (_10304_, _10303_, _03777_);
  and _61783_ (_10305_, _10304_, _10299_);
  nor _61784_ (_10306_, _08522_, _06075_);
  or _61785_ (_10307_, _10306_, _08581_);
  or _61786_ (_10308_, _10307_, _10208_);
  and _61787_ (_10309_, _10308_, _03776_);
  or _61788_ (_10310_, _10309_, _08506_);
  or _61789_ (_10311_, _10310_, _10305_);
  nor _61790_ (_10312_, _07921_, _06075_);
  or _61791_ (_10313_, _10312_, _08611_);
  or _61792_ (_10314_, _10232_, _08589_);
  or _61793_ (_10315_, _10314_, _10313_);
  and _61794_ (_10316_, _10315_, _08588_);
  and _61795_ (_10317_, _10316_, _10311_);
  nor _61796_ (_10318_, _08070_, _03949_);
  and _61797_ (_10319_, _04474_, _03202_);
  nor _61798_ (_10320_, _10319_, _10318_);
  nor _61799_ (_10321_, _04488_, _04066_);
  or _61800_ (_10322_, _10321_, _03949_);
  nand _61801_ (_10323_, _10322_, _10320_);
  and _61802_ (_10324_, _08587_, \oc8051_golden_model_1.ACC [7]);
  or _61803_ (_10325_, _10324_, _10323_);
  or _61804_ (_10326_, _10325_, _10317_);
  and _61805_ (_10327_, _04058_, _03202_);
  not _61806_ (_10328_, _10327_);
  nor _61807_ (_10329_, _08662_, _08375_);
  not _61808_ (_10330_, _10329_);
  or _61809_ (_10331_, _10330_, _08692_);
  and _61810_ (_10332_, _10331_, _08451_);
  and _61811_ (_10333_, _10332_, _10328_);
  or _61812_ (_10334_, _10333_, _08617_);
  and _61813_ (_10335_, _10334_, _10326_);
  and _61814_ (_10336_, _10332_, _10327_);
  or _61815_ (_10337_, _10336_, _08620_);
  or _61816_ (_10338_, _10337_, _10335_);
  and _61817_ (_10339_, _08656_, _08400_);
  nor _61818_ (_10340_, _08625_, _08399_);
  nor _61819_ (_10341_, _10340_, _08398_);
  or _61820_ (_10342_, _10341_, _08624_);
  or _61821_ (_10343_, _10342_, _10339_);
  and _61822_ (_10344_, _10343_, _08702_);
  and _61823_ (_10345_, _10344_, _10338_);
  not _61824_ (_10346_, _08406_);
  not _61825_ (_10347_, _08405_);
  nand _61826_ (_10348_, _08765_, _10347_);
  and _61827_ (_10349_, _10348_, _08701_);
  and _61828_ (_10350_, _10349_, _10346_);
  or _61829_ (_10351_, _10350_, _03815_);
  not _61830_ (_10352_, _08189_);
  nand _61831_ (_10353_, _08725_, _10352_);
  and _61832_ (_10354_, _10353_, _03517_);
  nor _61833_ (_10355_, _08701_, _08188_);
  and _61834_ (_10356_, _10355_, _10354_);
  or _61835_ (_10357_, _10356_, _10351_);
  or _61836_ (_10358_, _10357_, _10345_);
  not _61837_ (_10359_, _08780_);
  or _61838_ (_10360_, _09880_, _04246_);
  and _61839_ (_10361_, _10360_, _10359_);
  and _61840_ (_10362_, _10361_, _10358_);
  or _61841_ (_10363_, _10362_, _09656_);
  and _61842_ (_10364_, _10363_, _03823_);
  and _61843_ (_10365_, _09914_, _03453_);
  or _61844_ (_10366_, _10365_, _03447_);
  or _61845_ (_10367_, _10366_, _10364_);
  and _61846_ (_10368_, _05831_, _05245_);
  or _61847_ (_10369_, _09657_, _03514_);
  or _61848_ (_10370_, _10369_, _10368_);
  and _61849_ (_10371_, _10370_, _10367_);
  or _61850_ (_10372_, _10371_, _43004_);
  or _61851_ (_10373_, _43000_, \oc8051_golden_model_1.PSW [7]);
  and _61852_ (_10374_, _10373_, _41806_);
  and _61853_ (_40578_, _10374_, _10372_);
  not _61854_ (_10375_, \oc8051_golden_model_1.PCON [7]);
  nor _61855_ (_10376_, _05212_, _10375_);
  not _61856_ (_10377_, _05212_);
  nor _61857_ (_10378_, _06377_, _10377_);
  nor _61858_ (_10379_, _10378_, _10376_);
  nor _61859_ (_10380_, _10379_, _07793_);
  and _61860_ (_10381_, _06171_, _05212_);
  nor _61861_ (_10382_, _10381_, _10376_);
  and _61862_ (_10383_, _10382_, _03601_);
  nor _61863_ (_10384_, _10377_, _05204_);
  nor _61864_ (_10385_, _10384_, _10376_);
  and _61865_ (_10386_, _10385_, _07390_);
  and _61866_ (_10387_, _05212_, \oc8051_golden_model_1.ACC [7]);
  nor _61867_ (_10388_, _10387_, _10376_);
  nor _61868_ (_10389_, _10388_, _03737_);
  nor _61869_ (_10390_, _10388_, _09029_);
  nor _61870_ (_10391_, _04409_, _10375_);
  or _61871_ (_10392_, _10391_, _10390_);
  and _61872_ (_10393_, _10392_, _04081_);
  and _61873_ (_10394_, _05964_, _05212_);
  nor _61874_ (_10395_, _10394_, _10376_);
  nor _61875_ (_10396_, _10395_, _04081_);
  or _61876_ (_10397_, _10396_, _10393_);
  and _61877_ (_10398_, _10397_, _03996_);
  nor _61878_ (_10399_, _10385_, _03996_);
  nor _61879_ (_10400_, _10399_, _10398_);
  nor _61880_ (_10401_, _10400_, _03729_);
  or _61881_ (_10402_, _10401_, _07390_);
  nor _61882_ (_10403_, _10402_, _10389_);
  nor _61883_ (_10404_, _10403_, _10386_);
  nor _61884_ (_10405_, _10404_, _04481_);
  and _61885_ (_10406_, _06069_, _05212_);
  nor _61886_ (_10407_, _10376_, _07400_);
  not _61887_ (_10408_, _10407_);
  nor _61888_ (_10409_, _10408_, _10406_);
  or _61889_ (_10410_, _10409_, _03222_);
  nor _61890_ (_10411_, _10410_, _10405_);
  nor _61891_ (_10412_, _06363_, _10377_);
  nor _61892_ (_10413_, _10412_, _10376_);
  nor _61893_ (_10414_, _10413_, _03589_);
  or _61894_ (_10415_, _10414_, _03601_);
  nor _61895_ (_10416_, _10415_, _10411_);
  nor _61896_ (_10417_, _10416_, _10383_);
  or _61897_ (_10418_, _10417_, _03600_);
  and _61898_ (_10419_, _05884_, _05212_);
  or _61899_ (_10420_, _10419_, _10376_);
  or _61900_ (_10421_, _10420_, _07766_);
  and _61901_ (_10422_, _10421_, _07778_);
  and _61902_ (_10423_, _10422_, _10418_);
  and _61903_ (_10424_, _06378_, _05212_);
  nor _61904_ (_10425_, _10424_, _10376_);
  nor _61905_ (_10426_, _10425_, _07778_);
  nor _61906_ (_10427_, _10426_, _10423_);
  nor _61907_ (_10428_, _10427_, _03622_);
  nor _61908_ (_10429_, _10376_, _05310_);
  not _61909_ (_10430_, _10429_);
  nor _61910_ (_10431_, _10382_, _07777_);
  and _61911_ (_10432_, _10431_, _10430_);
  nor _61912_ (_10433_, _10432_, _10428_);
  nor _61913_ (_10434_, _10433_, _03790_);
  nor _61914_ (_10435_, _10388_, _06828_);
  and _61915_ (_10436_, _10435_, _10430_);
  or _61916_ (_10437_, _10436_, _10434_);
  and _61917_ (_10438_, _10437_, _07795_);
  nor _61918_ (_10439_, _05882_, _10377_);
  nor _61919_ (_10440_, _10439_, _10376_);
  nor _61920_ (_10441_, _10440_, _07795_);
  or _61921_ (_10442_, _10441_, _10438_);
  and _61922_ (_10443_, _10442_, _07793_);
  nor _61923_ (_10444_, _10443_, _10380_);
  nor _61924_ (_10445_, _10444_, _03815_);
  nor _61925_ (_10446_, _10395_, _04246_);
  or _61926_ (_10447_, _10446_, _03447_);
  nor _61927_ (_10448_, _10447_, _10445_);
  and _61928_ (_10449_, _05831_, _05212_);
  or _61929_ (_10450_, _10376_, _03514_);
  nor _61930_ (_10451_, _10450_, _10449_);
  nor _61931_ (_10452_, _10451_, _10448_);
  or _61932_ (_10453_, _10452_, _43004_);
  or _61933_ (_10454_, _43000_, \oc8051_golden_model_1.PCON [7]);
  and _61934_ (_10455_, _10454_, _41806_);
  and _61935_ (_40579_, _10455_, _10453_);
  not _61936_ (_10456_, \oc8051_golden_model_1.SBUF [7]);
  nor _61937_ (_10457_, _05221_, _10456_);
  not _61938_ (_10458_, _05221_);
  nor _61939_ (_10459_, _06377_, _10458_);
  nor _61940_ (_10460_, _10459_, _10457_);
  nor _61941_ (_10461_, _10460_, _07793_);
  and _61942_ (_10462_, _06171_, _05221_);
  nor _61943_ (_10463_, _10462_, _10457_);
  and _61944_ (_10464_, _10463_, _03601_);
  and _61945_ (_10465_, _05221_, \oc8051_golden_model_1.ACC [7]);
  nor _61946_ (_10466_, _10465_, _10457_);
  nor _61947_ (_10467_, _10466_, _03737_);
  nor _61948_ (_10468_, _10466_, _09029_);
  nor _61949_ (_10469_, _04409_, _10456_);
  or _61950_ (_10470_, _10469_, _10468_);
  and _61951_ (_10471_, _10470_, _04081_);
  and _61952_ (_10472_, _05964_, _05221_);
  nor _61953_ (_10473_, _10472_, _10457_);
  nor _61954_ (_10474_, _10473_, _04081_);
  or _61955_ (_10475_, _10474_, _10471_);
  and _61956_ (_10476_, _10475_, _03996_);
  nor _61957_ (_10477_, _10458_, _05204_);
  nor _61958_ (_10478_, _10477_, _10457_);
  nor _61959_ (_10479_, _10478_, _03996_);
  nor _61960_ (_10480_, _10479_, _10476_);
  nor _61961_ (_10481_, _10480_, _03729_);
  or _61962_ (_10482_, _10481_, _07390_);
  nor _61963_ (_10483_, _10482_, _10467_);
  and _61964_ (_10484_, _10478_, _07390_);
  nor _61965_ (_10485_, _10484_, _10483_);
  nor _61966_ (_10486_, _10485_, _04481_);
  and _61967_ (_10487_, _06069_, _05221_);
  nor _61968_ (_10488_, _10457_, _07400_);
  not _61969_ (_10489_, _10488_);
  nor _61970_ (_10490_, _10489_, _10487_);
  or _61971_ (_10491_, _10490_, _03222_);
  nor _61972_ (_10492_, _10491_, _10486_);
  nor _61973_ (_10493_, _06363_, _10458_);
  nor _61974_ (_10494_, _10493_, _10457_);
  nor _61975_ (_10495_, _10494_, _03589_);
  or _61976_ (_10496_, _10495_, _03601_);
  nor _61977_ (_10497_, _10496_, _10492_);
  nor _61978_ (_10498_, _10497_, _10464_);
  or _61979_ (_10499_, _10498_, _03600_);
  and _61980_ (_10500_, _05884_, _05221_);
  or _61981_ (_10501_, _10500_, _10457_);
  or _61982_ (_10502_, _10501_, _07766_);
  and _61983_ (_10503_, _10502_, _07778_);
  and _61984_ (_10504_, _10503_, _10499_);
  and _61985_ (_10505_, _06378_, _05221_);
  nor _61986_ (_10506_, _10505_, _10457_);
  nor _61987_ (_10507_, _10506_, _07778_);
  nor _61988_ (_10508_, _10507_, _10504_);
  nor _61989_ (_10509_, _10508_, _03622_);
  nor _61990_ (_10510_, _10457_, _05310_);
  not _61991_ (_10511_, _10510_);
  nor _61992_ (_10512_, _10463_, _07777_);
  and _61993_ (_10513_, _10512_, _10511_);
  nor _61994_ (_10514_, _10513_, _10509_);
  nor _61995_ (_10515_, _10514_, _03790_);
  nor _61996_ (_10516_, _10466_, _06828_);
  and _61997_ (_10517_, _10516_, _10511_);
  or _61998_ (_10518_, _10517_, _10515_);
  and _61999_ (_10519_, _10518_, _07795_);
  nor _62000_ (_10520_, _05882_, _10458_);
  nor _62001_ (_10521_, _10520_, _10457_);
  nor _62002_ (_10522_, _10521_, _07795_);
  or _62003_ (_10523_, _10522_, _10519_);
  and _62004_ (_10524_, _10523_, _07793_);
  nor _62005_ (_10525_, _10524_, _10461_);
  nor _62006_ (_10526_, _10525_, _03815_);
  nor _62007_ (_10527_, _10473_, _04246_);
  or _62008_ (_10528_, _10527_, _03447_);
  nor _62009_ (_10529_, _10528_, _10526_);
  and _62010_ (_10530_, _05831_, _05221_);
  or _62011_ (_10531_, _10457_, _03514_);
  nor _62012_ (_10532_, _10531_, _10530_);
  nor _62013_ (_10533_, _10532_, _10529_);
  or _62014_ (_10534_, _10533_, _43004_);
  or _62015_ (_10535_, _43000_, \oc8051_golden_model_1.SBUF [7]);
  and _62016_ (_10536_, _10535_, _41806_);
  and _62017_ (_40580_, _10536_, _10534_);
  not _62018_ (_10537_, \oc8051_golden_model_1.SCON [7]);
  nor _62019_ (_10538_, _05275_, _10537_);
  not _62020_ (_10539_, _05275_);
  nor _62021_ (_10540_, _10539_, _05204_);
  nor _62022_ (_10541_, _10540_, _10538_);
  and _62023_ (_10542_, _10541_, _07390_);
  nor _62024_ (_10543_, _05922_, _10537_);
  and _62025_ (_10544_, _05952_, _05922_);
  nor _62026_ (_10545_, _10544_, _10543_);
  nor _62027_ (_10546_, _10545_, _03736_);
  and _62028_ (_10547_, _05275_, \oc8051_golden_model_1.ACC [7]);
  nor _62029_ (_10548_, _10547_, _10538_);
  nor _62030_ (_10549_, _10548_, _09029_);
  nor _62031_ (_10550_, _04409_, _10537_);
  or _62032_ (_10551_, _10550_, _10549_);
  and _62033_ (_10552_, _10551_, _04081_);
  and _62034_ (_10553_, _05964_, _05275_);
  nor _62035_ (_10554_, _10553_, _10538_);
  nor _62036_ (_10555_, _10554_, _04081_);
  or _62037_ (_10556_, _10555_, _10552_);
  and _62038_ (_10557_, _10556_, _04055_);
  and _62039_ (_10558_, _06095_, _05922_);
  nor _62040_ (_10559_, _10558_, _10543_);
  nor _62041_ (_10560_, _10559_, _04055_);
  or _62042_ (_10561_, _10560_, _03723_);
  or _62043_ (_10562_, _10561_, _10557_);
  nand _62044_ (_10563_, _10541_, _03723_);
  and _62045_ (_10564_, _10563_, _10562_);
  and _62046_ (_10565_, _10564_, _03737_);
  nor _62047_ (_10566_, _10548_, _03737_);
  or _62048_ (_10567_, _10566_, _10565_);
  and _62049_ (_10568_, _10567_, _03736_);
  nor _62050_ (_10569_, _10568_, _10546_);
  nor _62051_ (_10570_, _10569_, _03719_);
  nor _62052_ (_10571_, _10543_, _06138_);
  or _62053_ (_10572_, _10559_, _06840_);
  nor _62054_ (_10573_, _10572_, _10571_);
  nor _62055_ (_10574_, _10573_, _10570_);
  nor _62056_ (_10575_, _10574_, _03505_);
  not _62057_ (_10576_, _05922_);
  nor _62058_ (_10577_, _05938_, _10576_);
  nor _62059_ (_10578_, _10577_, _10543_);
  nor _62060_ (_10579_, _10578_, _03710_);
  nor _62061_ (_10580_, _10579_, _07390_);
  not _62062_ (_10581_, _10580_);
  nor _62063_ (_10582_, _10581_, _10575_);
  nor _62064_ (_10583_, _10582_, _10542_);
  nor _62065_ (_10584_, _10583_, _04481_);
  and _62066_ (_10585_, _06069_, _05275_);
  nor _62067_ (_10586_, _10538_, _07400_);
  not _62068_ (_10587_, _10586_);
  nor _62069_ (_10588_, _10587_, _10585_);
  nor _62070_ (_10589_, _10588_, _03222_);
  not _62071_ (_10590_, _10589_);
  nor _62072_ (_10591_, _10590_, _10584_);
  nor _62073_ (_10592_, _06363_, _10539_);
  nor _62074_ (_10593_, _10592_, _10538_);
  nor _62075_ (_10594_, _10593_, _03589_);
  or _62076_ (_10595_, _10594_, _08828_);
  or _62077_ (_10596_, _10595_, _10591_);
  and _62078_ (_10597_, _05884_, _05275_);
  or _62079_ (_10598_, _10538_, _07766_);
  or _62080_ (_10599_, _10598_, _10597_);
  and _62081_ (_10600_, _06171_, _05275_);
  nor _62082_ (_10601_, _10600_, _10538_);
  and _62083_ (_10602_, _10601_, _03601_);
  nor _62084_ (_10603_, _10602_, _03780_);
  and _62085_ (_10604_, _10603_, _10599_);
  and _62086_ (_10605_, _10604_, _10596_);
  and _62087_ (_10606_, _06378_, _05275_);
  nor _62088_ (_10607_, _10606_, _10538_);
  nor _62089_ (_10608_, _10607_, _07778_);
  nor _62090_ (_10609_, _10608_, _10605_);
  nor _62091_ (_10610_, _10609_, _03622_);
  nor _62092_ (_10611_, _10538_, _05310_);
  not _62093_ (_10612_, _10611_);
  nor _62094_ (_10613_, _10601_, _07777_);
  and _62095_ (_10614_, _10613_, _10612_);
  nor _62096_ (_10615_, _10614_, _10610_);
  nor _62097_ (_10616_, _10615_, _03790_);
  nor _62098_ (_10617_, _10548_, _06828_);
  and _62099_ (_10618_, _10617_, _10612_);
  nor _62100_ (_10619_, _10618_, _03624_);
  not _62101_ (_10620_, _10619_);
  nor _62102_ (_10621_, _10620_, _10616_);
  nor _62103_ (_10622_, _05882_, _10539_);
  or _62104_ (_10623_, _10538_, _07795_);
  nor _62105_ (_10624_, _10623_, _10622_);
  or _62106_ (_10625_, _10624_, _03785_);
  nor _62107_ (_10626_, _10625_, _10621_);
  nor _62108_ (_10627_, _06377_, _10539_);
  nor _62109_ (_10628_, _10627_, _10538_);
  nor _62110_ (_10629_, _10628_, _07793_);
  or _62111_ (_10630_, _10629_, _10626_);
  and _62112_ (_10631_, _10630_, _04246_);
  nor _62113_ (_10632_, _10554_, _04246_);
  or _62114_ (_10633_, _10632_, _10631_);
  and _62115_ (_10634_, _10633_, _03823_);
  nor _62116_ (_10635_, _10545_, _03823_);
  or _62117_ (_10636_, _10635_, _10634_);
  and _62118_ (_10637_, _10636_, _03514_);
  and _62119_ (_10638_, _05831_, _05275_);
  nor _62120_ (_10639_, _10638_, _10538_);
  nor _62121_ (_10640_, _10639_, _03514_);
  or _62122_ (_10641_, _10640_, _10637_);
  or _62123_ (_10642_, _10641_, _43004_);
  or _62124_ (_10643_, _43000_, \oc8051_golden_model_1.SCON [7]);
  and _62125_ (_10644_, _10643_, _41806_);
  and _62126_ (_40581_, _10644_, _10642_);
  and _62127_ (_10645_, _05010_, \oc8051_golden_model_1.SP [4]);
  and _62128_ (_10646_, _10645_, \oc8051_golden_model_1.SP [5]);
  and _62129_ (_10647_, _10646_, \oc8051_golden_model_1.SP [6]);
  nor _62130_ (_10648_, _10647_, \oc8051_golden_model_1.SP [7]);
  and _62131_ (_10649_, _10647_, \oc8051_golden_model_1.SP [7]);
  nor _62132_ (_10650_, _10649_, _10648_);
  nor _62133_ (_10651_, _10650_, _04540_);
  not _62134_ (_10652_, _03798_);
  not _62135_ (_10653_, \oc8051_golden_model_1.SP [7]);
  nor _62136_ (_10654_, _05300_, _10653_);
  and _62137_ (_10655_, _06378_, _05300_);
  nor _62138_ (_10656_, _10655_, _10654_);
  nor _62139_ (_10657_, _10656_, _07778_);
  not _62140_ (_10658_, _06837_);
  nor _62141_ (_10659_, _10650_, _04767_);
  nor _62142_ (_10660_, _04409_, _10653_);
  and _62143_ (_10661_, _05300_, \oc8051_golden_model_1.ACC [7]);
  nor _62144_ (_10662_, _10661_, _10654_);
  nor _62145_ (_10663_, _10662_, _09029_);
  or _62146_ (_10664_, _10663_, _10660_);
  and _62147_ (_10665_, _10664_, _04763_);
  and _62148_ (_10666_, _10650_, _03980_);
  nor _62149_ (_10667_, _10666_, _10665_);
  nor _62150_ (_10668_, _10667_, _03610_);
  and _62151_ (_10669_, _05964_, _05300_);
  nor _62152_ (_10670_, _10669_, _10654_);
  nor _62153_ (_10671_, _10670_, _04081_);
  or _62154_ (_10672_, _10671_, _10668_);
  and _62155_ (_10673_, _10672_, _03230_);
  and _62156_ (_10674_, _10650_, _04768_);
  or _62157_ (_10675_, _10674_, _10673_);
  and _62158_ (_10676_, _10675_, _03996_);
  not _62159_ (_10677_, \oc8051_golden_model_1.SP [6]);
  not _62160_ (_10678_, \oc8051_golden_model_1.SP [5]);
  not _62161_ (_10679_, \oc8051_golden_model_1.SP [4]);
  and _62162_ (_10680_, _05971_, _10679_);
  and _62163_ (_10681_, _10680_, _10678_);
  and _62164_ (_10682_, _10681_, _10677_);
  and _62165_ (_10683_, _10682_, _03498_);
  nor _62166_ (_10684_, _10683_, _10653_);
  and _62167_ (_10685_, _10683_, _10653_);
  nor _62168_ (_10686_, _10685_, _10684_);
  nor _62169_ (_10687_, _10686_, _03996_);
  or _62170_ (_10688_, _10687_, _10676_);
  and _62171_ (_10689_, _10688_, _03737_);
  nor _62172_ (_10691_, _10662_, _03737_);
  or _62173_ (_10692_, _10691_, _10689_);
  and _62174_ (_10693_, _10692_, _03510_);
  not _62175_ (_10694_, _04767_);
  and _62176_ (_10695_, _10647_, \oc8051_golden_model_1.SP [0]);
  nor _62177_ (_10696_, _10695_, _10653_);
  and _62178_ (_10697_, _10695_, _10653_);
  nor _62179_ (_10698_, _10697_, _10696_);
  nor _62180_ (_10699_, _10698_, _03510_);
  nor _62181_ (_10700_, _10699_, _10694_);
  not _62182_ (_10702_, _10700_);
  nor _62183_ (_10703_, _10702_, _10693_);
  nor _62184_ (_10704_, _10703_, _10659_);
  nor _62185_ (_10705_, _10704_, _10658_);
  not _62186_ (_10706_, _05300_);
  nor _62187_ (_10707_, _10706_, _05204_);
  nor _62188_ (_10708_, _10707_, _10654_);
  and _62189_ (_10709_, _10708_, _10658_);
  nor _62190_ (_10710_, _10709_, _06833_);
  not _62191_ (_10711_, _10710_);
  nor _62192_ (_10713_, _10711_, _10705_);
  nor _62193_ (_10714_, _10708_, _06834_);
  nor _62194_ (_10715_, _10714_, _04481_);
  not _62195_ (_10716_, _10715_);
  nor _62196_ (_10717_, _10716_, _10713_);
  and _62197_ (_10718_, _06069_, _05300_);
  nor _62198_ (_10719_, _10654_, _07400_);
  not _62199_ (_10720_, _10719_);
  nor _62200_ (_10721_, _10720_, _10718_);
  nor _62201_ (_10722_, _10721_, _10717_);
  nor _62202_ (_10724_, _10722_, _03222_);
  nor _62203_ (_10725_, _06363_, _10706_);
  or _62204_ (_10726_, _10654_, _03589_);
  nor _62205_ (_10727_, _10726_, _10725_);
  or _62206_ (_10728_, _10727_, _03601_);
  nor _62207_ (_10729_, _10728_, _10724_);
  and _62208_ (_10730_, _06171_, _05300_);
  nor _62209_ (_10731_, _10730_, _10654_);
  nor _62210_ (_10732_, _10731_, _05886_);
  or _62211_ (_10733_, _10732_, _03178_);
  or _62212_ (_10735_, _10733_, _10729_);
  not _62213_ (_10736_, _03178_);
  or _62214_ (_10737_, _10650_, _10736_);
  and _62215_ (_10738_, _10737_, _10735_);
  nor _62216_ (_10739_, _10738_, _03600_);
  and _62217_ (_10740_, _05884_, _05300_);
  or _62218_ (_10741_, _10654_, _07766_);
  nor _62219_ (_10742_, _10741_, _10740_);
  or _62220_ (_10743_, _10742_, _03780_);
  nor _62221_ (_10744_, _10743_, _10739_);
  nor _62222_ (_10746_, _10744_, _10657_);
  nor _62223_ (_10747_, _10746_, _03622_);
  nor _62224_ (_10748_, _10654_, _05310_);
  not _62225_ (_10749_, _10748_);
  nor _62226_ (_10750_, _10731_, _07777_);
  and _62227_ (_10751_, _10750_, _10749_);
  nor _62228_ (_10752_, _10751_, _10747_);
  nor _62229_ (_10753_, _03790_, _03192_);
  not _62230_ (_10754_, _10753_);
  nor _62231_ (_10755_, _10754_, _10752_);
  and _62232_ (_10757_, _10650_, _03192_);
  or _62233_ (_10758_, _10748_, _06828_);
  nor _62234_ (_10759_, _10758_, _10662_);
  nor _62235_ (_10760_, _10759_, _10757_);
  and _62236_ (_10761_, _10760_, _07795_);
  not _62237_ (_10762_, _10761_);
  nor _62238_ (_10763_, _10762_, _10755_);
  nor _62239_ (_10764_, _05882_, _10706_);
  nor _62240_ (_10765_, _10764_, _10654_);
  and _62241_ (_10766_, _10765_, _03624_);
  nor _62242_ (_10767_, _10766_, _10763_);
  and _62243_ (_10768_, _10767_, _07793_);
  nor _62244_ (_10769_, _06377_, _10706_);
  nor _62245_ (_10770_, _10769_, _10654_);
  nor _62246_ (_10771_, _10770_, _07793_);
  or _62247_ (_10772_, _10771_, _10768_);
  and _62248_ (_10773_, _10772_, _10652_);
  nor _62249_ (_10774_, _03798_, _03188_);
  nor _62250_ (_10775_, _10682_, \oc8051_golden_model_1.SP [7]);
  and _62251_ (_10776_, _10682_, \oc8051_golden_model_1.SP [7]);
  nor _62252_ (_10777_, _10776_, _10775_);
  nor _62253_ (_10778_, _10777_, _03188_);
  nor _62254_ (_10779_, _10778_, _10774_);
  nor _62255_ (_10780_, _10779_, _10773_);
  nor _62256_ (_10781_, _10650_, _06399_);
  nor _62257_ (_10782_, _10781_, _10780_);
  and _62258_ (_10783_, _10782_, _03516_);
  and _62259_ (_10784_, _10777_, _03515_);
  or _62260_ (_10785_, _10784_, _10783_);
  and _62261_ (_10786_, _10785_, _04246_);
  nor _62262_ (_10787_, _10670_, _04246_);
  nor _62263_ (_10788_, _10787_, _05103_);
  not _62264_ (_10789_, _10788_);
  nor _62265_ (_10790_, _10789_, _10786_);
  nor _62266_ (_10791_, _10790_, _10651_);
  and _62267_ (_10792_, _10791_, _03514_);
  and _62268_ (_10793_, _05831_, _05300_);
  nor _62269_ (_10794_, _10793_, _10654_);
  nor _62270_ (_10795_, _10794_, _03514_);
  or _62271_ (_10796_, _10795_, _10792_);
  or _62272_ (_10797_, _10796_, _43004_);
  or _62273_ (_10798_, _43000_, \oc8051_golden_model_1.SP [7]);
  and _62274_ (_10799_, _10798_, _41806_);
  and _62275_ (_40583_, _10799_, _10797_);
  not _62276_ (_10800_, \oc8051_golden_model_1.TCON [7]);
  nor _62277_ (_10801_, _05258_, _10800_);
  not _62278_ (_10802_, _05258_);
  nor _62279_ (_10803_, _10802_, _05204_);
  nor _62280_ (_10804_, _10803_, _10801_);
  and _62281_ (_10805_, _10804_, _07390_);
  nor _62282_ (_10806_, _05927_, _10800_);
  and _62283_ (_10807_, _05952_, _05927_);
  nor _62284_ (_10808_, _10807_, _10806_);
  nor _62285_ (_10809_, _10808_, _03736_);
  and _62286_ (_10810_, _05258_, \oc8051_golden_model_1.ACC [7]);
  nor _62287_ (_10811_, _10810_, _10801_);
  nor _62288_ (_10812_, _10811_, _09029_);
  nor _62289_ (_10813_, _04409_, _10800_);
  or _62290_ (_10814_, _10813_, _10812_);
  and _62291_ (_10815_, _10814_, _04081_);
  and _62292_ (_10816_, _05964_, _05258_);
  nor _62293_ (_10817_, _10816_, _10801_);
  nor _62294_ (_10818_, _10817_, _04081_);
  or _62295_ (_10819_, _10818_, _10815_);
  and _62296_ (_10820_, _10819_, _04055_);
  and _62297_ (_10821_, _06095_, _05927_);
  nor _62298_ (_10822_, _10821_, _10806_);
  nor _62299_ (_10823_, _10822_, _04055_);
  or _62300_ (_10824_, _10823_, _03723_);
  or _62301_ (_10825_, _10824_, _10820_);
  nand _62302_ (_10826_, _10804_, _03723_);
  and _62303_ (_10827_, _10826_, _10825_);
  and _62304_ (_10828_, _10827_, _03737_);
  nor _62305_ (_10829_, _10811_, _03737_);
  or _62306_ (_10830_, _10829_, _10828_);
  and _62307_ (_10831_, _10830_, _03736_);
  nor _62308_ (_10832_, _10831_, _10809_);
  nor _62309_ (_10833_, _10832_, _03719_);
  and _62310_ (_10834_, _06139_, _05927_);
  nor _62311_ (_10835_, _10834_, _10806_);
  nor _62312_ (_10836_, _10835_, _06840_);
  nor _62313_ (_10837_, _10836_, _10833_);
  nor _62314_ (_10838_, _10837_, _03505_);
  not _62315_ (_10839_, _05927_);
  nor _62316_ (_10840_, _05938_, _10839_);
  nor _62317_ (_10841_, _10840_, _10806_);
  nor _62318_ (_10842_, _10841_, _03710_);
  nor _62319_ (_10843_, _10842_, _07390_);
  not _62320_ (_10844_, _10843_);
  nor _62321_ (_10845_, _10844_, _10838_);
  nor _62322_ (_10846_, _10845_, _10805_);
  nor _62323_ (_10847_, _10846_, _04481_);
  and _62324_ (_10848_, _06069_, _05258_);
  nor _62325_ (_10849_, _10801_, _07400_);
  not _62326_ (_10850_, _10849_);
  nor _62327_ (_10851_, _10850_, _10848_);
  nor _62328_ (_10852_, _10851_, _03222_);
  not _62329_ (_10853_, _10852_);
  nor _62330_ (_10854_, _10853_, _10847_);
  nor _62331_ (_10855_, _06363_, _10802_);
  nor _62332_ (_10856_, _10855_, _10801_);
  nor _62333_ (_10857_, _10856_, _03589_);
  or _62334_ (_10858_, _10857_, _08828_);
  or _62335_ (_10859_, _10858_, _10854_);
  and _62336_ (_10860_, _05884_, _05258_);
  or _62337_ (_10861_, _10801_, _07766_);
  or _62338_ (_10862_, _10861_, _10860_);
  and _62339_ (_10863_, _06171_, _05258_);
  nor _62340_ (_10864_, _10863_, _10801_);
  and _62341_ (_10865_, _10864_, _03601_);
  nor _62342_ (_10866_, _10865_, _03780_);
  and _62343_ (_10867_, _10866_, _10862_);
  and _62344_ (_10868_, _10867_, _10859_);
  and _62345_ (_10869_, _06378_, _05258_);
  nor _62346_ (_10870_, _10869_, _10801_);
  nor _62347_ (_10871_, _10870_, _07778_);
  nor _62348_ (_10872_, _10871_, _10868_);
  nor _62349_ (_10873_, _10872_, _03622_);
  nor _62350_ (_10874_, _10801_, _05310_);
  not _62351_ (_10875_, _10874_);
  nor _62352_ (_10876_, _10864_, _07777_);
  and _62353_ (_10877_, _10876_, _10875_);
  nor _62354_ (_10878_, _10877_, _10873_);
  nor _62355_ (_10879_, _10878_, _03790_);
  nor _62356_ (_10880_, _10811_, _06828_);
  and _62357_ (_10881_, _10880_, _10875_);
  or _62358_ (_10882_, _10881_, _10879_);
  and _62359_ (_10883_, _10882_, _07795_);
  nor _62360_ (_10884_, _05882_, _10802_);
  nor _62361_ (_10885_, _10884_, _10801_);
  nor _62362_ (_10886_, _10885_, _07795_);
  or _62363_ (_10887_, _10886_, _10883_);
  and _62364_ (_10888_, _10887_, _07793_);
  nor _62365_ (_10889_, _06377_, _10802_);
  nor _62366_ (_10890_, _10889_, _10801_);
  nor _62367_ (_10891_, _10890_, _07793_);
  or _62368_ (_10892_, _10891_, _10888_);
  and _62369_ (_10893_, _10892_, _04246_);
  nor _62370_ (_10894_, _10817_, _04246_);
  or _62371_ (_10895_, _10894_, _10893_);
  and _62372_ (_10896_, _10895_, _03823_);
  nor _62373_ (_10897_, _10808_, _03823_);
  or _62374_ (_10898_, _10897_, _10896_);
  and _62375_ (_10899_, _10898_, _03514_);
  and _62376_ (_10900_, _05831_, _05258_);
  nor _62377_ (_10901_, _10900_, _10801_);
  nor _62378_ (_10902_, _10901_, _03514_);
  or _62379_ (_10903_, _10902_, _10899_);
  or _62380_ (_10904_, _10903_, _43004_);
  or _62381_ (_10905_, _43000_, \oc8051_golden_model_1.TCON [7]);
  and _62382_ (_10906_, _10905_, _41806_);
  and _62383_ (_40584_, _10906_, _10904_);
  not _62384_ (_10907_, \oc8051_golden_model_1.TH0 [7]);
  nor _62385_ (_10908_, _05263_, _10907_);
  not _62386_ (_10909_, _05263_);
  nor _62387_ (_10910_, _06377_, _10909_);
  nor _62388_ (_10911_, _10910_, _10908_);
  nor _62389_ (_10912_, _10911_, _07793_);
  and _62390_ (_10913_, _06171_, _05263_);
  nor _62391_ (_10914_, _10913_, _10908_);
  and _62392_ (_10915_, _10914_, _03601_);
  nor _62393_ (_10916_, _10909_, _05204_);
  nor _62394_ (_10917_, _10916_, _10908_);
  and _62395_ (_10918_, _10917_, _07390_);
  and _62396_ (_10919_, _05263_, \oc8051_golden_model_1.ACC [7]);
  nor _62397_ (_10920_, _10919_, _10908_);
  nor _62398_ (_10921_, _10920_, _03737_);
  nor _62399_ (_10922_, _10920_, _09029_);
  nor _62400_ (_10923_, _04409_, _10907_);
  or _62401_ (_10924_, _10923_, _10922_);
  and _62402_ (_10925_, _10924_, _04081_);
  and _62403_ (_10926_, _05964_, _05263_);
  nor _62404_ (_10927_, _10926_, _10908_);
  nor _62405_ (_10928_, _10927_, _04081_);
  or _62406_ (_10929_, _10928_, _10925_);
  and _62407_ (_10930_, _10929_, _03996_);
  nor _62408_ (_10931_, _10917_, _03996_);
  nor _62409_ (_10932_, _10931_, _10930_);
  nor _62410_ (_10933_, _10932_, _03729_);
  or _62411_ (_10934_, _10933_, _07390_);
  nor _62412_ (_10935_, _10934_, _10921_);
  nor _62413_ (_10936_, _10935_, _10918_);
  nor _62414_ (_10937_, _10936_, _04481_);
  and _62415_ (_10938_, _06069_, _05263_);
  nor _62416_ (_10939_, _10908_, _07400_);
  not _62417_ (_10940_, _10939_);
  nor _62418_ (_10941_, _10940_, _10938_);
  or _62419_ (_10942_, _10941_, _03222_);
  nor _62420_ (_10943_, _10942_, _10937_);
  nor _62421_ (_10944_, _06363_, _10909_);
  nor _62422_ (_10945_, _10944_, _10908_);
  nor _62423_ (_10946_, _10945_, _03589_);
  or _62424_ (_10947_, _10946_, _03601_);
  nor _62425_ (_10948_, _10947_, _10943_);
  nor _62426_ (_10949_, _10948_, _10915_);
  or _62427_ (_10950_, _10949_, _03600_);
  and _62428_ (_10951_, _05884_, _05263_);
  or _62429_ (_10952_, _10951_, _10908_);
  or _62430_ (_10953_, _10952_, _07766_);
  and _62431_ (_10954_, _10953_, _07778_);
  and _62432_ (_10955_, _10954_, _10950_);
  and _62433_ (_10956_, _06378_, _05263_);
  nor _62434_ (_10957_, _10956_, _10908_);
  nor _62435_ (_10958_, _10957_, _07778_);
  nor _62436_ (_10959_, _10958_, _10955_);
  nor _62437_ (_10960_, _10959_, _03622_);
  nor _62438_ (_10961_, _10908_, _05310_);
  not _62439_ (_10962_, _10961_);
  nor _62440_ (_10963_, _10914_, _07777_);
  and _62441_ (_10964_, _10963_, _10962_);
  nor _62442_ (_10965_, _10964_, _10960_);
  nor _62443_ (_10966_, _10965_, _03790_);
  nor _62444_ (_10967_, _10920_, _06828_);
  and _62445_ (_10968_, _10967_, _10962_);
  nor _62446_ (_10969_, _10968_, _03624_);
  not _62447_ (_10970_, _10969_);
  nor _62448_ (_10971_, _10970_, _10966_);
  nor _62449_ (_10972_, _05882_, _10909_);
  or _62450_ (_10973_, _10908_, _07795_);
  nor _62451_ (_10974_, _10973_, _10972_);
  or _62452_ (_10975_, _10974_, _03785_);
  nor _62453_ (_10976_, _10975_, _10971_);
  nor _62454_ (_10977_, _10976_, _10912_);
  nor _62455_ (_10978_, _10977_, _03815_);
  nor _62456_ (_10979_, _10927_, _04246_);
  or _62457_ (_10980_, _10979_, _03447_);
  nor _62458_ (_10981_, _10980_, _10978_);
  and _62459_ (_10982_, _05831_, _05263_);
  or _62460_ (_10983_, _10908_, _03514_);
  nor _62461_ (_10984_, _10983_, _10982_);
  nor _62462_ (_10985_, _10984_, _10981_);
  or _62463_ (_10986_, _10985_, _43004_);
  or _62464_ (_10987_, _43000_, \oc8051_golden_model_1.TH0 [7]);
  and _62465_ (_10988_, _10987_, _41806_);
  and _62466_ (_40585_, _10988_, _10986_);
  not _62467_ (_10989_, \oc8051_golden_model_1.TH1 [7]);
  nor _62468_ (_10990_, _05278_, _10989_);
  not _62469_ (_10991_, _05278_);
  nor _62470_ (_10992_, _06377_, _10991_);
  nor _62471_ (_10993_, _10992_, _10990_);
  nor _62472_ (_10994_, _10993_, _07793_);
  and _62473_ (_10995_, _06171_, _05278_);
  nor _62474_ (_10996_, _10995_, _10990_);
  and _62475_ (_10997_, _10996_, _03601_);
  and _62476_ (_10998_, _05278_, \oc8051_golden_model_1.ACC [7]);
  nor _62477_ (_10999_, _10998_, _10990_);
  nor _62478_ (_11000_, _10999_, _03737_);
  nor _62479_ (_11001_, _10999_, _09029_);
  nor _62480_ (_11002_, _04409_, _10989_);
  or _62481_ (_11003_, _11002_, _11001_);
  and _62482_ (_11004_, _11003_, _04081_);
  and _62483_ (_11005_, _05964_, _05278_);
  nor _62484_ (_11006_, _11005_, _10990_);
  nor _62485_ (_11007_, _11006_, _04081_);
  or _62486_ (_11008_, _11007_, _11004_);
  and _62487_ (_11009_, _11008_, _03996_);
  nor _62488_ (_11010_, _10991_, _05204_);
  nor _62489_ (_11011_, _11010_, _10990_);
  nor _62490_ (_11012_, _11011_, _03996_);
  nor _62491_ (_11013_, _11012_, _11009_);
  nor _62492_ (_11014_, _11013_, _03729_);
  or _62493_ (_11015_, _11014_, _07390_);
  nor _62494_ (_11016_, _11015_, _11000_);
  and _62495_ (_11017_, _11011_, _07390_);
  nor _62496_ (_11018_, _11017_, _11016_);
  nor _62497_ (_11019_, _11018_, _04481_);
  and _62498_ (_11020_, _06069_, _05278_);
  nor _62499_ (_11021_, _10990_, _07400_);
  not _62500_ (_11022_, _11021_);
  nor _62501_ (_11023_, _11022_, _11020_);
  or _62502_ (_11024_, _11023_, _03222_);
  nor _62503_ (_11025_, _11024_, _11019_);
  nor _62504_ (_11026_, _06363_, _10991_);
  nor _62505_ (_11027_, _11026_, _10990_);
  nor _62506_ (_11028_, _11027_, _03589_);
  or _62507_ (_11029_, _11028_, _03601_);
  nor _62508_ (_11030_, _11029_, _11025_);
  nor _62509_ (_11031_, _11030_, _10997_);
  or _62510_ (_11032_, _11031_, _03600_);
  and _62511_ (_11033_, _05884_, _05278_);
  or _62512_ (_11034_, _11033_, _10990_);
  or _62513_ (_11035_, _11034_, _07766_);
  and _62514_ (_11036_, _11035_, _07778_);
  and _62515_ (_11037_, _11036_, _11032_);
  and _62516_ (_11038_, _06378_, _05278_);
  nor _62517_ (_11039_, _11038_, _10990_);
  nor _62518_ (_11040_, _11039_, _07778_);
  nor _62519_ (_11041_, _11040_, _11037_);
  nor _62520_ (_11042_, _11041_, _03622_);
  nor _62521_ (_11043_, _10990_, _05310_);
  not _62522_ (_11044_, _11043_);
  nor _62523_ (_11045_, _10996_, _07777_);
  and _62524_ (_11046_, _11045_, _11044_);
  nor _62525_ (_11047_, _11046_, _11042_);
  nor _62526_ (_11048_, _11047_, _03790_);
  nor _62527_ (_11049_, _10999_, _06828_);
  and _62528_ (_11050_, _11049_, _11044_);
  or _62529_ (_11051_, _11050_, _11048_);
  and _62530_ (_11052_, _11051_, _07795_);
  nor _62531_ (_11053_, _05882_, _10991_);
  nor _62532_ (_11054_, _11053_, _10990_);
  nor _62533_ (_11055_, _11054_, _07795_);
  or _62534_ (_11056_, _11055_, _11052_);
  and _62535_ (_11057_, _11056_, _07793_);
  nor _62536_ (_11058_, _11057_, _10994_);
  nor _62537_ (_11059_, _11058_, _03815_);
  nor _62538_ (_11060_, _11006_, _04246_);
  or _62539_ (_11061_, _11060_, _03447_);
  nor _62540_ (_11062_, _11061_, _11059_);
  and _62541_ (_11063_, _05831_, _05278_);
  or _62542_ (_11064_, _10990_, _03514_);
  nor _62543_ (_11065_, _11064_, _11063_);
  nor _62544_ (_11066_, _11065_, _11062_);
  or _62545_ (_11067_, _11066_, _43004_);
  or _62546_ (_11068_, _43000_, \oc8051_golden_model_1.TH1 [7]);
  and _62547_ (_11069_, _11068_, _41806_);
  and _62548_ (_40586_, _11069_, _11067_);
  not _62549_ (_11070_, \oc8051_golden_model_1.TL0 [7]);
  nor _62550_ (_11071_, _05284_, _11070_);
  not _62551_ (_11072_, _05284_);
  nor _62552_ (_11073_, _06377_, _11072_);
  nor _62553_ (_11074_, _11073_, _11071_);
  nor _62554_ (_11075_, _11074_, _07793_);
  and _62555_ (_11076_, _06171_, _05284_);
  nor _62556_ (_11077_, _11076_, _11071_);
  and _62557_ (_11078_, _11077_, _03601_);
  and _62558_ (_11079_, _05284_, \oc8051_golden_model_1.ACC [7]);
  nor _62559_ (_11080_, _11079_, _11071_);
  nor _62560_ (_11081_, _11080_, _03737_);
  nor _62561_ (_11082_, _11080_, _09029_);
  nor _62562_ (_11083_, _04409_, _11070_);
  or _62563_ (_11084_, _11083_, _11082_);
  and _62564_ (_11085_, _11084_, _04081_);
  and _62565_ (_11086_, _05964_, _05284_);
  nor _62566_ (_11087_, _11086_, _11071_);
  nor _62567_ (_11088_, _11087_, _04081_);
  or _62568_ (_11089_, _11088_, _11085_);
  and _62569_ (_11090_, _11089_, _03996_);
  nor _62570_ (_11091_, _11072_, _05204_);
  nor _62571_ (_11092_, _11091_, _11071_);
  nor _62572_ (_11093_, _11092_, _03996_);
  nor _62573_ (_11094_, _11093_, _11090_);
  nor _62574_ (_11095_, _11094_, _03729_);
  or _62575_ (_11096_, _11095_, _07390_);
  nor _62576_ (_11097_, _11096_, _11081_);
  and _62577_ (_11098_, _11092_, _07390_);
  nor _62578_ (_11099_, _11098_, _11097_);
  nor _62579_ (_11100_, _11099_, _04481_);
  and _62580_ (_11101_, _06069_, _05284_);
  nor _62581_ (_11102_, _11071_, _07400_);
  not _62582_ (_11103_, _11102_);
  nor _62583_ (_11104_, _11103_, _11101_);
  or _62584_ (_11105_, _11104_, _03222_);
  nor _62585_ (_11106_, _11105_, _11100_);
  nor _62586_ (_11107_, _06363_, _11072_);
  nor _62587_ (_11108_, _11107_, _11071_);
  nor _62588_ (_11109_, _11108_, _03589_);
  or _62589_ (_11110_, _11109_, _03601_);
  nor _62590_ (_11111_, _11110_, _11106_);
  nor _62591_ (_11112_, _11111_, _11078_);
  or _62592_ (_11113_, _11112_, _03600_);
  and _62593_ (_11114_, _05884_, _05284_);
  or _62594_ (_11115_, _11114_, _11071_);
  or _62595_ (_11116_, _11115_, _07766_);
  and _62596_ (_11117_, _11116_, _07778_);
  and _62597_ (_11118_, _11117_, _11113_);
  and _62598_ (_11119_, _06378_, _05284_);
  nor _62599_ (_11120_, _11119_, _11071_);
  nor _62600_ (_11121_, _11120_, _07778_);
  nor _62601_ (_11122_, _11121_, _11118_);
  nor _62602_ (_11123_, _11122_, _03622_);
  nor _62603_ (_11124_, _11071_, _05310_);
  not _62604_ (_11125_, _11124_);
  nor _62605_ (_11126_, _11077_, _07777_);
  and _62606_ (_11127_, _11126_, _11125_);
  nor _62607_ (_11128_, _11127_, _11123_);
  nor _62608_ (_11129_, _11128_, _03790_);
  nor _62609_ (_11130_, _11080_, _06828_);
  and _62610_ (_11131_, _11130_, _11125_);
  nor _62611_ (_11132_, _11131_, _03624_);
  not _62612_ (_11133_, _11132_);
  nor _62613_ (_11134_, _11133_, _11129_);
  nor _62614_ (_11135_, _05882_, _11072_);
  or _62615_ (_11136_, _11071_, _07795_);
  nor _62616_ (_11137_, _11136_, _11135_);
  or _62617_ (_11138_, _11137_, _03785_);
  nor _62618_ (_11139_, _11138_, _11134_);
  nor _62619_ (_11140_, _11139_, _11075_);
  nor _62620_ (_11141_, _11140_, _03815_);
  nor _62621_ (_11142_, _11087_, _04246_);
  or _62622_ (_11143_, _11142_, _03447_);
  nor _62623_ (_11144_, _11143_, _11141_);
  and _62624_ (_11145_, _05831_, _05284_);
  nor _62625_ (_11146_, _11145_, _11071_);
  and _62626_ (_11147_, _11146_, _03447_);
  nor _62627_ (_11148_, _11147_, _11144_);
  or _62628_ (_11149_, _11148_, _43004_);
  or _62629_ (_11150_, _43000_, \oc8051_golden_model_1.TL0 [7]);
  and _62630_ (_11151_, _11150_, _41806_);
  and _62631_ (_40587_, _11151_, _11149_);
  not _62632_ (_11152_, \oc8051_golden_model_1.TL1 [7]);
  nor _62633_ (_11153_, _05271_, _11152_);
  not _62634_ (_11154_, _05271_);
  nor _62635_ (_11155_, _06377_, _11154_);
  nor _62636_ (_11156_, _11155_, _11153_);
  nor _62637_ (_11157_, _11156_, _07793_);
  and _62638_ (_11158_, _06171_, _05271_);
  nor _62639_ (_11159_, _11158_, _11153_);
  and _62640_ (_11160_, _11159_, _03601_);
  and _62641_ (_11161_, _05271_, \oc8051_golden_model_1.ACC [7]);
  nor _62642_ (_11162_, _11161_, _11153_);
  nor _62643_ (_11163_, _11162_, _03737_);
  nor _62644_ (_11164_, _11162_, _09029_);
  nor _62645_ (_11165_, _04409_, _11152_);
  or _62646_ (_11166_, _11165_, _11164_);
  and _62647_ (_11167_, _11166_, _04081_);
  and _62648_ (_11168_, _05964_, _05271_);
  nor _62649_ (_11169_, _11168_, _11153_);
  nor _62650_ (_11170_, _11169_, _04081_);
  or _62651_ (_11171_, _11170_, _11167_);
  and _62652_ (_11172_, _11171_, _03996_);
  nor _62653_ (_11173_, _11154_, _05204_);
  nor _62654_ (_11174_, _11173_, _11153_);
  nor _62655_ (_11175_, _11174_, _03996_);
  nor _62656_ (_11176_, _11175_, _11172_);
  nor _62657_ (_11177_, _11176_, _03729_);
  or _62658_ (_11178_, _11177_, _07390_);
  nor _62659_ (_11179_, _11178_, _11163_);
  and _62660_ (_11180_, _11174_, _07390_);
  nor _62661_ (_11181_, _11180_, _11179_);
  nor _62662_ (_11182_, _11181_, _04481_);
  and _62663_ (_11183_, _06069_, _05271_);
  nor _62664_ (_11184_, _11153_, _07400_);
  not _62665_ (_11185_, _11184_);
  nor _62666_ (_11186_, _11185_, _11183_);
  or _62667_ (_11187_, _11186_, _03222_);
  nor _62668_ (_11188_, _11187_, _11182_);
  nor _62669_ (_11189_, _06363_, _11154_);
  nor _62670_ (_11190_, _11189_, _11153_);
  nor _62671_ (_11191_, _11190_, _03589_);
  or _62672_ (_11192_, _11191_, _03601_);
  nor _62673_ (_11193_, _11192_, _11188_);
  nor _62674_ (_11194_, _11193_, _11160_);
  or _62675_ (_11195_, _11194_, _03600_);
  and _62676_ (_11196_, _05884_, _05271_);
  or _62677_ (_11197_, _11196_, _11153_);
  or _62678_ (_11198_, _11197_, _07766_);
  and _62679_ (_11199_, _11198_, _07778_);
  and _62680_ (_11200_, _11199_, _11195_);
  and _62681_ (_11201_, _06378_, _05271_);
  nor _62682_ (_11202_, _11201_, _11153_);
  nor _62683_ (_11203_, _11202_, _07778_);
  nor _62684_ (_11204_, _11203_, _11200_);
  nor _62685_ (_11205_, _11204_, _03622_);
  nor _62686_ (_11206_, _11153_, _05310_);
  not _62687_ (_11207_, _11206_);
  nor _62688_ (_11208_, _11159_, _07777_);
  and _62689_ (_11209_, _11208_, _11207_);
  nor _62690_ (_11210_, _11209_, _11205_);
  nor _62691_ (_11211_, _11210_, _03790_);
  nor _62692_ (_11212_, _11162_, _06828_);
  and _62693_ (_11213_, _11212_, _11207_);
  nor _62694_ (_11214_, _11213_, _03624_);
  not _62695_ (_11215_, _11214_);
  nor _62696_ (_11216_, _11215_, _11211_);
  nor _62697_ (_11217_, _05882_, _11154_);
  or _62698_ (_11218_, _11153_, _07795_);
  nor _62699_ (_11219_, _11218_, _11217_);
  or _62700_ (_11220_, _11219_, _03785_);
  nor _62701_ (_11221_, _11220_, _11216_);
  nor _62702_ (_11222_, _11221_, _11157_);
  nor _62703_ (_11223_, _11222_, _03815_);
  nor _62704_ (_11224_, _11169_, _04246_);
  or _62705_ (_11225_, _11224_, _03447_);
  nor _62706_ (_11226_, _11225_, _11223_);
  and _62707_ (_11227_, _05831_, _05271_);
  or _62708_ (_11228_, _11153_, _03514_);
  nor _62709_ (_11229_, _11228_, _11227_);
  nor _62710_ (_11230_, _11229_, _11226_);
  or _62711_ (_11231_, _11230_, _43004_);
  or _62712_ (_11232_, _43000_, \oc8051_golden_model_1.TL1 [7]);
  and _62713_ (_11233_, _11232_, _41806_);
  and _62714_ (_40589_, _11233_, _11231_);
  not _62715_ (_11234_, \oc8051_golden_model_1.TMOD [7]);
  nor _62716_ (_11235_, _05286_, _11234_);
  not _62717_ (_11236_, _05286_);
  nor _62718_ (_11237_, _06377_, _11236_);
  nor _62719_ (_11238_, _11237_, _11235_);
  nor _62720_ (_11239_, _11238_, _07793_);
  and _62721_ (_11240_, _06171_, _05286_);
  nor _62722_ (_11241_, _11240_, _11235_);
  and _62723_ (_11242_, _11241_, _03601_);
  and _62724_ (_11243_, _05286_, \oc8051_golden_model_1.ACC [7]);
  nor _62725_ (_11244_, _11243_, _11235_);
  nor _62726_ (_11245_, _11244_, _03737_);
  nor _62727_ (_11246_, _11244_, _09029_);
  nor _62728_ (_11247_, _04409_, _11234_);
  or _62729_ (_11248_, _11247_, _11246_);
  and _62730_ (_11249_, _11248_, _04081_);
  and _62731_ (_11250_, _05964_, _05286_);
  nor _62732_ (_11251_, _11250_, _11235_);
  nor _62733_ (_11252_, _11251_, _04081_);
  or _62734_ (_11253_, _11252_, _11249_);
  and _62735_ (_11254_, _11253_, _03996_);
  nor _62736_ (_11255_, _11236_, _05204_);
  nor _62737_ (_11256_, _11255_, _11235_);
  nor _62738_ (_11257_, _11256_, _03996_);
  nor _62739_ (_11258_, _11257_, _11254_);
  nor _62740_ (_11259_, _11258_, _03729_);
  or _62741_ (_11260_, _11259_, _07390_);
  nor _62742_ (_11261_, _11260_, _11245_);
  and _62743_ (_11262_, _11256_, _07390_);
  nor _62744_ (_11263_, _11262_, _11261_);
  nor _62745_ (_11264_, _11263_, _04481_);
  and _62746_ (_11265_, _06069_, _05286_);
  nor _62747_ (_11266_, _11235_, _07400_);
  not _62748_ (_11267_, _11266_);
  nor _62749_ (_11268_, _11267_, _11265_);
  or _62750_ (_11269_, _11268_, _03222_);
  nor _62751_ (_11270_, _11269_, _11264_);
  nor _62752_ (_11271_, _06363_, _11236_);
  nor _62753_ (_11272_, _11271_, _11235_);
  nor _62754_ (_11273_, _11272_, _03589_);
  or _62755_ (_11274_, _11273_, _03601_);
  nor _62756_ (_11275_, _11274_, _11270_);
  nor _62757_ (_11276_, _11275_, _11242_);
  or _62758_ (_11277_, _11276_, _03600_);
  and _62759_ (_11278_, _05884_, _05286_);
  or _62760_ (_11279_, _11278_, _11235_);
  or _62761_ (_11280_, _11279_, _07766_);
  and _62762_ (_11281_, _11280_, _07778_);
  and _62763_ (_11282_, _11281_, _11277_);
  and _62764_ (_11283_, _06378_, _05286_);
  nor _62765_ (_11284_, _11283_, _11235_);
  nor _62766_ (_11285_, _11284_, _07778_);
  nor _62767_ (_11286_, _11285_, _11282_);
  nor _62768_ (_11287_, _11286_, _03622_);
  nor _62769_ (_11288_, _11235_, _05310_);
  not _62770_ (_11289_, _11288_);
  nor _62771_ (_11290_, _11241_, _07777_);
  and _62772_ (_11291_, _11290_, _11289_);
  nor _62773_ (_11292_, _11291_, _11287_);
  nor _62774_ (_11293_, _11292_, _03790_);
  nor _62775_ (_11294_, _11244_, _06828_);
  and _62776_ (_11295_, _11294_, _11289_);
  or _62777_ (_11296_, _11295_, _11293_);
  and _62778_ (_11297_, _11296_, _07795_);
  nor _62779_ (_11298_, _05882_, _11236_);
  nor _62780_ (_11299_, _11298_, _11235_);
  nor _62781_ (_11300_, _11299_, _07795_);
  or _62782_ (_11301_, _11300_, _11297_);
  and _62783_ (_11302_, _11301_, _07793_);
  nor _62784_ (_11303_, _11302_, _11239_);
  nor _62785_ (_11304_, _11303_, _03815_);
  nor _62786_ (_11305_, _11251_, _04246_);
  or _62787_ (_11306_, _11305_, _03447_);
  nor _62788_ (_11307_, _11306_, _11304_);
  and _62789_ (_11308_, _05831_, _05286_);
  or _62790_ (_11309_, _11235_, _03514_);
  nor _62791_ (_11310_, _11309_, _11308_);
  nor _62792_ (_11311_, _11310_, _11307_);
  or _62793_ (_11312_, _11311_, _43004_);
  or _62794_ (_11313_, _43000_, \oc8051_golden_model_1.TMOD [7]);
  and _62795_ (_11314_, _11313_, _41806_);
  and _62796_ (_40590_, _11314_, _11312_);
  not _62797_ (_11315_, _02892_);
  and _62798_ (_11316_, _06078_, _11315_);
  and _62799_ (_11317_, _11316_, \oc8051_golden_model_1.PC [7]);
  and _62800_ (_11318_, _11317_, \oc8051_golden_model_1.PC [8]);
  and _62801_ (_11319_, _11318_, \oc8051_golden_model_1.PC [9]);
  and _62802_ (_11320_, _11319_, \oc8051_golden_model_1.PC [10]);
  and _62803_ (_11321_, _11320_, \oc8051_golden_model_1.PC [11]);
  and _62804_ (_11322_, _11321_, \oc8051_golden_model_1.PC [12]);
  and _62805_ (_11323_, _11322_, \oc8051_golden_model_1.PC [13]);
  and _62806_ (_11324_, _11323_, \oc8051_golden_model_1.PC [14]);
  or _62807_ (_11325_, _11324_, \oc8051_golden_model_1.PC [15]);
  nand _62808_ (_11326_, _11324_, \oc8051_golden_model_1.PC [15]);
  and _62809_ (_11327_, _11326_, _11325_);
  nor _62810_ (_11328_, _08620_, _08618_);
  or _62811_ (_11329_, _11328_, _11327_);
  and _62812_ (_11330_, _08477_, _07898_);
  or _62813_ (_11331_, _11330_, _11327_);
  nor _62814_ (_11332_, _08441_, _04306_);
  and _62815_ (_11333_, _03494_, _03200_);
  nor _62816_ (_11334_, _08450_, _11333_);
  and _62817_ (_11335_, _11334_, _11332_);
  or _62818_ (_11336_, _11335_, _11327_);
  and _62819_ (_11337_, _03191_, _03452_);
  not _62820_ (_11338_, _11337_);
  or _62821_ (_11339_, _10753_, _06813_);
  and _62822_ (_11340_, _11339_, _11338_);
  nor _62823_ (_11341_, _07904_, _03778_);
  not _62824_ (_11342_, _11341_);
  nand _62825_ (_11343_, _03181_, _02962_);
  not _62826_ (_11344_, _11343_);
  nor _62827_ (_11345_, _11344_, _08392_);
  or _62828_ (_11346_, _11345_, _11327_);
  and _62829_ (_11347_, _03599_, _03176_);
  not _62830_ (_11348_, _11347_);
  and _62831_ (_11349_, _06821_, _03222_);
  and _62832_ (_11350_, _08059_, _10201_);
  or _62833_ (_11351_, _11350_, _11327_);
  and _62834_ (_11352_, _03751_, _03221_);
  not _62835_ (_11353_, _11352_);
  nor _62836_ (_11354_, _08847_, _06869_);
  and _62837_ (_11355_, _11354_, _11353_);
  not _62838_ (_11356_, _11355_);
  and _62839_ (_11357_, _11356_, _11327_);
  not _62840_ (_11358_, _10025_);
  and _62841_ (_11359_, _06813_, _03729_);
  and _62842_ (_11360_, _03730_, _03230_);
  or _62843_ (_11361_, _11360_, _06813_);
  nor _62844_ (_11362_, _09895_, _08089_);
  and _62845_ (_11363_, _05666_, _05617_);
  and _62846_ (_11364_, _05958_, _11363_);
  and _62847_ (_11365_, _05411_, _05309_);
  and _62848_ (_11366_, _11365_, _05955_);
  nand _62849_ (_11367_, _11366_, _11364_);
  or _62850_ (_11368_, _11367_, _06821_);
  and _62851_ (_11369_, _11366_, _11364_);
  and _62852_ (_11370_, _06746_, \oc8051_golden_model_1.PC [8]);
  and _62853_ (_11371_, _11370_, \oc8051_golden_model_1.PC [9]);
  and _62854_ (_11372_, _11371_, \oc8051_golden_model_1.PC [10]);
  and _62855_ (_11373_, _11372_, \oc8051_golden_model_1.PC [11]);
  and _62856_ (_11374_, _11373_, \oc8051_golden_model_1.PC [12]);
  and _62857_ (_11375_, _11374_, \oc8051_golden_model_1.PC [13]);
  and _62858_ (_11376_, _11375_, \oc8051_golden_model_1.PC [14]);
  nor _62859_ (_11377_, _11375_, \oc8051_golden_model_1.PC [14]);
  nor _62860_ (_11378_, _11377_, _11376_);
  not _62861_ (_11379_, _11378_);
  nor _62862_ (_11380_, _11379_, _05881_);
  and _62863_ (_11381_, _11379_, _05881_);
  nor _62864_ (_11382_, _11381_, _11380_);
  not _62865_ (_11383_, _11382_);
  nor _62866_ (_11384_, _11374_, \oc8051_golden_model_1.PC [13]);
  nor _62867_ (_11385_, _11384_, _11375_);
  not _62868_ (_11386_, _11385_);
  nor _62869_ (_11387_, _11386_, _05881_);
  and _62870_ (_11388_, _11386_, _05881_);
  nor _62871_ (_11389_, _11373_, \oc8051_golden_model_1.PC [12]);
  nor _62872_ (_11390_, _11389_, _11374_);
  not _62873_ (_11391_, _11390_);
  nor _62874_ (_11392_, _11391_, _05881_);
  nor _62875_ (_11393_, _11371_, \oc8051_golden_model_1.PC [10]);
  nor _62876_ (_11394_, _11393_, _11372_);
  not _62877_ (_11395_, _11394_);
  nor _62878_ (_11396_, _11395_, _05881_);
  not _62879_ (_11397_, _11396_);
  nor _62880_ (_11398_, _11372_, \oc8051_golden_model_1.PC [11]);
  nor _62881_ (_11399_, _11398_, _11373_);
  not _62882_ (_11400_, _11399_);
  nor _62883_ (_11401_, _11400_, _05881_);
  and _62884_ (_11402_, _11400_, _05881_);
  nor _62885_ (_11403_, _11402_, _11401_);
  and _62886_ (_11404_, _11395_, _05881_);
  nor _62887_ (_11405_, _11404_, _11396_);
  and _62888_ (_11406_, _11405_, _11403_);
  nor _62889_ (_11407_, _11370_, \oc8051_golden_model_1.PC [9]);
  nor _62890_ (_11408_, _11407_, _11371_);
  not _62891_ (_11409_, _11408_);
  nor _62892_ (_11410_, _11409_, _05881_);
  and _62893_ (_11411_, _11409_, _05881_);
  nor _62894_ (_11412_, _11411_, _11410_);
  nor _62895_ (_11413_, _06749_, _05881_);
  and _62896_ (_11414_, _06749_, _05881_);
  and _62897_ (_11415_, _06744_, _06077_);
  nor _62898_ (_11416_, _11415_, \oc8051_golden_model_1.PC [6]);
  nor _62899_ (_11417_, _11416_, _06745_);
  not _62900_ (_11418_, _11417_);
  nor _62901_ (_11419_, _11418_, _06204_);
  and _62902_ (_11420_, _11418_, _06204_);
  nor _62903_ (_11421_, _11420_, _11419_);
  not _62904_ (_11422_, _11421_);
  and _62905_ (_11423_, _06744_, \oc8051_golden_model_1.PC [4]);
  nor _62906_ (_11424_, _11423_, \oc8051_golden_model_1.PC [5]);
  nor _62907_ (_11425_, _11424_, _11415_);
  not _62908_ (_11426_, _11425_);
  nor _62909_ (_11427_, _11426_, _06267_);
  and _62910_ (_11428_, _11426_, _06267_);
  nor _62911_ (_11429_, _06744_, \oc8051_golden_model_1.PC [4]);
  nor _62912_ (_11430_, _11429_, _11423_);
  not _62913_ (_11431_, _11430_);
  nor _62914_ (_11432_, _11431_, _06236_);
  nor _62915_ (_11433_, _06743_, \oc8051_golden_model_1.PC [3]);
  nor _62916_ (_11434_, _11433_, _06744_);
  not _62917_ (_11435_, _11434_);
  nor _62918_ (_11436_, _11435_, _03708_);
  and _62919_ (_11437_, _11435_, _03708_);
  nor _62920_ (_11438_, _02909_, \oc8051_golden_model_1.PC [2]);
  nor _62921_ (_11439_, _11438_, _06743_);
  not _62922_ (_11440_, _11439_);
  nor _62923_ (_11441_, _11440_, _03946_);
  not _62924_ (_11442_, _03275_);
  nor _62925_ (_11443_, _04303_, _11442_);
  nor _62926_ (_11444_, _04163_, \oc8051_golden_model_1.PC [0]);
  and _62927_ (_11445_, _04303_, _11442_);
  nor _62928_ (_11446_, _11445_, _11443_);
  and _62929_ (_11447_, _11446_, _11444_);
  nor _62930_ (_11448_, _11447_, _11443_);
  and _62931_ (_11449_, _11440_, _03946_);
  nor _62932_ (_11450_, _11449_, _11441_);
  not _62933_ (_11451_, _11450_);
  nor _62934_ (_11452_, _11451_, _11448_);
  nor _62935_ (_11453_, _11452_, _11441_);
  nor _62936_ (_11454_, _11453_, _11437_);
  nor _62937_ (_11455_, _11454_, _11436_);
  and _62938_ (_11456_, _11431_, _06236_);
  nor _62939_ (_11457_, _11456_, _11432_);
  not _62940_ (_11458_, _11457_);
  nor _62941_ (_11459_, _11458_, _11455_);
  nor _62942_ (_11460_, _11459_, _11432_);
  nor _62943_ (_11461_, _11460_, _11428_);
  nor _62944_ (_11462_, _11461_, _11427_);
  nor _62945_ (_11463_, _11462_, _11422_);
  nor _62946_ (_11464_, _11463_, _11419_);
  nor _62947_ (_11465_, _11464_, _11414_);
  or _62948_ (_11466_, _11465_, _11413_);
  nor _62949_ (_11467_, _06746_, \oc8051_golden_model_1.PC [8]);
  nor _62950_ (_11468_, _11467_, _11370_);
  not _62951_ (_11469_, _11468_);
  nor _62952_ (_11470_, _11469_, _05881_);
  and _62953_ (_11471_, _11469_, _05881_);
  nor _62954_ (_11472_, _11471_, _11470_);
  and _62955_ (_11473_, _11472_, _11466_);
  and _62956_ (_11474_, _11473_, _11412_);
  and _62957_ (_11475_, _11474_, _11406_);
  nor _62958_ (_11476_, _11470_, _11410_);
  not _62959_ (_11477_, _11476_);
  and _62960_ (_11478_, _11477_, _11406_);
  or _62961_ (_11479_, _11478_, _11401_);
  nor _62962_ (_11480_, _11479_, _11475_);
  and _62963_ (_11481_, _11480_, _11397_);
  and _62964_ (_11482_, _11391_, _05881_);
  nor _62965_ (_11483_, _11482_, _11392_);
  not _62966_ (_11484_, _11483_);
  nor _62967_ (_11485_, _11484_, _11481_);
  nor _62968_ (_11486_, _11485_, _11392_);
  nor _62969_ (_11487_, _11486_, _11388_);
  nor _62970_ (_11488_, _11487_, _11387_);
  nor _62971_ (_11489_, _11488_, _11383_);
  nor _62972_ (_11490_, _11489_, _11380_);
  not _62973_ (_11491_, _06821_);
  and _62974_ (_11492_, _11491_, _05881_);
  nor _62975_ (_11493_, _11491_, _05881_);
  nor _62976_ (_11494_, _11493_, _11492_);
  and _62977_ (_11495_, _11494_, _11490_);
  nor _62978_ (_11496_, _11494_, _11490_);
  or _62979_ (_11497_, _11496_, _11495_);
  or _62980_ (_11498_, _11497_, _11369_);
  and _62981_ (_11499_, _11498_, _03610_);
  and _62982_ (_11500_, _11499_, _11368_);
  and _62983_ (_11501_, _05836_, _05834_);
  and _62984_ (_11502_, _04406_, _04620_);
  and _62985_ (_11503_, _06770_, _11502_);
  and _62986_ (_11504_, _11503_, _11501_);
  and _62987_ (_11505_, _11504_, _06813_);
  and _62988_ (_11506_, _06080_, \oc8051_golden_model_1.PC [8]);
  and _62989_ (_11507_, _11506_, \oc8051_golden_model_1.PC [9]);
  and _62990_ (_11508_, _11507_, \oc8051_golden_model_1.PC [10]);
  and _62991_ (_11509_, _11508_, \oc8051_golden_model_1.PC [11]);
  and _62992_ (_11510_, _11509_, \oc8051_golden_model_1.PC [12]);
  and _62993_ (_11511_, _11510_, \oc8051_golden_model_1.PC [13]);
  and _62994_ (_11512_, _11511_, \oc8051_golden_model_1.PC [14]);
  nor _62995_ (_11513_, _11511_, \oc8051_golden_model_1.PC [14]);
  nor _62996_ (_11514_, _11513_, _11512_);
  not _62997_ (_11515_, _11514_);
  nor _62998_ (_11516_, _11515_, _03446_);
  and _62999_ (_11517_, _11515_, _03446_);
  nor _63000_ (_11518_, _11517_, _11516_);
  not _63001_ (_11519_, _11518_);
  nor _63002_ (_11520_, _11510_, \oc8051_golden_model_1.PC [13]);
  nor _63003_ (_11521_, _11520_, _11511_);
  and _63004_ (_11522_, _11521_, _03454_);
  nor _63005_ (_11523_, _11521_, _03454_);
  nor _63006_ (_11524_, _11509_, \oc8051_golden_model_1.PC [12]);
  nor _63007_ (_11525_, _11524_, _11510_);
  not _63008_ (_11526_, _11525_);
  nor _63009_ (_11527_, _11526_, _03446_);
  nor _63010_ (_11528_, _11507_, \oc8051_golden_model_1.PC [10]);
  nor _63011_ (_11529_, _11528_, _11508_);
  and _63012_ (_11530_, _11529_, _03454_);
  not _63013_ (_11531_, _11530_);
  nor _63014_ (_11532_, _11508_, \oc8051_golden_model_1.PC [11]);
  nor _63015_ (_11533_, _11532_, _11509_);
  not _63016_ (_11534_, _11533_);
  nor _63017_ (_11535_, _11534_, _03446_);
  and _63018_ (_11536_, _11534_, _03446_);
  nor _63019_ (_11537_, _11536_, _11535_);
  nor _63020_ (_11538_, _11529_, _03454_);
  nor _63021_ (_11539_, _11538_, _11530_);
  and _63022_ (_11540_, _11539_, _11537_);
  nor _63023_ (_11541_, _11506_, \oc8051_golden_model_1.PC [9]);
  nor _63024_ (_11542_, _11541_, _11507_);
  not _63025_ (_11543_, _11542_);
  nor _63026_ (_11544_, _11543_, _03446_);
  and _63027_ (_11545_, _11543_, _03446_);
  nor _63028_ (_11546_, _11545_, _11544_);
  nor _63029_ (_11547_, _06143_, _03446_);
  and _63030_ (_11548_, _06143_, _03446_);
  and _63031_ (_11549_, _06077_, _03295_);
  nor _63032_ (_11550_, _11549_, \oc8051_golden_model_1.PC [6]);
  nor _63033_ (_11551_, _11550_, _06079_);
  not _63034_ (_11552_, _11551_);
  nor _63035_ (_11553_, _11552_, _03549_);
  and _63036_ (_11554_, _11552_, _03549_);
  nor _63037_ (_11555_, _11554_, _11553_);
  not _63038_ (_11556_, _11555_);
  and _63039_ (_11557_, _03295_, \oc8051_golden_model_1.PC [4]);
  nor _63040_ (_11558_, _11557_, \oc8051_golden_model_1.PC [5]);
  nor _63041_ (_11559_, _11558_, _11549_);
  not _63042_ (_11560_, _11559_);
  nor _63043_ (_11561_, _11560_, _03860_);
  and _63044_ (_11562_, _11560_, _03860_);
  nor _63045_ (_11563_, _03295_, \oc8051_golden_model_1.PC [4]);
  nor _63046_ (_11564_, _11563_, _11557_);
  not _63047_ (_11565_, _11564_);
  nor _63048_ (_11566_, _11565_, _03486_);
  nor _63049_ (_11567_, _03581_, _03648_);
  and _63050_ (_11568_, _03581_, _03648_);
  nor _63051_ (_11569_, _03904_, _03245_);
  nor _63052_ (_11570_, _03414_, \oc8051_golden_model_1.PC [1]);
  nor _63053_ (_11571_, _04048_, _02905_);
  and _63054_ (_11572_, _03414_, \oc8051_golden_model_1.PC [1]);
  nor _63055_ (_11573_, _11572_, _11570_);
  and _63056_ (_11574_, _11573_, _11571_);
  nor _63057_ (_11575_, _11574_, _11570_);
  and _63058_ (_11576_, _03904_, _03245_);
  nor _63059_ (_11577_, _11576_, _11569_);
  not _63060_ (_11578_, _11577_);
  nor _63061_ (_11579_, _11578_, _11575_);
  nor _63062_ (_11580_, _11579_, _11569_);
  nor _63063_ (_11581_, _11580_, _11568_);
  nor _63064_ (_11582_, _11581_, _11567_);
  and _63065_ (_11583_, _11565_, _03486_);
  nor _63066_ (_11584_, _11583_, _11566_);
  not _63067_ (_11585_, _11584_);
  nor _63068_ (_11586_, _11585_, _11582_);
  nor _63069_ (_11587_, _11586_, _11566_);
  nor _63070_ (_11588_, _11587_, _11562_);
  nor _63071_ (_11589_, _11588_, _11561_);
  nor _63072_ (_11590_, _11589_, _11556_);
  nor _63073_ (_11591_, _11590_, _11553_);
  nor _63074_ (_11592_, _11591_, _11548_);
  or _63075_ (_11593_, _11592_, _11547_);
  nor _63076_ (_11594_, _06080_, \oc8051_golden_model_1.PC [8]);
  nor _63077_ (_11595_, _11594_, _11506_);
  not _63078_ (_11596_, _11595_);
  nor _63079_ (_11597_, _11596_, _03446_);
  and _63080_ (_11598_, _11596_, _03446_);
  nor _63081_ (_11599_, _11598_, _11597_);
  and _63082_ (_11600_, _11599_, _11593_);
  and _63083_ (_11601_, _11600_, _11546_);
  and _63084_ (_11602_, _11601_, _11540_);
  nor _63085_ (_11603_, _11597_, _11544_);
  not _63086_ (_11604_, _11603_);
  and _63087_ (_11605_, _11604_, _11540_);
  or _63088_ (_11606_, _11605_, _11535_);
  nor _63089_ (_11607_, _11606_, _11602_);
  and _63090_ (_11608_, _11607_, _11531_);
  and _63091_ (_11609_, _11526_, _03446_);
  nor _63092_ (_11610_, _11609_, _11527_);
  not _63093_ (_11611_, _11610_);
  nor _63094_ (_11612_, _11611_, _11608_);
  nor _63095_ (_11613_, _11612_, _11527_);
  nor _63096_ (_11614_, _11613_, _11523_);
  nor _63097_ (_11615_, _11614_, _11522_);
  nor _63098_ (_11616_, _11615_, _11519_);
  nor _63099_ (_11617_, _11616_, _11516_);
  and _63100_ (_11618_, _06814_, _03446_);
  nor _63101_ (_11619_, _06814_, _03446_);
  nor _63102_ (_11620_, _11619_, _11618_);
  and _63103_ (_11621_, _11620_, _11617_);
  nor _63104_ (_11622_, _11620_, _11617_);
  or _63105_ (_11623_, _11622_, _11621_);
  nand _63106_ (_11624_, _11503_, _11501_);
  and _63107_ (_11625_, _11624_, _11623_);
  or _63108_ (_11626_, _11625_, _06072_);
  or _63109_ (_11627_, _11626_, _11505_);
  nor _63110_ (_11628_, _04622_, _03234_);
  not _63111_ (_11629_, _11628_);
  and _63112_ (_11630_, _11629_, _08078_);
  not _63113_ (_11631_, _11630_);
  and _63114_ (_11632_, _03979_, _02994_);
  nand _63115_ (_11633_, _06814_, _03979_);
  nor _63116_ (_11634_, _04729_, _03980_);
  nor _63117_ (_11635_, _04409_, \oc8051_golden_model_1.PC [15]);
  nand _63118_ (_11636_, _11635_, _11634_);
  and _63119_ (_11637_, _11636_, _11633_);
  or _63120_ (_11638_, _11637_, _11632_);
  nand _63121_ (_11639_, _06814_, _03980_);
  and _63122_ (_11640_, _11639_, _11638_);
  or _63123_ (_11641_, _11640_, _11631_);
  nor _63124_ (_11642_, _04729_, _11632_);
  and _63125_ (_11643_, _11642_, _11630_);
  or _63126_ (_11644_, _11643_, _11327_);
  and _63127_ (_11645_, _11644_, _11641_);
  or _63128_ (_11646_, _11645_, _06073_);
  nor _63129_ (_11647_, _04422_, _03610_);
  and _63130_ (_11648_, _11647_, _11646_);
  and _63131_ (_11649_, _11648_, _11627_);
  or _63132_ (_11650_, _11649_, _11500_);
  and _63133_ (_11651_, _11650_, _11362_);
  not _63134_ (_11652_, _11360_);
  and _63135_ (_11653_, _11362_, _05966_);
  not _63136_ (_11654_, _11653_);
  and _63137_ (_11655_, _11654_, _11327_);
  or _63138_ (_11656_, _11655_, _11652_);
  or _63139_ (_11657_, _11656_, _11651_);
  and _63140_ (_11658_, _11657_, _11361_);
  and _63141_ (_11659_, _08063_, _08128_);
  not _63142_ (_11660_, _11659_);
  or _63143_ (_11661_, _11660_, _11658_);
  or _63144_ (_11662_, _11659_, _11327_);
  and _63145_ (_11663_, _11662_, _03737_);
  and _63146_ (_11664_, _11663_, _11661_);
  or _63147_ (_11665_, _11664_, _11359_);
  nor _63148_ (_11666_, _09909_, _08132_);
  and _63149_ (_11667_, _11666_, _11665_);
  not _63150_ (_11668_, _11666_);
  and _63151_ (_11669_, _11668_, _11327_);
  not _63152_ (_11670_, _03233_);
  nor _63153_ (_11671_, _03508_, _11670_);
  and _63154_ (_11672_, _11671_, _03736_);
  not _63155_ (_11673_, _11672_);
  or _63156_ (_11674_, _11673_, _11669_);
  or _63157_ (_11675_, _11674_, _11667_);
  or _63158_ (_11676_, _11672_, _06813_);
  and _63159_ (_11677_, _11676_, _09921_);
  and _63160_ (_11678_, _11677_, _11675_);
  or _63161_ (_11679_, _11497_, _09969_);
  nand _63162_ (_11680_, _09969_, _11491_);
  and _63163_ (_11681_, _11680_, _09917_);
  and _63164_ (_11682_, _11681_, _11679_);
  or _63165_ (_11683_, _11682_, _09919_);
  or _63166_ (_11684_, _11683_, _11678_);
  and _63167_ (_11685_, _10017_, _10006_);
  and _63168_ (_11686_, _11685_, _06821_);
  and _63169_ (_11687_, _11497_, _10018_);
  or _63170_ (_11688_, _11687_, _11686_);
  or _63171_ (_11689_, _11688_, _09920_);
  and _63172_ (_11690_, _11689_, _11684_);
  or _63173_ (_11691_, _11690_, _03615_);
  and _63174_ (_11692_, _09876_, _06821_);
  not _63175_ (_11693_, _09876_);
  and _63176_ (_11694_, _11497_, _11693_);
  or _63177_ (_11695_, _11694_, _04107_);
  or _63178_ (_11696_, _11695_, _11692_);
  and _63179_ (_11697_, _11696_, _09856_);
  and _63180_ (_11698_, _11697_, _11691_);
  or _63181_ (_11699_, _11497_, _10061_);
  nand _63182_ (_11700_, _10061_, _11491_);
  and _63183_ (_11701_, _11700_, _03604_);
  and _63184_ (_11702_, _11701_, _11699_);
  or _63185_ (_11703_, _11702_, _11698_);
  and _63186_ (_11704_, _11703_, _11358_);
  nand _63187_ (_11705_, _11327_, _10025_);
  nor _63188_ (_11706_, _04746_, _03718_);
  and _63189_ (_11707_, _11706_, _03227_);
  and _63190_ (_11708_, _03593_, _03751_);
  not _63191_ (_11709_, _11708_);
  and _63192_ (_11710_, _11709_, _11707_);
  nor _63193_ (_11711_, _08070_, _03237_);
  not _63194_ (_11712_, _11711_);
  nor _63195_ (_11713_, _03616_, _03494_);
  nor _63196_ (_11714_, _11713_, _03237_);
  and _63197_ (_11715_, _04066_, _03751_);
  or _63198_ (_11716_, _04115_, _03719_);
  or _63199_ (_11717_, _11716_, _11715_);
  nor _63200_ (_11718_, _11717_, _11714_);
  and _63201_ (_11719_, _11718_, _11712_);
  and _63202_ (_11720_, _11719_, _11710_);
  nand _63203_ (_11721_, _11720_, _11705_);
  or _63204_ (_11722_, _11721_, _11704_);
  or _63205_ (_11723_, _11720_, _06813_);
  and _63206_ (_11724_, _11723_, _11355_);
  and _63207_ (_11725_, _11724_, _11722_);
  or _63208_ (_11726_, _11725_, _11357_);
  not _63209_ (_11727_, _03238_);
  nor _63210_ (_11728_, _03752_, _11727_);
  and _63211_ (_11729_, _11728_, _09669_);
  and _63212_ (_11730_, _11729_, _11726_);
  or _63213_ (_11731_, _11729_, _06814_);
  nand _63214_ (_11732_, _11731_, _11350_);
  or _63215_ (_11733_, _11732_, _11730_);
  and _63216_ (_11734_, _11733_, _11351_);
  or _63217_ (_11735_, _11734_, _08187_);
  or _63218_ (_11736_, _08186_, _06813_);
  and _63219_ (_11737_, _11736_, _03248_);
  and _63220_ (_11738_, _11737_, _11735_);
  and _63221_ (_11739_, _11327_, _07912_);
  nor _63222_ (_11740_, _03505_, _03224_);
  not _63223_ (_11741_, _11740_);
  or _63224_ (_11742_, _11741_, _11739_);
  or _63225_ (_11743_, _11742_, _11738_);
  or _63226_ (_11744_, _11740_, _06813_);
  and _63227_ (_11745_, _11744_, _08832_);
  and _63228_ (_11746_, _11745_, _11743_);
  nand _63229_ (_11747_, _06821_, _03625_);
  nor _63230_ (_11748_, _04481_, _06833_);
  and _63231_ (_11749_, _11748_, _06837_);
  nand _63232_ (_11750_, _11749_, _11747_);
  or _63233_ (_11751_, _11750_, _11746_);
  or _63234_ (_11752_, _11749_, _06813_);
  and _63235_ (_11753_, _11752_, _03589_);
  and _63236_ (_11754_, _11753_, _11751_);
  or _63237_ (_11755_, _11754_, _11349_);
  nor _63238_ (_11756_, _07405_, _03216_);
  and _63239_ (_11757_, _11756_, _11755_);
  not _63240_ (_11758_, _11756_);
  and _63241_ (_11759_, _11758_, _11327_);
  nor _63242_ (_11760_, _03585_, _03169_);
  not _63243_ (_11761_, _11760_);
  or _63244_ (_11762_, _11761_, _11759_);
  or _63245_ (_11763_, _11762_, _11757_);
  and _63246_ (_11764_, _03168_, _03452_);
  not _63247_ (_11765_, _11764_);
  or _63248_ (_11766_, _11760_, _06813_);
  and _63249_ (_11767_, _11766_, _11765_);
  and _63250_ (_11768_, _11767_, _11763_);
  and _63251_ (_11769_, _11764_, _11623_);
  or _63252_ (_11770_, _11769_, _06168_);
  or _63253_ (_11771_, _11770_, _11768_);
  or _63254_ (_11772_, _06813_, _05894_);
  and _63255_ (_11773_, _11772_, _11771_);
  or _63256_ (_11774_, _11773_, _03601_);
  nand _63257_ (_11775_, _11491_, _03601_);
  and _63258_ (_11776_, _11775_, _08364_);
  and _63259_ (_11777_, _11776_, _11774_);
  and _63260_ (_11778_, _08363_, _06813_);
  or _63261_ (_11779_, _11778_, _11777_);
  and _63262_ (_11780_, _11779_, _11348_);
  and _63263_ (_11781_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor _63264_ (_11782_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and _63265_ (_11783_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63266_ (_11784_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63267_ (_11785_, _11784_, _11783_);
  not _63268_ (_11786_, _11785_);
  and _63269_ (_11787_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63270_ (_11788_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63271_ (_11789_, _11788_, _11787_);
  not _63272_ (_11790_, _11789_);
  and _63273_ (_11791_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63274_ (_11792_, _03305_, _03301_);
  nor _63275_ (_11793_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63276_ (_11794_, _11793_, _11791_);
  not _63277_ (_11795_, _11794_);
  nor _63278_ (_11796_, _11795_, _11792_);
  nor _63279_ (_11797_, _11796_, _11791_);
  nor _63280_ (_11798_, _11797_, _11790_);
  nor _63281_ (_11799_, _11798_, _11787_);
  nor _63282_ (_11800_, _11799_, _11786_);
  nor _63283_ (_11801_, _11800_, _11783_);
  nor _63284_ (_11802_, _11801_, _11782_);
  or _63285_ (_11803_, _11802_, _11781_);
  and _63286_ (_11804_, _11803_, \oc8051_golden_model_1.DPH [0]);
  and _63287_ (_11805_, _11804_, \oc8051_golden_model_1.DPH [1]);
  and _63288_ (_11806_, _11805_, \oc8051_golden_model_1.DPH [2]);
  and _63289_ (_11807_, _11806_, \oc8051_golden_model_1.DPH [3]);
  and _63290_ (_11808_, _11807_, \oc8051_golden_model_1.DPH [4]);
  and _63291_ (_11809_, _11808_, \oc8051_golden_model_1.DPH [5]);
  and _63292_ (_11810_, _11809_, \oc8051_golden_model_1.DPH [6]);
  nand _63293_ (_11811_, _11810_, \oc8051_golden_model_1.DPH [7]);
  or _63294_ (_11812_, _11810_, \oc8051_golden_model_1.DPH [7]);
  and _63295_ (_11813_, _11812_, _11347_);
  and _63296_ (_11814_, _11813_, _11811_);
  nor _63297_ (_11815_, _03584_, _03178_);
  not _63298_ (_11816_, _11815_);
  or _63299_ (_11817_, _11816_, _11814_);
  or _63300_ (_11818_, _11817_, _11780_);
  and _63301_ (_11819_, _03176_, _03452_);
  not _63302_ (_11820_, _11819_);
  or _63303_ (_11821_, _11815_, _06813_);
  and _63304_ (_11822_, _11821_, _11820_);
  and _63305_ (_11823_, _11822_, _11818_);
  not _63306_ (_11824_, _11345_);
  or _63307_ (_11825_, _11623_, _08786_);
  not _63308_ (_11826_, _08786_);
  or _63309_ (_11827_, _11826_, _06813_);
  and _63310_ (_11828_, _11827_, _11819_);
  and _63311_ (_11829_, _11828_, _11825_);
  or _63312_ (_11830_, _11829_, _11824_);
  or _63313_ (_11831_, _11830_, _11823_);
  and _63314_ (_11832_, _11831_, _11346_);
  or _63315_ (_11833_, _11832_, _11342_);
  or _63316_ (_11834_, _11341_, _06813_);
  and _63317_ (_11835_, _11834_, _07766_);
  and _63318_ (_11836_, _11835_, _11833_);
  nand _63319_ (_11837_, _06821_, _03600_);
  nor _63320_ (_11838_, _03780_, _03182_);
  nand _63321_ (_11839_, _11838_, _11837_);
  or _63322_ (_11840_, _11839_, _11836_);
  and _63323_ (_11841_, _03181_, _03452_);
  not _63324_ (_11842_, _11841_);
  or _63325_ (_11843_, _11838_, _06813_);
  and _63326_ (_11844_, _11843_, _11842_);
  and _63327_ (_11845_, _11844_, _11840_);
  or _63328_ (_11846_, _11623_, _11826_);
  or _63329_ (_11847_, _08786_, _06813_);
  and _63330_ (_11848_, _11847_, _11841_);
  and _63331_ (_11849_, _11848_, _11846_);
  or _63332_ (_11850_, _11849_, _11845_);
  and _63333_ (_11851_, _08425_, _08417_);
  and _63334_ (_11852_, _11851_, _11850_);
  not _63335_ (_11853_, _11851_);
  and _63336_ (_11854_, _11853_, _11327_);
  or _63337_ (_11855_, _11854_, _08431_);
  or _63338_ (_11856_, _11855_, _11852_);
  or _63339_ (_11857_, _08430_, _06813_);
  and _63340_ (_11858_, _11857_, _07777_);
  and _63341_ (_11859_, _11858_, _11856_);
  nand _63342_ (_11860_, _06821_, _03622_);
  nand _63343_ (_11861_, _11860_, _10753_);
  or _63344_ (_11862_, _11861_, _11859_);
  and _63345_ (_11863_, _11862_, _11340_);
  not _63346_ (_11864_, _11335_);
  or _63347_ (_11865_, _11623_, \oc8051_golden_model_1.PSW [7]);
  or _63348_ (_11866_, _06813_, _07871_);
  and _63349_ (_11867_, _11866_, _11337_);
  and _63350_ (_11868_, _11867_, _11865_);
  or _63351_ (_11869_, _11868_, _11864_);
  or _63352_ (_11870_, _11869_, _11863_);
  and _63353_ (_11871_, _11870_, _11336_);
  or _63354_ (_11872_, _11871_, _08460_);
  or _63355_ (_11873_, _08459_, _06813_);
  and _63356_ (_11874_, _11873_, _07795_);
  and _63357_ (_11875_, _11874_, _11872_);
  nand _63358_ (_11876_, _06821_, _03624_);
  nor _63359_ (_11877_, _03785_, _03201_);
  nand _63360_ (_11878_, _11877_, _11876_);
  or _63361_ (_11879_, _11878_, _11875_);
  and _63362_ (_11880_, _03200_, _03452_);
  not _63363_ (_11881_, _11880_);
  or _63364_ (_11882_, _11877_, _06813_);
  and _63365_ (_11883_, _11882_, _11881_);
  and _63366_ (_11884_, _11883_, _11879_);
  not _63367_ (_11885_, _11330_);
  or _63368_ (_11886_, _11623_, _07871_);
  or _63369_ (_11887_, _06813_, \oc8051_golden_model_1.PSW [7]);
  and _63370_ (_11888_, _11887_, _11880_);
  and _63371_ (_11889_, _11888_, _11886_);
  or _63372_ (_11890_, _11889_, _11885_);
  or _63373_ (_11891_, _11890_, _11884_);
  and _63374_ (_11892_, _11891_, _11331_);
  or _63375_ (_11893_, _11892_, _08508_);
  or _63376_ (_11894_, _08507_, _06813_);
  and _63377_ (_11895_, _11894_, _08588_);
  and _63378_ (_11896_, _11895_, _11893_);
  and _63379_ (_11897_, _11327_, _08587_);
  or _63380_ (_11898_, _11897_, _03798_);
  or _63381_ (_11899_, _11898_, _11896_);
  nand _63382_ (_11900_, _05204_, _03798_);
  and _63383_ (_11901_, _11900_, _11899_);
  or _63384_ (_11902_, _11901_, _03188_);
  not _63385_ (_11903_, _03621_);
  nand _63386_ (_11904_, _06814_, _03188_);
  and _63387_ (_11905_, _11904_, _11903_);
  and _63388_ (_11906_, _11905_, _11902_);
  not _63389_ (_11907_, _11328_);
  not _63390_ (_11908_, _09854_);
  or _63391_ (_11909_, _11497_, _11908_);
  or _63392_ (_11910_, _09854_, _06821_);
  and _63393_ (_11911_, _11910_, _03621_);
  and _63394_ (_11912_, _11911_, _11909_);
  or _63395_ (_11913_, _11912_, _11907_);
  or _63396_ (_11914_, _11913_, _11906_);
  and _63397_ (_11915_, _11914_, _11329_);
  or _63398_ (_11916_, _11915_, _08703_);
  or _63399_ (_11917_, _08702_, _06813_);
  and _63400_ (_11918_, _11917_, _08733_);
  and _63401_ (_11919_, _11918_, _11916_);
  and _63402_ (_11920_, _11327_, _08732_);
  or _63403_ (_11921_, _11920_, _03515_);
  or _63404_ (_11922_, _11921_, _11919_);
  nand _63405_ (_11923_, _05204_, _03515_);
  and _63406_ (_11924_, _11923_, _11922_);
  or _63407_ (_11925_, _11924_, _03203_);
  nand _63408_ (_11926_, _06814_, _03203_);
  and _63409_ (_11927_, _11926_, _03816_);
  and _63410_ (_11928_, _11927_, _11925_);
  or _63411_ (_11929_, _11497_, _09854_);
  nand _63412_ (_11930_, _09854_, _11491_);
  and _63413_ (_11931_, _11930_, _11929_);
  and _63414_ (_11932_, _11931_, _03628_);
  and _63415_ (_11933_, _05848_, _06409_);
  not _63416_ (_11934_, _11933_);
  or _63417_ (_11935_, _11934_, _11932_);
  or _63418_ (_11936_, _11935_, _11928_);
  or _63419_ (_11937_, _11933_, _11327_);
  and _63420_ (_11938_, _11937_, _04246_);
  and _63421_ (_11939_, _11938_, _11936_);
  nor _63422_ (_11940_, _08780_, _08775_);
  nand _63423_ (_11941_, _06813_, _03815_);
  nand _63424_ (_11942_, _11941_, _11940_);
  or _63425_ (_11943_, _11942_, _11939_);
  not _63426_ (_11944_, _03629_);
  or _63427_ (_11945_, _11327_, _11940_);
  and _63428_ (_11946_, _11945_, _11944_);
  and _63429_ (_11947_, _11946_, _11943_);
  nor _63430_ (_11948_, _11944_, _03446_);
  or _63431_ (_11949_, _11948_, _03198_);
  or _63432_ (_11950_, _11949_, _11947_);
  nand _63433_ (_11951_, _06814_, _03198_);
  and _63434_ (_11952_, _11951_, _03823_);
  and _63435_ (_11953_, _11952_, _11950_);
  and _63436_ (_11954_, _11931_, _03453_);
  nand _63437_ (_11955_, _03195_, _02962_);
  not _63438_ (_11956_, _11955_);
  nor _63439_ (_11957_, _11956_, _04552_);
  not _63440_ (_11958_, _11957_);
  or _63441_ (_11959_, _11958_, _11954_);
  or _63442_ (_11960_, _11959_, _11953_);
  or _63443_ (_11961_, _11957_, _11327_);
  and _63444_ (_11962_, _11961_, _03514_);
  and _63445_ (_11963_, _11962_, _11960_);
  nor _63446_ (_11964_, _08805_, _08798_);
  nand _63447_ (_11965_, _06813_, _03447_);
  nand _63448_ (_11966_, _11965_, _11964_);
  or _63449_ (_11967_, _11966_, _11963_);
  not _63450_ (_11968_, _03631_);
  or _63451_ (_11969_, _11327_, _11964_);
  and _63452_ (_11970_, _11969_, _11968_);
  and _63453_ (_11971_, _11970_, _11967_);
  nor _63454_ (_11972_, _11968_, _03446_);
  or _63455_ (_11973_, _11972_, _03196_);
  or _63456_ (_11974_, _11973_, _11971_);
  and _63457_ (_11975_, _03195_, _03452_);
  not _63458_ (_11976_, _11975_);
  nand _63459_ (_11977_, _06814_, _03196_);
  and _63460_ (_11978_, _11977_, _11976_);
  and _63461_ (_11979_, _11978_, _11974_);
  and _63462_ (_11980_, _11975_, _11327_);
  or _63463_ (_11981_, _11980_, _11979_);
  or _63464_ (_11982_, _11981_, _43004_);
  or _63465_ (_11983_, _43000_, \oc8051_golden_model_1.PC [15]);
  and _63466_ (_11984_, _11983_, _41806_);
  and _63467_ (_40591_, _11984_, _11982_);
  and _63468_ (_11985_, _43004_, \oc8051_golden_model_1.P0INREG [7]);
  or _63469_ (_11986_, _11985_, _01195_);
  and _63470_ (_40592_, _11986_, _41806_);
  and _63471_ (_11987_, _43004_, \oc8051_golden_model_1.P1INREG [7]);
  or _63472_ (_11988_, _11987_, _01092_);
  and _63473_ (_40593_, _11988_, _41806_);
  and _63474_ (_11989_, _43004_, \oc8051_golden_model_1.P2INREG [7]);
  or _63475_ (_11990_, _11989_, _00908_);
  and _63476_ (_40595_, _11990_, _41806_);
  and _63477_ (_11991_, _43004_, \oc8051_golden_model_1.P3INREG [7]);
  or _63478_ (_11992_, _11991_, _01028_);
  and _63479_ (_40596_, _11992_, _41806_);
  nor _63480_ (_11993_, _04797_, _04556_);
  nor _63481_ (_11994_, _11993_, _04798_);
  nor _63482_ (_11995_, _04797_, _04951_);
  nor _63483_ (_11996_, _11995_, _05123_);
  and _63484_ (_11997_, _11996_, _04796_);
  and _63485_ (_11998_, _11997_, _11994_);
  not _63486_ (_11999_, _11998_);
  nand _63487_ (_12000_, _03198_, _02905_);
  or _63488_ (_12001_, _04533_, _04634_);
  and _63489_ (_12002_, _12001_, _11934_);
  nor _63490_ (_12003_, _05666_, \oc8051_golden_model_1.ACC [0]);
  nand _63491_ (_12004_, _12003_, _06394_);
  and _63492_ (_12005_, _05666_, \oc8051_golden_model_1.ACC [0]);
  or _63493_ (_12006_, _12005_, _06382_);
  or _63494_ (_12007_, _04480_, _04620_);
  nand _63495_ (_12008_, _08285_, _03745_);
  nor _63496_ (_12009_, _10122_, _05224_);
  or _63497_ (_12010_, _12009_, _05940_);
  or _63498_ (_12011_, _06072_, _04634_);
  nand _63499_ (_12012_, _03980_, _02905_);
  or _63500_ (_12013_, _03980_, \oc8051_golden_model_1.ACC [0]);
  and _63501_ (_12014_, _12013_, _12012_);
  nor _63502_ (_12015_, _12014_, _06073_);
  nor _63503_ (_12016_, _12015_, _04421_);
  and _63504_ (_12017_, _12016_, _12011_);
  nor _63505_ (_12018_, _05666_, _06071_);
  or _63506_ (_12019_, _12018_, _12017_);
  and _63507_ (_12020_, _12019_, _05954_);
  nand _63508_ (_12021_, _10122_, _09750_);
  and _63509_ (_12022_, _12021_, _04428_);
  or _63510_ (_12023_, _12022_, _04768_);
  or _63511_ (_12024_, _12023_, _12020_);
  nor _63512_ (_12025_, _03230_, \oc8051_golden_model_1.PC [0]);
  nor _63513_ (_12026_, _12025_, _04431_);
  and _63514_ (_12027_, _12026_, _12024_);
  and _63515_ (_12028_, _04431_, _04620_);
  or _63516_ (_12029_, _12028_, _04449_);
  or _63517_ (_12030_, _12029_, _12027_);
  and _63518_ (_12031_, _12030_, _12010_);
  or _63519_ (_12032_, _12031_, _03508_);
  nand _63520_ (_12033_, _08285_, _03508_);
  and _63521_ (_12034_, _12033_, _04562_);
  and _63522_ (_12035_, _12034_, _12032_);
  nor _63523_ (_12036_, _10123_, _04562_);
  and _63524_ (_12037_, _12036_, _12021_);
  or _63525_ (_12038_, _12037_, _12035_);
  and _63526_ (_12039_, _12038_, _03227_);
  nor _63527_ (_12040_, _03227_, _02905_);
  or _63528_ (_12041_, _03745_, _12040_);
  or _63529_ (_12042_, _12041_, _12039_);
  and _63530_ (_12043_, _12042_, _12008_);
  or _63531_ (_12044_, _12043_, _04463_);
  and _63532_ (_12045_, _06546_, _03446_);
  nand _63533_ (_12046_, _08284_, _04463_);
  or _63534_ (_12047_, _12046_, _12045_);
  and _63535_ (_12048_, _12047_, _12044_);
  or _63536_ (_12049_, _12048_, _04462_);
  nor _63537_ (_12050_, _09773_, _05224_);
  and _63538_ (_12051_, _05224_, \oc8051_golden_model_1.PSW [7]);
  nor _63539_ (_12052_, _12051_, _12050_);
  nand _63540_ (_12053_, _12052_, _04462_);
  and _63541_ (_12054_, _12053_, _05897_);
  and _63542_ (_12055_, _12054_, _12049_);
  nand _63543_ (_12056_, _03224_, \oc8051_golden_model_1.PC [0]);
  nand _63544_ (_12057_, _04480_, _12056_);
  or _63545_ (_12058_, _12057_, _12055_);
  and _63546_ (_12059_, _12058_, _12007_);
  or _63547_ (_12060_, _12059_, _04482_);
  or _63548_ (_12061_, _06546_, _06164_);
  and _63549_ (_12062_, _12061_, _06163_);
  and _63550_ (_12063_, _12062_, _12060_);
  and _63551_ (_12064_, _05881_, _04620_);
  and _63552_ (_12065_, _06340_, \oc8051_golden_model_1.P1INREG [0]);
  not _63553_ (_12066_, _12065_);
  and _63554_ (_12067_, _06343_, \oc8051_golden_model_1.P0INREG [0]);
  not _63555_ (_12068_, _12067_);
  and _63556_ (_12069_, _06346_, \oc8051_golden_model_1.P2INREG [0]);
  and _63557_ (_12070_, _06348_, \oc8051_golden_model_1.P3INREG [0]);
  nor _63558_ (_12071_, _12070_, _12069_);
  and _63559_ (_12072_, _12071_, _12068_);
  and _63560_ (_12073_, _12072_, _12066_);
  and _63561_ (_12074_, _06354_, \oc8051_golden_model_1.SP [0]);
  and _63562_ (_12075_, _06284_, \oc8051_golden_model_1.TL0 [0]);
  nor _63563_ (_12076_, _12075_, _12074_);
  and _63564_ (_12077_, _12076_, _12073_);
  and _63565_ (_12078_, _06315_, \oc8051_golden_model_1.IE [0]);
  and _63566_ (_12079_, _06319_, \oc8051_golden_model_1.SBUF [0]);
  and _63567_ (_12080_, _06321_, \oc8051_golden_model_1.SCON [0]);
  or _63568_ (_12081_, _12080_, _12079_);
  nor _63569_ (_12082_, _12081_, _12078_);
  and _63570_ (_12083_, _06296_, \oc8051_golden_model_1.IP [0]);
  and _63571_ (_12084_, _06310_, \oc8051_golden_model_1.B [0]);
  nor _63572_ (_12085_, _12084_, _12083_);
  and _63573_ (_12086_, _06303_, \oc8051_golden_model_1.PSW [0]);
  and _63574_ (_12087_, _06308_, \oc8051_golden_model_1.ACC [0]);
  nor _63575_ (_12088_, _12087_, _12086_);
  and _63576_ (_12089_, _12088_, _12085_);
  and _63577_ (_12090_, _12089_, _12082_);
  and _63578_ (_12091_, _12090_, _12077_);
  and _63579_ (_12092_, _06327_, \oc8051_golden_model_1.TH0 [0]);
  and _63580_ (_12093_, _06329_, \oc8051_golden_model_1.TL1 [0]);
  nor _63581_ (_12094_, _12093_, _12092_);
  and _63582_ (_12095_, _06334_, \oc8051_golden_model_1.PCON [0]);
  and _63583_ (_12096_, _06336_, \oc8051_golden_model_1.TCON [0]);
  nor _63584_ (_12097_, _12096_, _12095_);
  and _63585_ (_12098_, _12097_, _12094_);
  and _63586_ (_12099_, _06272_, \oc8051_golden_model_1.DPH [0]);
  and _63587_ (_12100_, _06279_, \oc8051_golden_model_1.TMOD [0]);
  nor _63588_ (_12101_, _12100_, _12099_);
  and _63589_ (_12102_, _06356_, \oc8051_golden_model_1.DPL [0]);
  and _63590_ (_12103_, _06288_, \oc8051_golden_model_1.TH1 [0]);
  nor _63591_ (_12104_, _12103_, _12102_);
  and _63592_ (_12105_, _12104_, _12101_);
  and _63593_ (_12106_, _12105_, _12098_);
  and _63594_ (_12107_, _12106_, _12091_);
  not _63595_ (_12108_, _12107_);
  nor _63596_ (_12109_, _12108_, _12064_);
  nor _63597_ (_12110_, _12109_, _06170_);
  or _63598_ (_12111_, _12110_, _06168_);
  or _63599_ (_12112_, _12111_, _12063_);
  and _63600_ (_12113_, _06168_, _04048_);
  nor _63601_ (_12114_, _12113_, _04500_);
  and _63602_ (_12115_, _12114_, _12112_);
  and _63603_ (_12116_, _04500_, _06274_);
  or _63604_ (_12117_, _12116_, _03178_);
  or _63605_ (_12118_, _12117_, _12115_);
  and _63606_ (_12119_, _03178_, _02905_);
  nor _63607_ (_12120_, _12119_, _04512_);
  and _63608_ (_12121_, _12120_, _12118_);
  nor _63609_ (_12122_, _05666_, _06274_);
  and _63610_ (_12123_, _05666_, _06274_);
  nor _63611_ (_12124_, _12123_, _12122_);
  nor _63612_ (_12125_, _12124_, _04511_);
  nor _63613_ (_12126_, _12125_, _04513_);
  or _63614_ (_12127_, _12126_, _12121_);
  nor _63615_ (_12128_, _12005_, _12003_);
  or _63616_ (_12129_, _12128_, _05850_);
  and _63617_ (_12130_, _12129_, _06383_);
  and _63618_ (_12131_, _12130_, _12127_);
  and _63619_ (_12132_, _12123_, _04515_);
  or _63620_ (_12133_, _12132_, _04514_);
  or _63621_ (_12134_, _12133_, _12131_);
  and _63622_ (_12135_, _12134_, _12006_);
  or _63623_ (_12136_, _12135_, _03192_);
  and _63624_ (_12137_, _03192_, _02905_);
  nor _63625_ (_12138_, _12137_, _06390_);
  and _63626_ (_12139_, _12138_, _12136_);
  nor _63627_ (_12140_, _12122_, _06395_);
  or _63628_ (_12141_, _12140_, _06394_);
  or _63629_ (_12142_, _12141_, _12139_);
  and _63630_ (_12143_, _12142_, _12004_);
  or _63631_ (_12144_, _12143_, _03188_);
  nand _63632_ (_12145_, _03188_, _02905_);
  and _63633_ (_12146_, _12145_, _05848_);
  and _63634_ (_12147_, _12146_, _12144_);
  or _63635_ (_12148_, _12147_, _12002_);
  nand _63636_ (_12149_, _06546_, _04533_);
  and _63637_ (_12150_, _12149_, _12148_);
  or _63638_ (_12151_, _12150_, _04531_);
  nand _63639_ (_12152_, _05666_, _04531_);
  and _63640_ (_12153_, _12152_, _11944_);
  and _63641_ (_12154_, _12153_, _12151_);
  and _63642_ (_12155_, _03629_, _02905_);
  or _63643_ (_12156_, _12155_, _03198_);
  or _63644_ (_12157_, _12156_, _12154_);
  and _63645_ (_12158_, _12157_, _12000_);
  or _63646_ (_12159_, _12158_, _04539_);
  or _63647_ (_12160_, _12050_, _04558_);
  and _63648_ (_12161_, _12160_, _11955_);
  and _63649_ (_12162_, _12161_, _12159_);
  or _63650_ (_12163_, _04552_, _04634_);
  and _63651_ (_12164_, _12163_, _11958_);
  or _63652_ (_12165_, _12164_, _12162_);
  nand _63653_ (_12166_, _06546_, _04552_);
  and _63654_ (_12167_, _12166_, _12165_);
  or _63655_ (_12168_, _12167_, _03448_);
  nand _63656_ (_12169_, _05666_, _03448_);
  and _63657_ (_12170_, _12169_, _04796_);
  and _63658_ (_12171_, _12170_, _12168_);
  or _63659_ (_12172_, _12171_, _11999_);
  not _63660_ (_12173_, _00000_);
  nor _63661_ (_12174_, _04793_, _12173_);
  not _63662_ (_12175_, _12174_);
  nor _63663_ (_12176_, _04951_, _12175_);
  nor _63664_ (_12177_, _05122_, _12175_);
  nor _63665_ (_12178_, _12177_, _12176_);
  nor _63666_ (_12179_, _12175_, _04556_);
  nor _63667_ (_12180_, _12175_, _04711_);
  nor _63668_ (_12181_, _12180_, _12179_);
  and _63669_ (_12182_, _12181_, _12174_);
  and _63670_ (_12183_, _12182_, _12178_);
  or _63671_ (_12184_, _12183_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _63672_ (_12185_, _05137_, _05129_);
  nor _63673_ (_12186_, _12185_, _05138_);
  and _63674_ (_12187_, _12186_, _05137_);
  nand _63675_ (_12188_, _12187_, _03499_);
  and _63676_ (_12189_, _12188_, _12184_);
  and _63677_ (_12190_, _12189_, _12172_);
  nor _63678_ (_12191_, _05136_, _12173_);
  not _63679_ (_12192_, _05129_);
  and _63680_ (_12193_, _12192_, _05132_);
  and _63681_ (_12194_, _12193_, _12191_);
  and _63682_ (_12195_, _12194_, _03499_);
  and _63683_ (_12196_, _11468_, _03629_);
  nor _63684_ (_12197_, _11596_, _03629_);
  or _63685_ (_12198_, _12197_, _12196_);
  and _63686_ (_12199_, _12198_, _12195_);
  or _63687_ (_40634_, _12199_, _12190_);
  not _63688_ (_12200_, _12195_);
  or _63689_ (_12201_, _12183_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _63690_ (_12202_, _12201_, _12200_);
  nor _63691_ (_12203_, _06786_, _06547_);
  or _63692_ (_12204_, _12203_, _06785_);
  nor _63693_ (_12205_, _06765_, _05835_);
  nand _63694_ (_12206_, _12205_, _03972_);
  nor _63695_ (_12207_, _05617_, _04303_);
  and _63696_ (_12208_, _12207_, _04515_);
  or _63697_ (_12209_, _06764_, _04480_);
  nand _63698_ (_12210_, _08271_, _03745_);
  nor _63699_ (_12211_, _10095_, _05216_);
  or _63700_ (_12212_, _12211_, _05940_);
  nor _63701_ (_12213_, _05957_, _05667_);
  nor _63702_ (_12214_, _12213_, _06071_);
  nand _63703_ (_12215_, _12205_, _06073_);
  and _63704_ (_12216_, _03980_, _02878_);
  nor _63705_ (_12217_, _03980_, _03274_);
  or _63706_ (_12218_, _12217_, _12216_);
  nor _63707_ (_12219_, _12218_, _06073_);
  nor _63708_ (_12220_, _12219_, _04421_);
  and _63709_ (_12221_, _12220_, _12215_);
  or _63710_ (_12222_, _12221_, _04428_);
  or _63711_ (_12223_, _12222_, _12214_);
  nand _63712_ (_12224_, _10095_, _09695_);
  or _63713_ (_12225_, _12224_, _05954_);
  and _63714_ (_12226_, _12225_, _12223_);
  or _63715_ (_12227_, _12226_, _04768_);
  nor _63716_ (_12228_, _03230_, _02878_);
  nor _63717_ (_12229_, _12228_, _04431_);
  and _63718_ (_12230_, _12229_, _12227_);
  and _63719_ (_12231_, _06764_, _04431_);
  or _63720_ (_12232_, _12231_, _04449_);
  or _63721_ (_12233_, _12232_, _12230_);
  and _63722_ (_12234_, _12233_, _12212_);
  or _63723_ (_12235_, _12234_, _03508_);
  nand _63724_ (_12236_, _08271_, _03508_);
  and _63725_ (_12237_, _12236_, _04562_);
  and _63726_ (_12238_, _12237_, _12235_);
  not _63727_ (_12239_, _10096_);
  and _63728_ (_12240_, _12224_, _12239_);
  and _63729_ (_12241_, _12240_, _04454_);
  or _63730_ (_12242_, _12241_, _12238_);
  and _63731_ (_12243_, _12242_, _03227_);
  nor _63732_ (_12244_, _03227_, \oc8051_golden_model_1.PC [1]);
  or _63733_ (_12245_, _03745_, _12244_);
  or _63734_ (_12246_, _12245_, _12243_);
  and _63735_ (_12247_, _12246_, _12210_);
  or _63736_ (_12248_, _12247_, _04463_);
  and _63737_ (_12249_, _06501_, _03446_);
  nand _63738_ (_12250_, _08270_, _04463_);
  or _63739_ (_12251_, _12250_, _12249_);
  and _63740_ (_12252_, _12251_, _12248_);
  or _63741_ (_12253_, _12252_, _04462_);
  nor _63742_ (_12254_, _09718_, _05216_);
  and _63743_ (_12255_, _05216_, \oc8051_golden_model_1.PSW [7]);
  nor _63744_ (_12256_, _12255_, _12254_);
  nand _63745_ (_12257_, _12256_, _04462_);
  and _63746_ (_12258_, _12257_, _05897_);
  and _63747_ (_12259_, _12258_, _12253_);
  nand _63748_ (_12260_, _03224_, _02878_);
  nand _63749_ (_12261_, _04480_, _12260_);
  or _63750_ (_12262_, _12261_, _12259_);
  and _63751_ (_12263_, _12262_, _12209_);
  or _63752_ (_12264_, _12263_, _04482_);
  or _63753_ (_12265_, _06501_, _06164_);
  and _63754_ (_12266_, _12265_, _06163_);
  and _63755_ (_12267_, _12266_, _12264_);
  and _63756_ (_12268_, _05881_, _06764_);
  and _63757_ (_12269_, _06340_, \oc8051_golden_model_1.P1INREG [1]);
  not _63758_ (_12270_, _12269_);
  and _63759_ (_12271_, _06343_, \oc8051_golden_model_1.P0INREG [1]);
  not _63760_ (_12272_, _12271_);
  and _63761_ (_12273_, _06346_, \oc8051_golden_model_1.P2INREG [1]);
  and _63762_ (_12274_, _06348_, \oc8051_golden_model_1.P3INREG [1]);
  nor _63763_ (_12275_, _12274_, _12273_);
  and _63764_ (_12276_, _12275_, _12272_);
  and _63765_ (_12277_, _12276_, _12270_);
  and _63766_ (_12278_, _06354_, \oc8051_golden_model_1.SP [1]);
  and _63767_ (_12279_, _06284_, \oc8051_golden_model_1.TL0 [1]);
  nor _63768_ (_12280_, _12279_, _12278_);
  and _63769_ (_12281_, _12280_, _12277_);
  and _63770_ (_12282_, _06315_, \oc8051_golden_model_1.IE [1]);
  and _63771_ (_12283_, _06319_, \oc8051_golden_model_1.SBUF [1]);
  and _63772_ (_12284_, _06321_, \oc8051_golden_model_1.SCON [1]);
  or _63773_ (_12285_, _12284_, _12283_);
  nor _63774_ (_12286_, _12285_, _12282_);
  and _63775_ (_12287_, _06296_, \oc8051_golden_model_1.IP [1]);
  and _63776_ (_12288_, _06310_, \oc8051_golden_model_1.B [1]);
  nor _63777_ (_12289_, _12288_, _12287_);
  and _63778_ (_12290_, _06303_, \oc8051_golden_model_1.PSW [1]);
  and _63779_ (_12291_, _06308_, \oc8051_golden_model_1.ACC [1]);
  nor _63780_ (_12292_, _12291_, _12290_);
  and _63781_ (_12293_, _12292_, _12289_);
  and _63782_ (_12294_, _12293_, _12286_);
  and _63783_ (_12295_, _12294_, _12281_);
  and _63784_ (_12296_, _06327_, \oc8051_golden_model_1.TH0 [1]);
  and _63785_ (_12297_, _06329_, \oc8051_golden_model_1.TL1 [1]);
  nor _63786_ (_12298_, _12297_, _12296_);
  and _63787_ (_12299_, _06334_, \oc8051_golden_model_1.PCON [1]);
  and _63788_ (_12300_, _06336_, \oc8051_golden_model_1.TCON [1]);
  nor _63789_ (_12301_, _12300_, _12299_);
  and _63790_ (_12302_, _12301_, _12298_);
  and _63791_ (_12303_, _06272_, \oc8051_golden_model_1.DPH [1]);
  and _63792_ (_12304_, _06279_, \oc8051_golden_model_1.TMOD [1]);
  nor _63793_ (_12305_, _12304_, _12303_);
  and _63794_ (_12306_, _06356_, \oc8051_golden_model_1.DPL [1]);
  and _63795_ (_12307_, _06288_, \oc8051_golden_model_1.TH1 [1]);
  nor _63796_ (_12308_, _12307_, _12306_);
  and _63797_ (_12309_, _12308_, _12305_);
  and _63798_ (_12310_, _12309_, _12302_);
  and _63799_ (_12311_, _12310_, _12295_);
  not _63800_ (_12312_, _12311_);
  nor _63801_ (_12313_, _12312_, _12268_);
  nor _63802_ (_12314_, _12313_, _06170_);
  or _63803_ (_12315_, _12314_, _06168_);
  or _63804_ (_12316_, _12315_, _12267_);
  and _63805_ (_12317_, _06168_, _03414_);
  nor _63806_ (_12318_, _12317_, _04500_);
  and _63807_ (_12319_, _12318_, _12316_);
  and _63808_ (_12320_, _04500_, _06282_);
  or _63809_ (_12321_, _12320_, _03178_);
  or _63810_ (_12322_, _12321_, _12319_);
  and _63811_ (_12323_, _03178_, \oc8051_golden_model_1.PC [1]);
  nor _63812_ (_12324_, _12323_, _04512_);
  and _63813_ (_12325_, _12324_, _12322_);
  and _63814_ (_12326_, _05617_, _04303_);
  nor _63815_ (_12327_, _12326_, _12207_);
  nor _63816_ (_12328_, _12327_, _04511_);
  nor _63817_ (_12329_, _12328_, _04513_);
  or _63818_ (_12330_, _12329_, _12325_);
  nor _63819_ (_12331_, _05617_, _03274_);
  and _63820_ (_12332_, _05617_, _03274_);
  nor _63821_ (_12333_, _12332_, _12331_);
  or _63822_ (_12334_, _12333_, _05850_);
  and _63823_ (_12335_, _12334_, _06383_);
  and _63824_ (_12336_, _12335_, _12330_);
  or _63825_ (_12337_, _12336_, _12208_);
  and _63826_ (_12338_, _12337_, _06382_);
  and _63827_ (_12339_, _12331_, _04514_);
  or _63828_ (_12340_, _12339_, _03192_);
  or _63829_ (_12341_, _12340_, _12338_);
  and _63830_ (_12342_, _03192_, \oc8051_golden_model_1.PC [1]);
  nor _63831_ (_12343_, _12342_, _06390_);
  and _63832_ (_12344_, _12343_, _12341_);
  nor _63833_ (_12345_, _12326_, _06395_);
  or _63834_ (_12346_, _12345_, _06394_);
  or _63835_ (_12347_, _12346_, _12344_);
  nand _63836_ (_12348_, _12332_, _06394_);
  and _63837_ (_12349_, _12348_, _06399_);
  and _63838_ (_12350_, _12349_, _12347_);
  and _63839_ (_12351_, _03188_, _02878_);
  or _63840_ (_12352_, _03972_, _12351_);
  or _63841_ (_12353_, _12352_, _12350_);
  and _63842_ (_12354_, _12353_, _12206_);
  or _63843_ (_12355_, _12354_, _03491_);
  and _63844_ (_12356_, _12205_, _03491_);
  nor _63845_ (_12357_, _12356_, _04322_);
  and _63846_ (_12358_, _12357_, _12355_);
  nand _63847_ (_12359_, _12205_, _03027_);
  and _63848_ (_12360_, _12359_, _04803_);
  or _63849_ (_12361_, _12360_, _12358_);
  nand _63850_ (_12362_, _12205_, _03495_);
  and _63851_ (_12363_, _12362_, _06409_);
  and _63852_ (_12364_, _12363_, _12361_);
  nor _63853_ (_12365_, _12203_, _06409_);
  or _63854_ (_12366_, _12365_, _04531_);
  or _63855_ (_12367_, _12366_, _12364_);
  nand _63856_ (_12368_, _12213_, _04531_);
  and _63857_ (_12369_, _12368_, _12367_);
  or _63858_ (_12370_, _12369_, _03629_);
  not _63859_ (_12371_, _03198_);
  nand _63860_ (_12372_, _03629_, _11442_);
  and _63861_ (_12373_, _12372_, _12371_);
  and _63862_ (_12374_, _12373_, _12370_);
  and _63863_ (_12375_, _03198_, _02878_);
  or _63864_ (_12376_, _04539_, _12375_);
  or _63865_ (_12377_, _12376_, _12374_);
  or _63866_ (_12378_, _12254_, _04558_);
  and _63867_ (_12379_, _12378_, _11955_);
  and _63868_ (_12380_, _12379_, _12377_);
  and _63869_ (_12381_, _12205_, _11956_);
  or _63870_ (_12382_, _12381_, _04552_);
  or _63871_ (_12383_, _12382_, _12380_);
  and _63872_ (_12384_, _12383_, _12204_);
  or _63873_ (_12385_, _12384_, _03448_);
  or _63874_ (_12386_, _12213_, _04713_);
  and _63875_ (_12387_, _12386_, _04796_);
  and _63876_ (_12388_, _12387_, _12385_);
  or _63877_ (_12389_, _12388_, _11999_);
  and _63878_ (_12390_, _12389_, _12202_);
  nor _63879_ (_12391_, _11543_, _03629_);
  and _63880_ (_12392_, _11408_, _03629_);
  or _63881_ (_12393_, _12392_, _12391_);
  and _63882_ (_12394_, _12393_, _12195_);
  or _63883_ (_40635_, _12394_, _12390_);
  or _63884_ (_12395_, _12183_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _63885_ (_12396_, _12395_, _12200_);
  not _63886_ (_12397_, _12183_);
  nor _63887_ (_12398_, _06765_, _07849_);
  nor _63888_ (_12399_, _12398_, _07850_);
  and _63889_ (_12400_, _12399_, _11956_);
  not _63890_ (_12401_, _06637_);
  and _63891_ (_12402_, _06547_, _12401_);
  nor _63892_ (_12403_, _06547_, _12401_);
  or _63893_ (_12404_, _12403_, _12402_);
  and _63894_ (_12405_, _12404_, _04242_);
  and _63895_ (_12406_, _03210_, _03188_);
  nor _63896_ (_12407_, _05717_, _03946_);
  and _63897_ (_12408_, _12407_, _04515_);
  nor _63898_ (_12409_, _10083_, _05302_);
  or _63899_ (_12410_, _12409_, _05940_);
  nand _63900_ (_12411_, _10083_, _09670_);
  or _63901_ (_12412_, _12411_, _05954_);
  and _63902_ (_12413_, _05717_, _05617_);
  and _63903_ (_12414_, _12413_, _05956_);
  nor _63904_ (_12415_, _05957_, _05717_);
  nor _63905_ (_12416_, _12415_, _12414_);
  nor _63906_ (_12417_, _12416_, _06071_);
  and _63907_ (_12418_, _05835_, _04875_);
  nor _63908_ (_12419_, _05835_, _04875_);
  or _63909_ (_12420_, _12419_, _12418_);
  or _63910_ (_12421_, _12420_, _06072_);
  and _63911_ (_12422_, _03980_, _03210_);
  nor _63912_ (_12423_, _03980_, _07584_);
  or _63913_ (_12424_, _12423_, _12422_);
  nor _63914_ (_12425_, _12424_, _06073_);
  nor _63915_ (_12426_, _12425_, _04421_);
  and _63916_ (_12427_, _12426_, _12421_);
  or _63917_ (_12428_, _12427_, _04428_);
  or _63918_ (_12429_, _12428_, _12417_);
  and _63919_ (_12430_, _12429_, _12412_);
  or _63920_ (_12431_, _12430_, _04768_);
  nor _63921_ (_12432_, _03210_, _03230_);
  nor _63922_ (_12433_, _12432_, _04431_);
  and _63923_ (_12434_, _12433_, _12431_);
  and _63924_ (_12435_, _07849_, _04431_);
  or _63925_ (_12436_, _12435_, _04449_);
  or _63926_ (_12437_, _12436_, _12434_);
  and _63927_ (_12438_, _12437_, _12410_);
  or _63928_ (_12439_, _12438_, _03508_);
  nand _63929_ (_12440_, _08260_, _03508_);
  and _63930_ (_12441_, _12440_, _04562_);
  and _63931_ (_12442_, _12441_, _12439_);
  not _63932_ (_12443_, _10084_);
  and _63933_ (_12444_, _12411_, _12443_);
  and _63934_ (_12445_, _12444_, _04454_);
  or _63935_ (_12446_, _12445_, _12442_);
  and _63936_ (_12447_, _12446_, _03227_);
  nor _63937_ (_12448_, _03245_, _03227_);
  or _63938_ (_12449_, _03745_, _12448_);
  or _63939_ (_12450_, _12449_, _12447_);
  nand _63940_ (_12451_, _08260_, _03745_);
  and _63941_ (_12452_, _12451_, _12450_);
  or _63942_ (_12453_, _12452_, _04463_);
  and _63943_ (_12454_, _06637_, _03446_);
  nand _63944_ (_12455_, _08259_, _04463_);
  or _63945_ (_12456_, _12455_, _12454_);
  and _63946_ (_12457_, _12456_, _12453_);
  or _63947_ (_12458_, _12457_, _04462_);
  nor _63948_ (_12459_, _09693_, _05302_);
  and _63949_ (_12460_, _05302_, \oc8051_golden_model_1.PSW [7]);
  nor _63950_ (_12461_, _12460_, _12459_);
  nand _63951_ (_12462_, _12461_, _04462_);
  and _63952_ (_12463_, _12462_, _05897_);
  and _63953_ (_12464_, _12463_, _12458_);
  nand _63954_ (_12465_, _03210_, _03224_);
  nand _63955_ (_12466_, _04480_, _12465_);
  or _63956_ (_12467_, _12466_, _12464_);
  or _63957_ (_12468_, _07849_, _04480_);
  and _63958_ (_12469_, _12468_, _12467_);
  or _63959_ (_12470_, _12469_, _04482_);
  or _63960_ (_12471_, _06637_, _06164_);
  and _63961_ (_12472_, _12471_, _06163_);
  and _63962_ (_12473_, _12472_, _12470_);
  nor _63963_ (_12474_, _06171_, _04875_);
  and _63964_ (_12475_, _06340_, \oc8051_golden_model_1.P1INREG [2]);
  not _63965_ (_12476_, _12475_);
  and _63966_ (_12477_, _06343_, \oc8051_golden_model_1.P0INREG [2]);
  not _63967_ (_12478_, _12477_);
  and _63968_ (_12479_, _06346_, \oc8051_golden_model_1.P2INREG [2]);
  and _63969_ (_12480_, _06348_, \oc8051_golden_model_1.P3INREG [2]);
  nor _63970_ (_12481_, _12480_, _12479_);
  and _63971_ (_12482_, _12481_, _12478_);
  and _63972_ (_12483_, _12482_, _12476_);
  and _63973_ (_12484_, _06284_, \oc8051_golden_model_1.TL0 [2]);
  and _63974_ (_12485_, _06279_, \oc8051_golden_model_1.TMOD [2]);
  nor _63975_ (_12486_, _12485_, _12484_);
  and _63976_ (_12487_, _12486_, _12483_);
  and _63977_ (_12488_, _06315_, \oc8051_golden_model_1.IE [2]);
  and _63978_ (_12489_, _06319_, \oc8051_golden_model_1.SBUF [2]);
  and _63979_ (_12490_, _06321_, \oc8051_golden_model_1.SCON [2]);
  or _63980_ (_12491_, _12490_, _12489_);
  nor _63981_ (_12492_, _12491_, _12488_);
  and _63982_ (_12493_, _06272_, \oc8051_golden_model_1.DPH [2]);
  and _63983_ (_12494_, _06288_, \oc8051_golden_model_1.TH1 [2]);
  nor _63984_ (_12495_, _12494_, _12493_);
  and _63985_ (_12496_, _12495_, _12492_);
  and _63986_ (_12497_, _12496_, _12487_);
  and _63987_ (_12498_, _06327_, \oc8051_golden_model_1.TH0 [2]);
  and _63988_ (_12499_, _06329_, \oc8051_golden_model_1.TL1 [2]);
  nor _63989_ (_12500_, _12499_, _12498_);
  and _63990_ (_12501_, _06334_, \oc8051_golden_model_1.PCON [2]);
  and _63991_ (_12502_, _06336_, \oc8051_golden_model_1.TCON [2]);
  nor _63992_ (_12503_, _12502_, _12501_);
  and _63993_ (_12504_, _12503_, _12500_);
  and _63994_ (_12505_, _06296_, \oc8051_golden_model_1.IP [2]);
  and _63995_ (_12506_, _06303_, \oc8051_golden_model_1.PSW [2]);
  nor _63996_ (_12507_, _12506_, _12505_);
  and _63997_ (_12508_, _06308_, \oc8051_golden_model_1.ACC [2]);
  and _63998_ (_12509_, _06310_, \oc8051_golden_model_1.B [2]);
  nor _63999_ (_12510_, _12509_, _12508_);
  and _64000_ (_12511_, _12510_, _12507_);
  and _64001_ (_12512_, _06354_, \oc8051_golden_model_1.SP [2]);
  and _64002_ (_12513_, _06356_, \oc8051_golden_model_1.DPL [2]);
  nor _64003_ (_12514_, _12513_, _12512_);
  and _64004_ (_12515_, _12514_, _12511_);
  and _64005_ (_12516_, _12515_, _12504_);
  and _64006_ (_12517_, _12516_, _12497_);
  not _64007_ (_12518_, _12517_);
  nor _64008_ (_12519_, _12518_, _12474_);
  nor _64009_ (_12520_, _12519_, _06170_);
  or _64010_ (_12521_, _12520_, _06168_);
  or _64011_ (_12522_, _12521_, _12473_);
  and _64012_ (_12523_, _06168_, _03904_);
  nor _64013_ (_12524_, _12523_, _04500_);
  and _64014_ (_12525_, _12524_, _12522_);
  and _64015_ (_12526_, _04500_, _06332_);
  or _64016_ (_12527_, _12526_, _03178_);
  or _64017_ (_12528_, _12527_, _12525_);
  and _64018_ (_12529_, _03245_, _03178_);
  nor _64019_ (_12530_, _12529_, _04512_);
  and _64020_ (_12531_, _12530_, _12528_);
  and _64021_ (_12532_, _05717_, _03946_);
  nor _64022_ (_12533_, _12532_, _12407_);
  nor _64023_ (_12534_, _12533_, _04511_);
  nor _64024_ (_12535_, _12534_, _04513_);
  or _64025_ (_12536_, _12535_, _12531_);
  nor _64026_ (_12537_, _05717_, _07584_);
  and _64027_ (_12538_, _05717_, _07584_);
  nor _64028_ (_12539_, _12538_, _12537_);
  or _64029_ (_12540_, _12539_, _05850_);
  and _64030_ (_12541_, _12540_, _06383_);
  and _64031_ (_12542_, _12541_, _12536_);
  or _64032_ (_12543_, _12542_, _12408_);
  and _64033_ (_12544_, _12543_, _06382_);
  and _64034_ (_12545_, _12537_, _04514_);
  or _64035_ (_12546_, _12545_, _03192_);
  or _64036_ (_12547_, _12546_, _12544_);
  and _64037_ (_12548_, _03245_, _03192_);
  nor _64038_ (_12549_, _12548_, _06390_);
  and _64039_ (_12550_, _12549_, _12547_);
  nor _64040_ (_12551_, _12532_, _06395_);
  or _64041_ (_12552_, _12551_, _06394_);
  or _64042_ (_12553_, _12552_, _12550_);
  nand _64043_ (_12554_, _12538_, _06394_);
  and _64044_ (_12555_, _12554_, _06399_);
  and _64045_ (_12556_, _12555_, _12553_);
  or _64046_ (_12557_, _12556_, _12406_);
  and _64047_ (_12558_, _12557_, _05848_);
  not _64048_ (_12559_, _02994_);
  and _64049_ (_12560_, _04533_, _12559_);
  not _64050_ (_12561_, _05848_);
  and _64051_ (_12562_, _12420_, _12561_);
  or _64052_ (_12563_, _12562_, _12560_);
  or _64053_ (_12564_, _12563_, _12558_);
  not _64054_ (_12565_, _04242_);
  nand _64055_ (_12566_, _04533_, _12559_);
  or _64056_ (_12567_, _12566_, _12404_);
  and _64057_ (_12568_, _12567_, _12565_);
  and _64058_ (_12569_, _12568_, _12564_);
  or _64059_ (_12570_, _12569_, _12405_);
  and _64060_ (_12571_, _12570_, _06408_);
  nor _64061_ (_12572_, _12416_, _06408_);
  or _64062_ (_12573_, _12572_, _03629_);
  or _64063_ (_12574_, _12573_, _12571_);
  nand _64064_ (_12575_, _11440_, _03629_);
  and _64065_ (_12576_, _12575_, _12371_);
  and _64066_ (_12577_, _12576_, _12574_);
  and _64067_ (_12578_, _03210_, _03198_);
  or _64068_ (_12579_, _04539_, _12578_);
  or _64069_ (_12580_, _12579_, _12577_);
  or _64070_ (_12581_, _12459_, _04558_);
  and _64071_ (_12582_, _12581_, _11955_);
  and _64072_ (_12583_, _12582_, _12580_);
  or _64073_ (_12584_, _12583_, _12400_);
  and _64074_ (_12585_, _12584_, _06785_);
  or _64075_ (_12586_, _06786_, _06637_);
  nor _64076_ (_12587_, _08016_, _06785_);
  and _64077_ (_12588_, _12587_, _12586_);
  or _64078_ (_12589_, _12588_, _03448_);
  or _64079_ (_12590_, _12589_, _12585_);
  nor _64080_ (_12591_, _05718_, _05667_);
  nor _64081_ (_12592_, _12591_, _05719_);
  or _64082_ (_12593_, _12592_, _04713_);
  and _64083_ (_12594_, _12593_, _12174_);
  and _64084_ (_12595_, _12594_, _12590_);
  or _64085_ (_12596_, _12595_, _12397_);
  and _64086_ (_12597_, _12596_, _12396_);
  and _64087_ (_12598_, _11394_, _03629_);
  and _64088_ (_12599_, _11529_, _11944_);
  or _64089_ (_12600_, _12599_, _12598_);
  and _64090_ (_12601_, _12600_, _12195_);
  or _64091_ (_40637_, _12601_, _12597_);
  or _64092_ (_12602_, _12183_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _64093_ (_12603_, _12602_, _12200_);
  nor _64094_ (_12604_, _12402_, _08636_);
  or _64095_ (_12605_, _12604_, _06639_);
  and _64096_ (_12606_, _12605_, _04533_);
  and _64097_ (_12607_, _03297_, _03188_);
  nor _64098_ (_12608_, _05566_, _03708_);
  and _64099_ (_12609_, _12608_, _04515_);
  and _64100_ (_12610_, _05296_, \oc8051_golden_model_1.PSW [7]);
  nor _64101_ (_12611_, _09825_, _05296_);
  nor _64102_ (_12612_, _12611_, _12610_);
  nor _64103_ (_12613_, _12612_, _05063_);
  or _64104_ (_12614_, _08636_, _03454_);
  nand _64105_ (_12615_, _12614_, _08247_);
  and _64106_ (_12616_, _12615_, _04463_);
  nor _64107_ (_12617_, _12418_, _05005_);
  or _64108_ (_12618_, _12617_, _05837_);
  or _64109_ (_12619_, _12618_, _06072_);
  and _64110_ (_12620_, _03980_, _03297_);
  nor _64111_ (_12621_, _03980_, _07578_);
  or _64112_ (_12622_, _12621_, _06073_);
  or _64113_ (_12623_, _12622_, _12620_);
  and _64114_ (_12624_, _12623_, _12619_);
  and _64115_ (_12625_, _12624_, _06071_);
  nor _64116_ (_12626_, _12414_, _05566_);
  nor _64117_ (_12627_, _12626_, _05959_);
  nor _64118_ (_12628_, _12627_, _06071_);
  or _64119_ (_12629_, _12628_, _12625_);
  or _64120_ (_12630_, _12629_, _04428_);
  nand _64121_ (_12631_, _10146_, _09802_);
  or _64122_ (_12632_, _12631_, _05954_);
  and _64123_ (_12633_, _12632_, _12630_);
  or _64124_ (_12634_, _12633_, _04768_);
  nor _64125_ (_12635_, _03297_, _03230_);
  nor _64126_ (_12636_, _12635_, _04431_);
  and _64127_ (_12637_, _12636_, _12634_);
  and _64128_ (_12638_, _07848_, _04431_);
  or _64129_ (_12639_, _12638_, _04449_);
  or _64130_ (_12640_, _12639_, _12637_);
  nor _64131_ (_12641_, _10146_, _05296_);
  or _64132_ (_12642_, _12641_, _05940_);
  and _64133_ (_12643_, _12642_, _12640_);
  or _64134_ (_12644_, _12643_, _03508_);
  nand _64135_ (_12645_, _08248_, _03508_);
  and _64136_ (_12646_, _12645_, _04562_);
  and _64137_ (_12647_, _12646_, _12644_);
  not _64138_ (_12648_, _10147_);
  and _64139_ (_12649_, _12631_, _12648_);
  and _64140_ (_12650_, _12649_, _04454_);
  or _64141_ (_12651_, _12650_, _12647_);
  and _64142_ (_12652_, _12651_, _03227_);
  nor _64143_ (_12653_, _03648_, _03227_);
  or _64144_ (_12654_, _03745_, _12653_);
  or _64145_ (_12655_, _12654_, _12652_);
  nand _64146_ (_12656_, _08248_, _03745_);
  and _64147_ (_12657_, _12656_, _05976_);
  and _64148_ (_12658_, _12657_, _12655_);
  or _64149_ (_12659_, _12658_, _12616_);
  and _64150_ (_12660_, _12659_, _05063_);
  or _64151_ (_12661_, _12660_, _12613_);
  and _64152_ (_12662_, _12661_, _05897_);
  nand _64153_ (_12663_, _03297_, _03224_);
  nand _64154_ (_12664_, _04480_, _12663_);
  or _64155_ (_12665_, _12664_, _12662_);
  or _64156_ (_12666_, _07848_, _04480_);
  and _64157_ (_12667_, _12666_, _12665_);
  or _64158_ (_12668_, _12667_, _04482_);
  or _64159_ (_12669_, _06592_, _06164_);
  and _64160_ (_12670_, _12669_, _06163_);
  and _64161_ (_12671_, _12670_, _12668_);
  nor _64162_ (_12672_, _06171_, _05005_);
  and _64163_ (_12673_, _06356_, \oc8051_golden_model_1.DPL [3]);
  and _64164_ (_12674_, _06284_, \oc8051_golden_model_1.TL0 [3]);
  nor _64165_ (_12675_, _12674_, _12673_);
  and _64166_ (_12676_, _06272_, \oc8051_golden_model_1.DPH [3]);
  and _64167_ (_12677_, _06288_, \oc8051_golden_model_1.TH1 [3]);
  nor _64168_ (_12678_, _12677_, _12676_);
  and _64169_ (_12679_, _12678_, _12675_);
  and _64170_ (_12680_, _06315_, \oc8051_golden_model_1.IE [3]);
  and _64171_ (_12681_, _06319_, \oc8051_golden_model_1.SBUF [3]);
  and _64172_ (_12682_, _06321_, \oc8051_golden_model_1.SCON [3]);
  or _64173_ (_12683_, _12682_, _12681_);
  nor _64174_ (_12684_, _12683_, _12680_);
  and _64175_ (_12685_, _06296_, \oc8051_golden_model_1.IP [3]);
  and _64176_ (_12686_, _06303_, \oc8051_golden_model_1.PSW [3]);
  nor _64177_ (_12687_, _12686_, _12685_);
  and _64178_ (_12688_, _06308_, \oc8051_golden_model_1.ACC [3]);
  and _64179_ (_12689_, _06310_, \oc8051_golden_model_1.B [3]);
  nor _64180_ (_12690_, _12689_, _12688_);
  and _64181_ (_12691_, _12690_, _12687_);
  and _64182_ (_12692_, _12691_, _12684_);
  and _64183_ (_12693_, _12692_, _12679_);
  and _64184_ (_12694_, _06327_, \oc8051_golden_model_1.TH0 [3]);
  and _64185_ (_12695_, _06329_, \oc8051_golden_model_1.TL1 [3]);
  nor _64186_ (_12696_, _12695_, _12694_);
  and _64187_ (_12697_, _06334_, \oc8051_golden_model_1.PCON [3]);
  and _64188_ (_12698_, _06336_, \oc8051_golden_model_1.TCON [3]);
  nor _64189_ (_12699_, _12698_, _12697_);
  and _64190_ (_12700_, _12699_, _12696_);
  and _64191_ (_12701_, _06340_, \oc8051_golden_model_1.P1INREG [3]);
  not _64192_ (_12703_, _12701_);
  and _64193_ (_12704_, _06343_, \oc8051_golden_model_1.P0INREG [3]);
  not _64194_ (_12705_, _12704_);
  and _64195_ (_12706_, _06346_, \oc8051_golden_model_1.P2INREG [3]);
  and _64196_ (_12707_, _06348_, \oc8051_golden_model_1.P3INREG [3]);
  nor _64197_ (_12708_, _12707_, _12706_);
  and _64198_ (_12709_, _12708_, _12705_);
  and _64199_ (_12710_, _12709_, _12703_);
  and _64200_ (_12711_, _06354_, \oc8051_golden_model_1.SP [3]);
  and _64201_ (_12712_, _06279_, \oc8051_golden_model_1.TMOD [3]);
  nor _64202_ (_12713_, _12712_, _12711_);
  and _64203_ (_12714_, _12713_, _12710_);
  and _64204_ (_12715_, _12714_, _12700_);
  and _64205_ (_12716_, _12715_, _12693_);
  not _64206_ (_12717_, _12716_);
  nor _64207_ (_12718_, _12717_, _12672_);
  nor _64208_ (_12719_, _12718_, _06170_);
  or _64209_ (_12720_, _12719_, _06168_);
  or _64210_ (_12721_, _12720_, _12671_);
  and _64211_ (_12722_, _06168_, _03581_);
  nor _64212_ (_12724_, _12722_, _04500_);
  and _64213_ (_12725_, _12724_, _12721_);
  and _64214_ (_12726_, _04500_, _06276_);
  or _64215_ (_12727_, _12726_, _03178_);
  or _64216_ (_12728_, _12727_, _12725_);
  and _64217_ (_12729_, _03648_, _03178_);
  nor _64218_ (_12730_, _12729_, _04512_);
  and _64219_ (_12731_, _12730_, _12728_);
  and _64220_ (_12732_, _05566_, _03708_);
  nor _64221_ (_12733_, _12732_, _12608_);
  nor _64222_ (_12734_, _12733_, _04511_);
  nor _64223_ (_12735_, _12734_, _04513_);
  or _64224_ (_12736_, _12735_, _12731_);
  nor _64225_ (_12737_, _05566_, _07578_);
  and _64226_ (_12738_, _05566_, _07578_);
  nor _64227_ (_12739_, _12738_, _12737_);
  or _64228_ (_12740_, _12739_, _05850_);
  and _64229_ (_12741_, _12740_, _06383_);
  and _64230_ (_12742_, _12741_, _12736_);
  or _64231_ (_12743_, _12742_, _12609_);
  and _64232_ (_12744_, _12743_, _06382_);
  and _64233_ (_12745_, _12737_, _04514_);
  or _64234_ (_12746_, _12745_, _03192_);
  or _64235_ (_12747_, _12746_, _12744_);
  and _64236_ (_12748_, _03648_, _03192_);
  nor _64237_ (_12749_, _12748_, _06390_);
  and _64238_ (_12750_, _12749_, _12747_);
  nor _64239_ (_12751_, _12732_, _06395_);
  or _64240_ (_12752_, _12751_, _06394_);
  or _64241_ (_12753_, _12752_, _12750_);
  nand _64242_ (_12754_, _12738_, _06394_);
  and _64243_ (_12755_, _12754_, _06399_);
  and _64244_ (_12756_, _12755_, _12753_);
  or _64245_ (_12757_, _12756_, _12607_);
  and _64246_ (_12758_, _12757_, _05847_);
  not _64247_ (_12759_, _05847_);
  and _64248_ (_12760_, _12618_, _12759_);
  or _64249_ (_12761_, _12760_, _03495_);
  or _64250_ (_12762_, _12761_, _12758_);
  or _64251_ (_12763_, _12618_, _04745_);
  and _64252_ (_12764_, _12763_, _06409_);
  and _64253_ (_12765_, _12764_, _12762_);
  or _64254_ (_12766_, _12765_, _12606_);
  and _64255_ (_12767_, _12766_, _06408_);
  nor _64256_ (_12768_, _12627_, _06408_);
  or _64257_ (_12769_, _12768_, _03629_);
  or _64258_ (_12770_, _12769_, _12767_);
  nand _64259_ (_12771_, _11435_, _03629_);
  and _64260_ (_12772_, _12771_, _12371_);
  and _64261_ (_12773_, _12772_, _12770_);
  and _64262_ (_12774_, _03297_, _03198_);
  or _64263_ (_12775_, _04539_, _12774_);
  or _64264_ (_12776_, _12775_, _12773_);
  or _64265_ (_12777_, _12611_, _04558_);
  and _64266_ (_12778_, _12777_, _06757_);
  and _64267_ (_12779_, _12778_, _12776_);
  nor _64268_ (_12780_, _07850_, _07848_);
  nor _64269_ (_12781_, _12780_, _06767_);
  and _64270_ (_12782_, _12781_, _06758_);
  or _64271_ (_12783_, _12782_, _04547_);
  or _64272_ (_12784_, _12783_, _12779_);
  or _64273_ (_12785_, _12781_, _06780_);
  and _64274_ (_12786_, _12785_, _06785_);
  and _64275_ (_12787_, _12786_, _12784_);
  or _64276_ (_12788_, _08016_, _06592_);
  nor _64277_ (_12789_, _06788_, _06785_);
  and _64278_ (_12790_, _12789_, _12788_);
  or _64279_ (_12791_, _12790_, _03448_);
  or _64280_ (_12792_, _12791_, _12787_);
  nor _64281_ (_12793_, _05719_, _05567_);
  nor _64282_ (_12794_, _12793_, _05720_);
  or _64283_ (_12795_, _12794_, _04713_);
  and _64284_ (_12796_, _12795_, _12174_);
  and _64285_ (_12797_, _12796_, _12792_);
  or _64286_ (_12798_, _12797_, _12397_);
  and _64287_ (_12799_, _12798_, _12603_);
  nor _64288_ (_12800_, _11534_, _03629_);
  and _64289_ (_12801_, _11399_, _03629_);
  or _64290_ (_12802_, _12801_, _12800_);
  and _64291_ (_12803_, _12802_, _12195_);
  or _64292_ (_40638_, _12803_, _12799_);
  or _64293_ (_12804_, _12183_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _64294_ (_12805_, _12804_, _12200_);
  not _64295_ (_12806_, _06730_);
  and _64296_ (_12807_, _06639_, _12806_);
  nor _64297_ (_12808_, _06639_, _12806_);
  or _64298_ (_12809_, _12808_, _12807_);
  and _64299_ (_12810_, _12809_, _04533_);
  nor _64300_ (_12811_, _05837_, _05777_);
  and _64301_ (_12812_, _05837_, _05777_);
  or _64302_ (_12813_, _12812_, _12811_);
  or _64303_ (_12814_, _12813_, _05847_);
  nor _64304_ (_12815_, _05824_, _07484_);
  and _64305_ (_12816_, _05824_, _07484_);
  nor _64306_ (_12817_, _12816_, _12815_);
  and _64307_ (_12818_, _12817_, _04511_);
  and _64308_ (_12819_, _06236_, _05824_);
  nor _64309_ (_12820_, _06236_, _05824_);
  nor _64310_ (_12821_, _12820_, _12819_);
  and _64311_ (_12822_, _12821_, _04512_);
  nor _64312_ (_12823_, _09745_, _09721_);
  and _64313_ (_12824_, _09721_, \oc8051_golden_model_1.PSW [7]);
  nor _64314_ (_12825_, _12824_, _12823_);
  nor _64315_ (_12826_, _12825_, _05063_);
  nor _64316_ (_12827_, _09721_, _10109_);
  or _64317_ (_12828_, _12827_, _05940_);
  and _64318_ (_12829_, _11564_, _03980_);
  nor _64319_ (_12830_, _03980_, _07484_);
  or _64320_ (_12831_, _12830_, _12829_);
  and _64321_ (_12832_, _12831_, _06072_);
  and _64322_ (_12833_, _12813_, _06073_);
  or _64323_ (_12834_, _12833_, _12832_);
  and _64324_ (_12835_, _12834_, _05966_);
  and _64325_ (_12836_, _06730_, _04422_);
  or _64326_ (_12837_, _12836_, _12835_);
  and _64327_ (_12838_, _12837_, _06071_);
  and _64328_ (_12839_, _05959_, _05824_);
  nor _64329_ (_12840_, _05959_, _05824_);
  nor _64330_ (_12841_, _12840_, _12839_);
  nor _64331_ (_12842_, _12841_, _06071_);
  or _64332_ (_12843_, _12842_, _12838_);
  and _64333_ (_12844_, _12843_, _05954_);
  nand _64334_ (_12845_, _09722_, _10109_);
  and _64335_ (_12846_, _12845_, _04428_);
  or _64336_ (_12847_, _12846_, _04768_);
  or _64337_ (_12848_, _12847_, _12844_);
  nor _64338_ (_12849_, _11564_, _03230_);
  nor _64339_ (_12850_, _12849_, _04431_);
  and _64340_ (_12851_, _12850_, _12848_);
  and _64341_ (_12852_, _06763_, _04431_);
  or _64342_ (_12853_, _12852_, _04449_);
  or _64343_ (_12854_, _12853_, _12851_);
  and _64344_ (_12855_, _12854_, _12828_);
  or _64345_ (_12856_, _12855_, _03508_);
  nand _64346_ (_12857_, _08235_, _03508_);
  and _64347_ (_12858_, _12857_, _04562_);
  and _64348_ (_12859_, _12858_, _12856_);
  not _64349_ (_12860_, _10110_);
  and _64350_ (_12861_, _12845_, _12860_);
  and _64351_ (_12862_, _12861_, _04454_);
  or _64352_ (_12863_, _12862_, _12859_);
  and _64353_ (_12864_, _12863_, _03227_);
  nor _64354_ (_12865_, _11565_, _03227_);
  or _64355_ (_12866_, _12865_, _03745_);
  or _64356_ (_12867_, _12866_, _12864_);
  nand _64357_ (_12868_, _08235_, _03745_);
  and _64358_ (_12869_, _12868_, _12867_);
  or _64359_ (_12870_, _12869_, _04463_);
  and _64360_ (_12871_, _06730_, _03446_);
  nand _64361_ (_12872_, _08234_, _04463_);
  or _64362_ (_12873_, _12872_, _12871_);
  and _64363_ (_12874_, _12873_, _05063_);
  and _64364_ (_12875_, _12874_, _12870_);
  or _64365_ (_12876_, _12875_, _12826_);
  and _64366_ (_12877_, _12876_, _05897_);
  nand _64367_ (_12878_, _11564_, _03224_);
  nand _64368_ (_12879_, _12878_, _04480_);
  or _64369_ (_12880_, _12879_, _12877_);
  or _64370_ (_12881_, _06763_, _04480_);
  and _64371_ (_12882_, _12881_, _12880_);
  or _64372_ (_12883_, _12882_, _04482_);
  or _64373_ (_12884_, _06730_, _06164_);
  and _64374_ (_12885_, _12884_, _06163_);
  and _64375_ (_12886_, _12885_, _12883_);
  nor _64376_ (_12887_, _06171_, _05777_);
  and _64377_ (_12888_, _06340_, \oc8051_golden_model_1.P1INREG [4]);
  not _64378_ (_12889_, _12888_);
  and _64379_ (_12890_, _06343_, \oc8051_golden_model_1.P0INREG [4]);
  not _64380_ (_12891_, _12890_);
  and _64381_ (_12892_, _06346_, \oc8051_golden_model_1.P2INREG [4]);
  and _64382_ (_12893_, _06348_, \oc8051_golden_model_1.P3INREG [4]);
  nor _64383_ (_12894_, _12893_, _12892_);
  and _64384_ (_12895_, _12894_, _12891_);
  and _64385_ (_12896_, _12895_, _12889_);
  and _64386_ (_12897_, _06354_, \oc8051_golden_model_1.SP [4]);
  and _64387_ (_12898_, _06284_, \oc8051_golden_model_1.TL0 [4]);
  nor _64388_ (_12899_, _12898_, _12897_);
  and _64389_ (_12900_, _12899_, _12896_);
  and _64390_ (_12901_, _06315_, \oc8051_golden_model_1.IE [4]);
  and _64391_ (_12902_, _06319_, \oc8051_golden_model_1.SBUF [4]);
  and _64392_ (_12903_, _06321_, \oc8051_golden_model_1.SCON [4]);
  or _64393_ (_12904_, _12903_, _12902_);
  nor _64394_ (_12905_, _12904_, _12901_);
  and _64395_ (_12906_, _06296_, \oc8051_golden_model_1.IP [4]);
  and _64396_ (_12907_, _06310_, \oc8051_golden_model_1.B [4]);
  nor _64397_ (_12908_, _12907_, _12906_);
  and _64398_ (_12909_, _06303_, \oc8051_golden_model_1.PSW [4]);
  and _64399_ (_12910_, _06308_, \oc8051_golden_model_1.ACC [4]);
  nor _64400_ (_12911_, _12910_, _12909_);
  and _64401_ (_12912_, _12911_, _12908_);
  and _64402_ (_12913_, _12912_, _12905_);
  and _64403_ (_12914_, _12913_, _12900_);
  and _64404_ (_12915_, _06272_, \oc8051_golden_model_1.DPH [4]);
  and _64405_ (_12916_, _06279_, \oc8051_golden_model_1.TMOD [4]);
  nor _64406_ (_12917_, _12916_, _12915_);
  and _64407_ (_12918_, _06356_, \oc8051_golden_model_1.DPL [4]);
  and _64408_ (_12919_, _06288_, \oc8051_golden_model_1.TH1 [4]);
  nor _64409_ (_12920_, _12919_, _12918_);
  and _64410_ (_12921_, _12920_, _12917_);
  and _64411_ (_12922_, _06293_, _06269_);
  and _64412_ (_12923_, _12922_, \oc8051_golden_model_1.TCON [4]);
  and _64413_ (_12924_, _06327_, \oc8051_golden_model_1.TH0 [4]);
  nor _64414_ (_12925_, _12924_, _12923_);
  and _64415_ (_12926_, _06334_, \oc8051_golden_model_1.PCON [4]);
  and _64416_ (_12927_, _06329_, \oc8051_golden_model_1.TL1 [4]);
  nor _64417_ (_12928_, _12927_, _12926_);
  and _64418_ (_12929_, _12928_, _12925_);
  and _64419_ (_12930_, _12929_, _12921_);
  and _64420_ (_12931_, _12930_, _12914_);
  not _64421_ (_12932_, _12931_);
  nor _64422_ (_12933_, _12932_, _12887_);
  nor _64423_ (_12934_, _12933_, _06170_);
  or _64424_ (_12935_, _12934_, _06168_);
  or _64425_ (_12936_, _12935_, _12886_);
  and _64426_ (_12937_, _06168_, _03486_);
  nor _64427_ (_12938_, _12937_, _04500_);
  and _64428_ (_12939_, _12938_, _12936_);
  and _64429_ (_12940_, _06298_, _04500_);
  or _64430_ (_12941_, _12940_, _03178_);
  or _64431_ (_12942_, _12941_, _12939_);
  and _64432_ (_12943_, _11565_, _03178_);
  nor _64433_ (_12944_, _12943_, _04512_);
  and _64434_ (_12945_, _12944_, _12942_);
  or _64435_ (_12946_, _12945_, _12822_);
  and _64436_ (_12947_, _12946_, _05850_);
  or _64437_ (_12948_, _12947_, _12818_);
  and _64438_ (_12949_, _12948_, _06383_);
  and _64439_ (_12950_, _12820_, _04515_);
  or _64440_ (_12951_, _12950_, _12949_);
  and _64441_ (_12952_, _12951_, _06382_);
  and _64442_ (_12953_, _12815_, _04514_);
  or _64443_ (_12954_, _12953_, _03192_);
  or _64444_ (_12955_, _12954_, _12952_);
  and _64445_ (_12956_, _11565_, _03192_);
  nor _64446_ (_12957_, _12956_, _06390_);
  and _64447_ (_12958_, _12957_, _12955_);
  nor _64448_ (_12959_, _12819_, _06395_);
  or _64449_ (_12960_, _12959_, _06394_);
  or _64450_ (_12961_, _12960_, _12958_);
  nand _64451_ (_12962_, _12816_, _06394_);
  and _64452_ (_12963_, _12962_, _06399_);
  and _64453_ (_12964_, _12963_, _12961_);
  nand _64454_ (_12965_, _11564_, _03188_);
  nand _64455_ (_12966_, _12965_, _05847_);
  or _64456_ (_12967_, _12966_, _12964_);
  and _64457_ (_12968_, _12967_, _12814_);
  or _64458_ (_12969_, _12968_, _03495_);
  or _64459_ (_12970_, _12813_, _04745_);
  and _64460_ (_12971_, _12970_, _06409_);
  and _64461_ (_12972_, _12971_, _12969_);
  or _64462_ (_12973_, _12972_, _12810_);
  and _64463_ (_12974_, _12973_, _06408_);
  nor _64464_ (_12975_, _12841_, _06408_);
  or _64465_ (_12976_, _12975_, _03629_);
  or _64466_ (_12977_, _12976_, _12974_);
  nand _64467_ (_12978_, _11431_, _03629_);
  and _64468_ (_12979_, _12978_, _12371_);
  and _64469_ (_12980_, _12979_, _12977_);
  and _64470_ (_12981_, _11564_, _03198_);
  or _64471_ (_12982_, _12981_, _04539_);
  or _64472_ (_12983_, _12982_, _12980_);
  or _64473_ (_12984_, _12823_, _04558_);
  and _64474_ (_12985_, _12984_, _11955_);
  and _64475_ (_12986_, _12985_, _12983_);
  and _64476_ (_12987_, _03616_, _03195_);
  or _64477_ (_12988_, _06767_, _06763_);
  nor _64478_ (_12989_, _11955_, _06768_);
  and _64479_ (_12990_, _12989_, _12988_);
  or _64480_ (_12991_, _12990_, _12987_);
  or _64481_ (_12992_, _12991_, _12986_);
  not _64482_ (_12993_, _12987_);
  nor _64483_ (_12994_, _06788_, _06730_);
  nor _64484_ (_12995_, _12994_, _07999_);
  nor _64485_ (_12996_, _12995_, _12993_);
  nor _64486_ (_12997_, _12996_, _04256_);
  and _64487_ (_12998_, _12997_, _12992_);
  and _64488_ (_12999_, _12995_, _04256_);
  or _64489_ (_13000_, _12999_, _03448_);
  or _64490_ (_13001_, _13000_, _12998_);
  nor _64491_ (_13002_, _05825_, _05720_);
  nor _64492_ (_13003_, _13002_, _05826_);
  or _64493_ (_13004_, _13003_, _04713_);
  and _64494_ (_13005_, _13004_, _12174_);
  and _64495_ (_13006_, _13005_, _13001_);
  or _64496_ (_13007_, _13006_, _12397_);
  and _64497_ (_13008_, _13007_, _12805_);
  and _64498_ (_13009_, _11390_, _03629_);
  nor _64499_ (_13010_, _11526_, _03629_);
  or _64500_ (_13011_, _13010_, _13009_);
  and _64501_ (_13012_, _13011_, _12195_);
  or _64502_ (_40640_, _13012_, _13008_);
  nor _64503_ (_13013_, _12839_, _05517_);
  nor _64504_ (_13014_, _13013_, _05960_);
  nand _64505_ (_13015_, _13014_, _04531_);
  nor _64506_ (_13016_, _06267_, _05517_);
  and _64507_ (_13017_, _13016_, _04515_);
  nor _64508_ (_13018_, _09850_, _09827_);
  and _64509_ (_13019_, _09827_, \oc8051_golden_model_1.PSW [7]);
  nor _64510_ (_13020_, _13019_, _13018_);
  nor _64511_ (_13021_, _13020_, _05063_);
  nor _64512_ (_13022_, _12812_, _05469_);
  or _64513_ (_13023_, _13022_, _05838_);
  and _64514_ (_13024_, _13023_, _06073_);
  nor _64515_ (_13025_, _03980_, _07478_);
  and _64516_ (_13026_, _11559_, _03980_);
  or _64517_ (_13027_, _13026_, _13025_);
  and _64518_ (_13028_, _13027_, _06072_);
  or _64519_ (_13029_, _13028_, _13024_);
  and _64520_ (_13030_, _13029_, _05966_);
  and _64521_ (_13031_, _06684_, _04422_);
  or _64522_ (_13032_, _13031_, _13030_);
  and _64523_ (_13033_, _13032_, _06071_);
  nor _64524_ (_13034_, _13014_, _06071_);
  or _64525_ (_13035_, _13034_, _13033_);
  and _64526_ (_13036_, _13035_, _05954_);
  nand _64527_ (_13037_, _09828_, _10158_);
  and _64528_ (_13038_, _13037_, _04428_);
  or _64529_ (_13039_, _13038_, _04768_);
  or _64530_ (_13040_, _13039_, _13036_);
  nor _64531_ (_13041_, _11559_, _03230_);
  nor _64532_ (_13042_, _13041_, _04431_);
  and _64533_ (_13043_, _13042_, _13040_);
  and _64534_ (_13044_, _06762_, _04431_);
  or _64535_ (_13045_, _13044_, _04449_);
  or _64536_ (_13046_, _13045_, _13043_);
  nor _64537_ (_13047_, _09827_, _10158_);
  or _64538_ (_13048_, _13047_, _05940_);
  and _64539_ (_13049_, _13048_, _13046_);
  or _64540_ (_13050_, _13049_, _03508_);
  nand _64541_ (_13051_, _08218_, _03508_);
  and _64542_ (_13052_, _13051_, _04562_);
  and _64543_ (_13053_, _13052_, _13050_);
  not _64544_ (_13054_, _10159_);
  and _64545_ (_13055_, _13037_, _13054_);
  and _64546_ (_13056_, _13055_, _04454_);
  or _64547_ (_13057_, _13056_, _13053_);
  and _64548_ (_13058_, _13057_, _03227_);
  nor _64549_ (_13059_, _11560_, _03227_);
  or _64550_ (_13060_, _13059_, _03745_);
  or _64551_ (_13061_, _13060_, _13058_);
  nand _64552_ (_13062_, _08218_, _03745_);
  and _64553_ (_13063_, _13062_, _13061_);
  or _64554_ (_13064_, _13063_, _04463_);
  and _64555_ (_13065_, _06684_, _03446_);
  nand _64556_ (_13066_, _08217_, _04463_);
  or _64557_ (_13067_, _13066_, _13065_);
  and _64558_ (_13068_, _13067_, _05063_);
  and _64559_ (_13069_, _13068_, _13064_);
  or _64560_ (_13070_, _13069_, _13021_);
  and _64561_ (_13071_, _13070_, _05897_);
  nand _64562_ (_13072_, _11559_, _03224_);
  nand _64563_ (_13073_, _13072_, _04480_);
  or _64564_ (_13074_, _13073_, _13071_);
  or _64565_ (_13075_, _06762_, _04480_);
  and _64566_ (_13076_, _13075_, _13074_);
  or _64567_ (_13077_, _13076_, _04482_);
  or _64568_ (_13078_, _06684_, _06164_);
  and _64569_ (_13079_, _13078_, _06163_);
  and _64570_ (_13080_, _13079_, _13077_);
  nor _64571_ (_13081_, _06171_, _05469_);
  and _64572_ (_13082_, _06296_, \oc8051_golden_model_1.IP [5]);
  and _64573_ (_13083_, _06310_, \oc8051_golden_model_1.B [5]);
  nor _64574_ (_13084_, _13083_, _13082_);
  and _64575_ (_13085_, _06303_, \oc8051_golden_model_1.PSW [5]);
  and _64576_ (_13086_, _06308_, \oc8051_golden_model_1.ACC [5]);
  nor _64577_ (_13087_, _13086_, _13085_);
  and _64578_ (_13088_, _13087_, _13084_);
  and _64579_ (_13089_, _06288_, \oc8051_golden_model_1.TH1 [5]);
  not _64580_ (_13090_, _13089_);
  and _64581_ (_13091_, _06354_, \oc8051_golden_model_1.SP [5]);
  and _64582_ (_13092_, _06284_, \oc8051_golden_model_1.TL0 [5]);
  nor _64583_ (_13093_, _13092_, _13091_);
  and _64584_ (_13094_, _13093_, _13090_);
  and _64585_ (_13095_, _13094_, _13088_);
  and _64586_ (_13096_, _06327_, \oc8051_golden_model_1.TH0 [5]);
  and _64587_ (_13097_, _06329_, \oc8051_golden_model_1.TL1 [5]);
  nor _64588_ (_13098_, _13097_, _13096_);
  and _64589_ (_13099_, _06334_, \oc8051_golden_model_1.PCON [5]);
  and _64590_ (_13100_, _06336_, \oc8051_golden_model_1.TCON [5]);
  nor _64591_ (_13101_, _13100_, _13099_);
  and _64592_ (_13102_, _13101_, _13098_);
  and _64593_ (_13103_, _06356_, \oc8051_golden_model_1.DPL [5]);
  not _64594_ (_13104_, _13103_);
  and _64595_ (_13105_, _06343_, \oc8051_golden_model_1.P0INREG [5]);
  not _64596_ (_13106_, _13105_);
  and _64597_ (_13107_, _06348_, \oc8051_golden_model_1.P3INREG [5]);
  and _64598_ (_13108_, _06340_, \oc8051_golden_model_1.P1INREG [5]);
  and _64599_ (_13109_, _06346_, \oc8051_golden_model_1.P2INREG [5]);
  or _64600_ (_13110_, _13109_, _13108_);
  nor _64601_ (_13111_, _13110_, _13107_);
  and _64602_ (_13112_, _13111_, _13106_);
  and _64603_ (_13113_, _13112_, _13104_);
  and _64604_ (_13114_, _06315_, \oc8051_golden_model_1.IE [5]);
  and _64605_ (_13115_, _06319_, \oc8051_golden_model_1.SBUF [5]);
  and _64606_ (_13116_, _06321_, \oc8051_golden_model_1.SCON [5]);
  or _64607_ (_13117_, _13116_, _13115_);
  nor _64608_ (_13118_, _13117_, _13114_);
  and _64609_ (_13119_, _06272_, \oc8051_golden_model_1.DPH [5]);
  and _64610_ (_13120_, _06279_, \oc8051_golden_model_1.TMOD [5]);
  nor _64611_ (_13121_, _13120_, _13119_);
  and _64612_ (_13122_, _13121_, _13118_);
  and _64613_ (_13123_, _13122_, _13113_);
  and _64614_ (_13124_, _13123_, _13102_);
  and _64615_ (_13125_, _13124_, _13095_);
  not _64616_ (_13126_, _13125_);
  nor _64617_ (_13127_, _13126_, _13081_);
  nor _64618_ (_13128_, _13127_, _06170_);
  or _64619_ (_13129_, _13128_, _06168_);
  or _64620_ (_13130_, _13129_, _13080_);
  and _64621_ (_13131_, _06168_, _03860_);
  nor _64622_ (_13132_, _13131_, _04500_);
  and _64623_ (_13133_, _13132_, _13130_);
  and _64624_ (_13134_, _06306_, _04500_);
  or _64625_ (_13135_, _13134_, _03178_);
  or _64626_ (_13136_, _13135_, _13133_);
  and _64627_ (_13137_, _11560_, _03178_);
  nor _64628_ (_13138_, _13137_, _04512_);
  and _64629_ (_13139_, _13138_, _13136_);
  and _64630_ (_13140_, _06267_, _05517_);
  nor _64631_ (_13141_, _13140_, _13016_);
  nor _64632_ (_13142_, _13141_, _04511_);
  nor _64633_ (_13143_, _13142_, _04513_);
  or _64634_ (_13144_, _13143_, _13139_);
  nor _64635_ (_13145_, _05517_, _07478_);
  and _64636_ (_13146_, _05517_, _07478_);
  nor _64637_ (_13147_, _13146_, _13145_);
  or _64638_ (_13148_, _13147_, _05850_);
  and _64639_ (_13149_, _13148_, _06383_);
  and _64640_ (_13150_, _13149_, _13144_);
  or _64641_ (_13151_, _13150_, _13017_);
  and _64642_ (_13152_, _13151_, _06382_);
  and _64643_ (_13153_, _13145_, _04514_);
  or _64644_ (_13154_, _13153_, _03192_);
  or _64645_ (_13155_, _13154_, _13152_);
  and _64646_ (_13156_, _11560_, _03192_);
  nor _64647_ (_13157_, _13156_, _06390_);
  and _64648_ (_13158_, _13157_, _13155_);
  nor _64649_ (_13159_, _13140_, _06395_);
  or _64650_ (_13160_, _13159_, _06394_);
  or _64651_ (_13161_, _13160_, _13158_);
  nand _64652_ (_13162_, _13146_, _06394_);
  and _64653_ (_13163_, _13162_, _06399_);
  and _64654_ (_13164_, _13163_, _13161_);
  nand _64655_ (_13165_, _11559_, _03188_);
  nand _64656_ (_13166_, _13165_, _05848_);
  or _64657_ (_13167_, _13166_, _13164_);
  and _64658_ (_13168_, _13023_, _06409_);
  or _64659_ (_13169_, _13168_, _11933_);
  and _64660_ (_13170_, _13169_, _13167_);
  not _64661_ (_13171_, _06684_);
  nor _64662_ (_13172_, _12807_, _13171_);
  or _64663_ (_13173_, _13172_, _06732_);
  and _64664_ (_13174_, _13173_, _04533_);
  or _64665_ (_13175_, _13174_, _04531_);
  or _64666_ (_13176_, _13175_, _13170_);
  and _64667_ (_13177_, _13176_, _13015_);
  or _64668_ (_13178_, _13177_, _03629_);
  nand _64669_ (_13179_, _11426_, _03629_);
  and _64670_ (_13180_, _13179_, _12371_);
  and _64671_ (_13181_, _13180_, _13178_);
  and _64672_ (_13182_, _11559_, _03198_);
  or _64673_ (_13183_, _13182_, _04539_);
  or _64674_ (_13184_, _13183_, _13181_);
  or _64675_ (_13185_, _13018_, _04558_);
  and _64676_ (_13186_, _13185_, _11955_);
  and _64677_ (_13187_, _13186_, _13184_);
  nor _64678_ (_13188_, _06768_, _06762_);
  or _64679_ (_13189_, _13188_, _06769_);
  nor _64680_ (_13190_, _13189_, _11955_);
  or _64681_ (_13191_, _13190_, _04552_);
  or _64682_ (_13192_, _13191_, _13187_);
  nor _64683_ (_13193_, _07999_, _06684_);
  nor _64684_ (_13194_, _13193_, _06790_);
  or _64685_ (_13195_, _13194_, _06785_);
  and _64686_ (_13196_, _13195_, _13192_);
  or _64687_ (_13197_, _13196_, _03448_);
  nor _64688_ (_13198_, _05826_, _05518_);
  nor _64689_ (_13199_, _13198_, _05827_);
  or _64690_ (_13200_, _13199_, _04713_);
  and _64691_ (_13201_, _13200_, _04796_);
  and _64692_ (_13202_, _13201_, _13197_);
  or _64693_ (_13203_, _13202_, _11999_);
  or _64694_ (_13204_, _11998_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _64695_ (_13205_, _13204_, _12188_);
  and _64696_ (_13206_, _13205_, _13203_);
  and _64697_ (_13207_, _11385_, _03629_);
  and _64698_ (_13208_, _11521_, _11944_);
  or _64699_ (_13209_, _13208_, _13207_);
  and _64700_ (_13210_, _13209_, _12195_);
  or _64701_ (_40641_, _13210_, _13206_);
  or _64702_ (_13211_, _12183_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _64703_ (_13212_, _13211_, _12200_);
  nor _64704_ (_13213_, _06790_, _06455_);
  nor _64705_ (_13214_, _13213_, _06791_);
  or _64706_ (_13215_, _13214_, _06785_);
  nor _64707_ (_13216_, _06732_, _06456_);
  or _64708_ (_13217_, _13216_, _06733_);
  and _64709_ (_13218_, _13217_, _04533_);
  nor _64710_ (_13219_, _05838_, _05363_);
  or _64711_ (_13220_, _13219_, _05839_);
  or _64712_ (_13221_, _13220_, _05847_);
  nor _64713_ (_13222_, _06204_, _05411_);
  and _64714_ (_13223_, _13222_, _04515_);
  nor _64715_ (_13224_, _09799_, _09775_);
  and _64716_ (_13225_, _09775_, \oc8051_golden_model_1.PSW [7]);
  nor _64717_ (_13226_, _13225_, _13224_);
  nor _64718_ (_13227_, _13226_, _05063_);
  and _64719_ (_13228_, _07818_, _04431_);
  nand _64720_ (_13229_, _09776_, _10133_);
  or _64721_ (_13230_, _13229_, _05954_);
  or _64722_ (_13231_, _13220_, _06072_);
  and _64723_ (_13232_, _11551_, _03980_);
  nor _64724_ (_13233_, _03980_, _07433_);
  or _64725_ (_13234_, _13233_, _06073_);
  or _64726_ (_13235_, _13234_, _13232_);
  and _64727_ (_13236_, _13235_, _13231_);
  or _64728_ (_13237_, _13236_, _04422_);
  or _64729_ (_13238_, _06455_, _05966_);
  and _64730_ (_13239_, _13238_, _13237_);
  or _64731_ (_13240_, _13239_, _04421_);
  nor _64732_ (_13241_, _05960_, _05411_);
  nor _64733_ (_13242_, _13241_, _05961_);
  nand _64734_ (_13243_, _13242_, _04421_);
  and _64735_ (_13244_, _13243_, _13240_);
  or _64736_ (_13245_, _13244_, _04428_);
  and _64737_ (_13246_, _13245_, _13230_);
  or _64738_ (_13247_, _13246_, _04768_);
  nor _64739_ (_13248_, _11551_, _03230_);
  nor _64740_ (_13249_, _13248_, _04431_);
  and _64741_ (_13250_, _13249_, _13247_);
  or _64742_ (_13251_, _13250_, _13228_);
  and _64743_ (_13252_, _13251_, _05940_);
  nor _64744_ (_13253_, _09775_, _10133_);
  and _64745_ (_13254_, _13253_, _04449_);
  or _64746_ (_13255_, _13254_, _03508_);
  or _64747_ (_13256_, _13255_, _13252_);
  nand _64748_ (_13257_, _08203_, _03508_);
  and _64749_ (_13258_, _13257_, _04562_);
  and _64750_ (_13259_, _13258_, _13256_);
  not _64751_ (_13260_, _10134_);
  and _64752_ (_13261_, _13229_, _13260_);
  and _64753_ (_13262_, _13261_, _04454_);
  or _64754_ (_13263_, _13262_, _13259_);
  and _64755_ (_13264_, _13263_, _03227_);
  nor _64756_ (_13265_, _11552_, _03227_);
  or _64757_ (_13266_, _13265_, _03745_);
  or _64758_ (_13267_, _13266_, _13264_);
  nand _64759_ (_13268_, _08203_, _03745_);
  and _64760_ (_13269_, _13268_, _13267_);
  or _64761_ (_13270_, _13269_, _04463_);
  and _64762_ (_13271_, _06455_, _03446_);
  nand _64763_ (_13272_, _08202_, _04463_);
  or _64764_ (_13273_, _13272_, _13271_);
  and _64765_ (_13274_, _13273_, _05063_);
  and _64766_ (_13275_, _13274_, _13270_);
  or _64767_ (_13276_, _13275_, _13227_);
  and _64768_ (_13277_, _13276_, _05897_);
  nand _64769_ (_13278_, _11551_, _03224_);
  nand _64770_ (_13279_, _13278_, _04480_);
  or _64771_ (_13280_, _13279_, _13277_);
  or _64772_ (_13281_, _07818_, _04480_);
  and _64773_ (_13282_, _13281_, _13280_);
  or _64774_ (_13283_, _13282_, _04482_);
  or _64775_ (_13284_, _06455_, _06164_);
  and _64776_ (_13285_, _13284_, _06163_);
  and _64777_ (_13286_, _13285_, _13283_);
  nor _64778_ (_13287_, _06171_, _05363_);
  and _64779_ (_13288_, _06272_, \oc8051_golden_model_1.DPH [6]);
  and _64780_ (_13289_, _06288_, \oc8051_golden_model_1.TH1 [6]);
  nor _64781_ (_13290_, _13289_, _13288_);
  and _64782_ (_13291_, _06340_, \oc8051_golden_model_1.P1INREG [6]);
  not _64783_ (_13292_, _13291_);
  and _64784_ (_13293_, _06343_, \oc8051_golden_model_1.P0INREG [6]);
  not _64785_ (_13294_, _13293_);
  and _64786_ (_13295_, _06346_, \oc8051_golden_model_1.P2INREG [6]);
  and _64787_ (_13296_, _06348_, \oc8051_golden_model_1.P3INREG [6]);
  nor _64788_ (_13297_, _13296_, _13295_);
  and _64789_ (_13298_, _13297_, _13294_);
  and _64790_ (_13299_, _13298_, _13292_);
  and _64791_ (_13300_, _13299_, _13290_);
  and _64792_ (_13301_, _06315_, \oc8051_golden_model_1.IE [6]);
  and _64793_ (_13302_, _06319_, \oc8051_golden_model_1.SBUF [6]);
  and _64794_ (_13303_, _06321_, \oc8051_golden_model_1.SCON [6]);
  or _64795_ (_13304_, _13303_, _13302_);
  nor _64796_ (_13305_, _13304_, _13301_);
  and _64797_ (_13306_, _06296_, \oc8051_golden_model_1.IP [6]);
  and _64798_ (_13307_, _06310_, \oc8051_golden_model_1.B [6]);
  nor _64799_ (_13308_, _13307_, _13306_);
  and _64800_ (_13309_, _06303_, \oc8051_golden_model_1.PSW [6]);
  and _64801_ (_13310_, _06308_, \oc8051_golden_model_1.ACC [6]);
  nor _64802_ (_13311_, _13310_, _13309_);
  and _64803_ (_13312_, _13311_, _13308_);
  and _64804_ (_13313_, _13312_, _13305_);
  and _64805_ (_13314_, _13313_, _13300_);
  and _64806_ (_13315_, _06327_, \oc8051_golden_model_1.TH0 [6]);
  and _64807_ (_13316_, _06329_, \oc8051_golden_model_1.TL1 [6]);
  nor _64808_ (_13317_, _13316_, _13315_);
  and _64809_ (_13318_, _06334_, \oc8051_golden_model_1.PCON [6]);
  and _64810_ (_13319_, _06336_, \oc8051_golden_model_1.TCON [6]);
  nor _64811_ (_13320_, _13319_, _13318_);
  and _64812_ (_13321_, _13320_, _13317_);
  and _64813_ (_13322_, _06354_, \oc8051_golden_model_1.SP [6]);
  and _64814_ (_13323_, _06356_, \oc8051_golden_model_1.DPL [6]);
  nor _64815_ (_13324_, _13323_, _13322_);
  and _64816_ (_13325_, _06284_, \oc8051_golden_model_1.TL0 [6]);
  and _64817_ (_13326_, _06279_, \oc8051_golden_model_1.TMOD [6]);
  nor _64818_ (_13327_, _13326_, _13325_);
  and _64819_ (_13328_, _13327_, _13324_);
  and _64820_ (_13329_, _13328_, _13321_);
  and _64821_ (_13330_, _13329_, _13314_);
  not _64822_ (_13331_, _13330_);
  nor _64823_ (_13332_, _13331_, _13287_);
  nor _64824_ (_13333_, _13332_, _06170_);
  or _64825_ (_13334_, _13333_, _06168_);
  or _64826_ (_13335_, _13334_, _13286_);
  and _64827_ (_13336_, _06168_, _03549_);
  nor _64828_ (_13337_, _13336_, _04500_);
  and _64829_ (_13338_, _13337_, _13335_);
  not _64830_ (_13339_, _06204_);
  and _64831_ (_13340_, _13339_, _04500_);
  or _64832_ (_13341_, _13340_, _03178_);
  or _64833_ (_13342_, _13341_, _13338_);
  and _64834_ (_13343_, _11552_, _03178_);
  nor _64835_ (_13344_, _13343_, _04512_);
  and _64836_ (_13345_, _13344_, _13342_);
  and _64837_ (_13346_, _06204_, _05411_);
  nor _64838_ (_13347_, _13346_, _13222_);
  nor _64839_ (_13348_, _13347_, _04511_);
  nor _64840_ (_13349_, _13348_, _04513_);
  or _64841_ (_13350_, _13349_, _13345_);
  nor _64842_ (_13351_, _05411_, _07433_);
  and _64843_ (_13352_, _05411_, _07433_);
  nor _64844_ (_13353_, _13352_, _13351_);
  or _64845_ (_13354_, _13353_, _05850_);
  and _64846_ (_13355_, _13354_, _06383_);
  and _64847_ (_13356_, _13355_, _13350_);
  or _64848_ (_13357_, _13356_, _13223_);
  and _64849_ (_13358_, _13357_, _06382_);
  and _64850_ (_13359_, _13351_, _04514_);
  or _64851_ (_13360_, _13359_, _03192_);
  or _64852_ (_13361_, _13360_, _13358_);
  and _64853_ (_13362_, _11552_, _03192_);
  nor _64854_ (_13363_, _13362_, _06390_);
  and _64855_ (_13364_, _13363_, _13361_);
  nor _64856_ (_13365_, _13346_, _06395_);
  or _64857_ (_13366_, _13365_, _06394_);
  or _64858_ (_13367_, _13366_, _13364_);
  nand _64859_ (_13368_, _13352_, _06394_);
  and _64860_ (_13369_, _13368_, _06399_);
  and _64861_ (_13370_, _13369_, _13367_);
  nand _64862_ (_13371_, _11551_, _03188_);
  nand _64863_ (_13372_, _13371_, _05847_);
  or _64864_ (_13373_, _13372_, _13370_);
  and _64865_ (_13374_, _13373_, _13221_);
  or _64866_ (_13375_, _13374_, _03495_);
  or _64867_ (_13376_, _13220_, _04745_);
  and _64868_ (_13377_, _13376_, _06409_);
  and _64869_ (_13378_, _13377_, _13375_);
  or _64870_ (_13379_, _13378_, _13218_);
  and _64871_ (_13380_, _13379_, _06408_);
  nor _64872_ (_13381_, _13242_, _06408_);
  or _64873_ (_13382_, _13381_, _03629_);
  or _64874_ (_13383_, _13382_, _13380_);
  nand _64875_ (_13384_, _11418_, _03629_);
  and _64876_ (_13385_, _13384_, _12371_);
  and _64877_ (_13386_, _13385_, _13383_);
  and _64878_ (_13387_, _11551_, _03198_);
  or _64879_ (_13388_, _13387_, _04539_);
  or _64880_ (_13389_, _13388_, _13386_);
  or _64881_ (_13390_, _13224_, _04558_);
  and _64882_ (_13391_, _13390_, _11955_);
  and _64883_ (_13392_, _13391_, _13389_);
  nand _64884_ (_13393_, _06769_, _07818_);
  or _64885_ (_13394_, _06769_, _07818_);
  and _64886_ (_13395_, _13394_, _11956_);
  and _64887_ (_13396_, _13395_, _13393_);
  or _64888_ (_13397_, _13396_, _04552_);
  or _64889_ (_13398_, _13397_, _13392_);
  and _64890_ (_13399_, _13398_, _13215_);
  or _64891_ (_13400_, _13399_, _03448_);
  nor _64892_ (_13401_, _05827_, _05412_);
  nor _64893_ (_13402_, _13401_, _05828_);
  or _64894_ (_13403_, _13402_, _04713_);
  and _64895_ (_13404_, _13403_, _12174_);
  and _64896_ (_13405_, _13404_, _13400_);
  or _64897_ (_13406_, _13405_, _12397_);
  and _64898_ (_13407_, _13406_, _13212_);
  and _64899_ (_13408_, _11514_, _11944_);
  and _64900_ (_13409_, _11378_, _03629_);
  or _64901_ (_13410_, _13409_, _13408_);
  and _64902_ (_13411_, _13410_, _12195_);
  or _64903_ (_40642_, _13411_, _13407_);
  nor _64904_ (_13412_, _12183_, _05144_);
  nor _64905_ (_13413_, _12397_, _06799_);
  or _64906_ (_13414_, _13413_, _13412_);
  and _64907_ (_13415_, _13414_, _12200_);
  and _64908_ (_13416_, _12195_, _06823_);
  or _64909_ (_40644_, _13416_, _13415_);
  and _64910_ (_13417_, _04798_, _04556_);
  and _64911_ (_13418_, _13417_, _11996_);
  not _64912_ (_13419_, _13418_);
  or _64913_ (_13420_, _13419_, _12171_);
  or _64914_ (_13421_, _13418_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand _64915_ (_13422_, _12187_, _04804_);
  and _64916_ (_13423_, _13422_, _13421_);
  and _64917_ (_13424_, _13423_, _13420_);
  and _64918_ (_13425_, _12194_, _04804_);
  and _64919_ (_13426_, _13425_, _12198_);
  or _64920_ (_40648_, _13426_, _13424_);
  not _64921_ (_13427_, _13425_);
  or _64922_ (_13428_, _13418_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _64923_ (_13429_, _13428_, _13427_);
  or _64924_ (_13430_, _13419_, _12388_);
  and _64925_ (_13431_, _13430_, _13429_);
  and _64926_ (_13432_, _13425_, _12393_);
  or _64927_ (_40649_, _13432_, _13431_);
  or _64928_ (_13433_, _13418_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _64929_ (_13434_, _13433_, _13427_);
  and _64930_ (_13435_, _12593_, _04796_);
  and _64931_ (_13436_, _13435_, _12590_);
  or _64932_ (_13437_, _13419_, _13436_);
  and _64933_ (_13438_, _13437_, _13434_);
  and _64934_ (_13439_, _13425_, _12600_);
  or _64935_ (_40650_, _13439_, _13438_);
  or _64936_ (_13440_, _13418_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _64937_ (_13441_, _13440_, _13427_);
  and _64938_ (_13442_, _12795_, _04796_);
  and _64939_ (_13443_, _13442_, _12792_);
  or _64940_ (_13444_, _13419_, _13443_);
  and _64941_ (_13445_, _13444_, _13441_);
  and _64942_ (_13446_, _13425_, _12802_);
  or _64943_ (_40651_, _13446_, _13445_);
  or _64944_ (_13447_, _13418_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _64945_ (_13448_, _13447_, _13427_);
  and _64946_ (_13449_, _13004_, _04796_);
  and _64947_ (_13450_, _13449_, _13001_);
  or _64948_ (_13451_, _13419_, _13450_);
  and _64949_ (_13452_, _13451_, _13448_);
  and _64950_ (_13453_, _13425_, _13011_);
  or _64951_ (_40653_, _13453_, _13452_);
  or _64952_ (_13454_, _13418_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _64953_ (_13455_, _13454_, _13427_);
  or _64954_ (_13456_, _13419_, _13202_);
  and _64955_ (_13457_, _13456_, _13455_);
  and _64956_ (_13458_, _13425_, _13209_);
  or _64957_ (_40654_, _13458_, _13457_);
  or _64958_ (_13459_, _13418_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _64959_ (_13460_, _13459_, _13427_);
  and _64960_ (_13461_, _13403_, _04796_);
  and _64961_ (_13462_, _13461_, _13400_);
  or _64962_ (_13463_, _13419_, _13462_);
  and _64963_ (_13464_, _13463_, _13460_);
  and _64964_ (_13465_, _13425_, _13410_);
  or _64965_ (_40655_, _13465_, _13464_);
  or _64966_ (_13466_, _13418_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _64967_ (_13467_, _13466_, _13427_);
  or _64968_ (_13468_, _13419_, _06800_);
  and _64969_ (_13469_, _13468_, _13467_);
  and _64970_ (_13470_, _13425_, _06823_);
  or _64971_ (_40656_, _13470_, _13469_);
  and _64972_ (_13471_, _11993_, _04711_);
  and _64973_ (_13472_, _13471_, _11996_);
  not _64974_ (_13473_, _13472_);
  or _64975_ (_13474_, _13473_, _12171_);
  and _64976_ (_13475_, _12187_, _05967_);
  not _64977_ (_13476_, _13475_);
  or _64978_ (_13477_, _13472_, \oc8051_golden_model_1.IRAM[2] [0]);
  and _64979_ (_13478_, _13477_, _13476_);
  and _64980_ (_13479_, _13478_, _13474_);
  and _64981_ (_13480_, _12198_, _05137_);
  and _64982_ (_13481_, _13480_, _13475_);
  or _64983_ (_40661_, _13481_, _13479_);
  or _64984_ (_13482_, _13473_, _12388_);
  or _64985_ (_13483_, _13472_, \oc8051_golden_model_1.IRAM[2] [1]);
  and _64986_ (_13484_, _13483_, _13476_);
  and _64987_ (_13485_, _13484_, _13482_);
  and _64988_ (_13486_, _12393_, _05137_);
  and _64989_ (_13487_, _13486_, _13475_);
  or _64990_ (_40662_, _13487_, _13485_);
  and _64991_ (_13488_, _12194_, _05967_);
  not _64992_ (_13489_, _13488_);
  and _64993_ (_13490_, _12179_, _04711_);
  and _64994_ (_13491_, _13490_, _12178_);
  or _64995_ (_13492_, _13491_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _64996_ (_13493_, _13492_, _13489_);
  not _64997_ (_13494_, _13491_);
  or _64998_ (_13495_, _13494_, _12595_);
  and _64999_ (_13496_, _13495_, _13493_);
  and _65000_ (_13497_, _12600_, _12191_);
  and _65001_ (_13498_, _13497_, _13488_);
  or _65002_ (_40663_, _13498_, _13496_);
  or _65003_ (_13499_, _13491_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _65004_ (_13500_, _13499_, _13489_);
  or _65005_ (_13501_, _13494_, _12797_);
  and _65006_ (_13502_, _13501_, _13500_);
  and _65007_ (_13503_, _12802_, _12191_);
  and _65008_ (_13504_, _13503_, _13488_);
  or _65009_ (_40664_, _13504_, _13502_);
  or _65010_ (_13505_, _13491_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _65011_ (_13506_, _13505_, _13489_);
  or _65012_ (_13507_, _13494_, _13006_);
  and _65013_ (_13508_, _13507_, _13506_);
  and _65014_ (_13509_, _13011_, _12191_);
  and _65015_ (_13510_, _13509_, _13488_);
  or _65016_ (_40665_, _13510_, _13508_);
  or _65017_ (_13511_, _13491_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _65018_ (_13512_, _13511_, _13489_);
  and _65019_ (_13513_, _13200_, _12174_);
  and _65020_ (_13514_, _13513_, _13197_);
  or _65021_ (_13515_, _13494_, _13514_);
  and _65022_ (_13516_, _13515_, _13512_);
  and _65023_ (_13517_, _13209_, _12191_);
  and _65024_ (_13518_, _13517_, _13488_);
  or _65025_ (_40667_, _13518_, _13516_);
  or _65026_ (_13519_, _13491_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _65027_ (_13520_, _13519_, _13489_);
  or _65028_ (_13521_, _13494_, _13405_);
  and _65029_ (_13522_, _13521_, _13520_);
  and _65030_ (_13523_, _13410_, _12191_);
  and _65031_ (_13524_, _13523_, _13488_);
  or _65032_ (_40668_, _13524_, _13522_);
  or _65033_ (_13525_, _13491_, \oc8051_golden_model_1.IRAM[2] [7]);
  and _65034_ (_13526_, _13525_, _13489_);
  nor _65035_ (_13527_, _06799_, _12175_);
  or _65036_ (_13528_, _13494_, _13527_);
  and _65037_ (_13529_, _13528_, _13526_);
  and _65038_ (_13530_, _06823_, _12191_);
  and _65039_ (_13531_, _13488_, _13530_);
  or _65040_ (_40669_, _13531_, _13529_);
  and _65041_ (_13532_, _11996_, _04799_);
  not _65042_ (_13533_, _13532_);
  or _65043_ (_13534_, _13533_, _12171_);
  and _65044_ (_13535_, _12187_, _03497_);
  not _65045_ (_13536_, _13535_);
  or _65046_ (_13537_, _13532_, \oc8051_golden_model_1.IRAM[3] [0]);
  and _65047_ (_13538_, _13537_, _13536_);
  and _65048_ (_13539_, _13538_, _13534_);
  and _65049_ (_13540_, _13535_, _13480_);
  or _65050_ (_40673_, _13540_, _13539_);
  or _65051_ (_13541_, _13533_, _12388_);
  or _65052_ (_13542_, _13532_, \oc8051_golden_model_1.IRAM[3] [1]);
  and _65053_ (_13543_, _13542_, _13536_);
  and _65054_ (_13544_, _13543_, _13541_);
  and _65055_ (_13545_, _13535_, _13486_);
  or _65056_ (_40674_, _13545_, _13544_);
  and _65057_ (_13546_, _12194_, _03497_);
  not _65058_ (_13547_, _13546_);
  not _65059_ (_13548_, _12179_);
  nor _65060_ (_13549_, _13548_, _04711_);
  and _65061_ (_13550_, _12178_, _13549_);
  or _65062_ (_13551_, _13550_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _65063_ (_13552_, _13551_, _13547_);
  not _65064_ (_13553_, _13550_);
  or _65065_ (_13554_, _13553_, _12595_);
  and _65066_ (_13555_, _13554_, _13552_);
  and _65067_ (_13556_, _13546_, _13497_);
  or _65068_ (_40675_, _13556_, _13555_);
  or _65069_ (_13557_, _13550_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _65070_ (_13558_, _13557_, _13547_);
  or _65071_ (_13559_, _13553_, _12797_);
  and _65072_ (_13560_, _13559_, _13558_);
  and _65073_ (_13561_, _13546_, _13503_);
  or _65074_ (_40676_, _13561_, _13560_);
  or _65075_ (_13562_, _13550_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _65076_ (_13563_, _13562_, _13547_);
  or _65077_ (_13564_, _13553_, _13006_);
  and _65078_ (_13565_, _13564_, _13563_);
  and _65079_ (_13566_, _13546_, _13509_);
  or _65080_ (_40678_, _13566_, _13565_);
  or _65081_ (_13567_, _13550_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _65082_ (_13568_, _13567_, _13547_);
  or _65083_ (_13569_, _13553_, _13514_);
  and _65084_ (_13570_, _13569_, _13568_);
  and _65085_ (_13571_, _13546_, _13517_);
  or _65086_ (_40679_, _13571_, _13570_);
  or _65087_ (_13572_, _13550_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _65088_ (_13573_, _13572_, _13547_);
  or _65089_ (_13574_, _13553_, _13405_);
  and _65090_ (_13575_, _13574_, _13573_);
  and _65091_ (_13576_, _13546_, _13523_);
  or _65092_ (_40680_, _13576_, _13575_);
  or _65093_ (_13577_, _13550_, \oc8051_golden_model_1.IRAM[3] [7]);
  and _65094_ (_13578_, _13577_, _13547_);
  or _65095_ (_13579_, _13553_, _13527_);
  and _65096_ (_13580_, _13579_, _13578_);
  and _65097_ (_13581_, _13546_, _13530_);
  or _65098_ (_40681_, _13581_, _13580_);
  and _65099_ (_13582_, _11995_, _05122_);
  and _65100_ (_13583_, _13582_, _11994_);
  not _65101_ (_13584_, _13583_);
  or _65102_ (_13585_, _13584_, _12171_);
  and _65103_ (_13586_, _12185_, _05132_);
  and _65104_ (_13587_, _13586_, _03499_);
  not _65105_ (_13588_, _13587_);
  or _65106_ (_13589_, _13583_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _65107_ (_13590_, _13589_, _13588_);
  and _65108_ (_13591_, _13590_, _13585_);
  and _65109_ (_13592_, _13587_, _13480_);
  or _65110_ (_40686_, _13592_, _13591_);
  or _65111_ (_13593_, _13584_, _12388_);
  or _65112_ (_13594_, _13583_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _65113_ (_13595_, _13594_, _13588_);
  and _65114_ (_13596_, _13595_, _13593_);
  and _65115_ (_13597_, _13587_, _13486_);
  or _65116_ (_40687_, _13597_, _13596_);
  and _65117_ (_13598_, _12191_, _05129_);
  and _65118_ (_13599_, _13598_, _05132_);
  and _65119_ (_13600_, _13599_, _03499_);
  not _65120_ (_13601_, _13600_);
  and _65121_ (_13602_, _12176_, _05122_);
  and _65122_ (_13603_, _13602_, _12181_);
  or _65123_ (_13604_, _13603_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _65124_ (_13605_, _13604_, _13601_);
  not _65125_ (_13606_, _13603_);
  or _65126_ (_13607_, _13606_, _12595_);
  and _65127_ (_13608_, _13607_, _13605_);
  and _65128_ (_13609_, _13600_, _13497_);
  or _65129_ (_40688_, _13609_, _13608_);
  or _65130_ (_13610_, _13603_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _65131_ (_13611_, _13610_, _13601_);
  or _65132_ (_13613_, _13606_, _12797_);
  and _65133_ (_13614_, _13613_, _13611_);
  and _65134_ (_13615_, _13600_, _13503_);
  or _65135_ (_40689_, _13615_, _13614_);
  or _65136_ (_13616_, _13603_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _65137_ (_13617_, _13616_, _13601_);
  or _65138_ (_13618_, _13606_, _13006_);
  and _65139_ (_13619_, _13618_, _13617_);
  and _65140_ (_13620_, _13600_, _13509_);
  or _65141_ (_40690_, _13620_, _13619_);
  or _65142_ (_13622_, _13603_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _65143_ (_13623_, _13622_, _13601_);
  or _65144_ (_13624_, _13606_, _13514_);
  and _65145_ (_13625_, _13624_, _13623_);
  and _65146_ (_13626_, _13600_, _13517_);
  or _65147_ (_40692_, _13626_, _13625_);
  or _65148_ (_13627_, _13603_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _65149_ (_13628_, _13627_, _13601_);
  or _65150_ (_13629_, _13606_, _13405_);
  and _65151_ (_13630_, _13629_, _13628_);
  and _65152_ (_13632_, _13600_, _13523_);
  or _65153_ (_40693_, _13632_, _13630_);
  or _65154_ (_13633_, _13603_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _65155_ (_13634_, _13633_, _13601_);
  or _65156_ (_13635_, _13606_, _13527_);
  and _65157_ (_13636_, _13635_, _13634_);
  and _65158_ (_13637_, _13600_, _13530_);
  or _65159_ (_40694_, _13637_, _13636_);
  and _65160_ (_13638_, _13582_, _13417_);
  not _65161_ (_13639_, _13638_);
  or _65162_ (_13641_, _13639_, _12171_);
  and _65163_ (_13642_, _12180_, _04556_);
  and _65164_ (_13643_, _13602_, _13642_);
  or _65165_ (_13644_, _13643_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _65166_ (_13645_, _13586_, _04804_);
  not _65167_ (_13646_, _13645_);
  and _65168_ (_13647_, _13646_, _13644_);
  and _65169_ (_13648_, _13647_, _13641_);
  and _65170_ (_13649_, _13645_, _13480_);
  or _65171_ (_40698_, _13649_, _13648_);
  or _65172_ (_13651_, _13639_, _12388_);
  or _65173_ (_13652_, _13638_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _65174_ (_13653_, _13652_, _13646_);
  and _65175_ (_13654_, _13653_, _13651_);
  and _65176_ (_13655_, _13645_, _13486_);
  or _65177_ (_40699_, _13655_, _13654_);
  and _65178_ (_13656_, _13599_, _04804_);
  not _65179_ (_13657_, _13656_);
  or _65180_ (_13658_, _13643_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _65181_ (_13659_, _13658_, _13657_);
  not _65182_ (_13661_, _13643_);
  or _65183_ (_13662_, _13661_, _12595_);
  and _65184_ (_13663_, _13662_, _13659_);
  and _65185_ (_13664_, _13656_, _13497_);
  or _65186_ (_40700_, _13664_, _13663_);
  or _65187_ (_13665_, _13643_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _65188_ (_13666_, _13665_, _13657_);
  or _65189_ (_13667_, _13661_, _12797_);
  and _65190_ (_13668_, _13667_, _13666_);
  and _65191_ (_13669_, _13656_, _13503_);
  or _65192_ (_40701_, _13669_, _13668_);
  or _65193_ (_13671_, _13643_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _65194_ (_13672_, _13671_, _13657_);
  or _65195_ (_13673_, _13661_, _13006_);
  and _65196_ (_13674_, _13673_, _13672_);
  and _65197_ (_13675_, _13656_, _13509_);
  or _65198_ (_40702_, _13675_, _13674_);
  or _65199_ (_13676_, _13643_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _65200_ (_13677_, _13676_, _13657_);
  or _65201_ (_13678_, _13661_, _13514_);
  and _65202_ (_13680_, _13678_, _13677_);
  and _65203_ (_13681_, _13656_, _13517_);
  or _65204_ (_40704_, _13681_, _13680_);
  or _65205_ (_13682_, _13643_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _65206_ (_13683_, _13682_, _13657_);
  or _65207_ (_13684_, _13661_, _13405_);
  and _65208_ (_13685_, _13684_, _13683_);
  and _65209_ (_13686_, _13656_, _13523_);
  or _65210_ (_40705_, _13686_, _13685_);
  and _65211_ (_13687_, _13643_, _13527_);
  nor _65212_ (_13689_, _13643_, _05166_);
  or _65213_ (_13690_, _13689_, _13656_);
  or _65214_ (_13691_, _13690_, _13687_);
  or _65215_ (_13692_, _13657_, _13530_);
  and _65216_ (_40706_, _13692_, _13691_);
  and _65217_ (_13693_, _13582_, _13471_);
  not _65218_ (_13694_, _13693_);
  or _65219_ (_13695_, _13694_, _12171_);
  and _65220_ (_13696_, _13586_, _05967_);
  not _65221_ (_13697_, _13696_);
  or _65222_ (_13699_, _13693_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _65223_ (_13700_, _13699_, _13697_);
  and _65224_ (_13701_, _13700_, _13695_);
  and _65225_ (_13702_, _13696_, _13480_);
  or _65226_ (_40710_, _13702_, _13701_);
  or _65227_ (_13703_, _13694_, _12388_);
  or _65228_ (_13704_, _13693_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _65229_ (_13705_, _13704_, _13697_);
  and _65230_ (_13706_, _13705_, _13703_);
  and _65231_ (_13707_, _13696_, _13486_);
  or _65232_ (_40711_, _13707_, _13706_);
  and _65233_ (_13709_, _13599_, _05967_);
  not _65234_ (_13710_, _13709_);
  and _65235_ (_13711_, _13602_, _13490_);
  or _65236_ (_13712_, _13711_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _65237_ (_13713_, _13712_, _13710_);
  not _65238_ (_13714_, _13711_);
  or _65239_ (_13715_, _13714_, _12595_);
  and _65240_ (_13716_, _13715_, _13713_);
  and _65241_ (_13717_, _13709_, _13497_);
  or _65242_ (_40712_, _13717_, _13716_);
  or _65243_ (_13719_, _13711_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _65244_ (_13720_, _13719_, _13710_);
  or _65245_ (_13721_, _13714_, _12797_);
  and _65246_ (_13722_, _13721_, _13720_);
  and _65247_ (_13723_, _13709_, _13503_);
  or _65248_ (_40713_, _13723_, _13722_);
  or _65249_ (_13724_, _13711_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _65250_ (_13725_, _13724_, _13710_);
  or _65251_ (_13726_, _13714_, _13006_);
  and _65252_ (_13728_, _13726_, _13725_);
  and _65253_ (_13729_, _13709_, _13509_);
  or _65254_ (_40715_, _13729_, _13728_);
  or _65255_ (_13730_, _13711_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _65256_ (_13731_, _13730_, _13710_);
  or _65257_ (_13732_, _13714_, _13514_);
  and _65258_ (_13733_, _13732_, _13731_);
  and _65259_ (_13734_, _13709_, _13517_);
  or _65260_ (_40716_, _13734_, _13733_);
  or _65261_ (_13735_, _13711_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _65262_ (_13737_, _13735_, _13710_);
  or _65263_ (_13738_, _13714_, _13405_);
  and _65264_ (_13739_, _13738_, _13737_);
  and _65265_ (_13740_, _13709_, _13523_);
  or _65266_ (_40717_, _13740_, _13739_);
  or _65267_ (_13741_, _13711_, \oc8051_golden_model_1.IRAM[6] [7]);
  and _65268_ (_13742_, _13741_, _13710_);
  or _65269_ (_13743_, _13714_, _13527_);
  and _65270_ (_13744_, _13743_, _13742_);
  and _65271_ (_13745_, _13709_, _13530_);
  or _65272_ (_40718_, _13745_, _13744_);
  and _65273_ (_13746_, _13582_, _04799_);
  not _65274_ (_13747_, _13746_);
  or _65275_ (_13748_, _13747_, _12171_);
  and _65276_ (_13749_, _13586_, _03497_);
  not _65277_ (_13750_, _13749_);
  or _65278_ (_13751_, _13746_, \oc8051_golden_model_1.IRAM[7] [0]);
  and _65279_ (_13752_, _13751_, _13750_);
  and _65280_ (_13753_, _13752_, _13748_);
  and _65281_ (_13754_, _13749_, _13480_);
  or _65282_ (_40722_, _13754_, _13753_);
  or _65283_ (_13755_, _13747_, _12388_);
  or _65284_ (_13756_, _13746_, \oc8051_golden_model_1.IRAM[7] [1]);
  and _65285_ (_13757_, _13756_, _13750_);
  and _65286_ (_13758_, _13757_, _13755_);
  and _65287_ (_13759_, _13749_, _13486_);
  or _65288_ (_40723_, _13759_, _13758_);
  and _65289_ (_13760_, _13599_, _03497_);
  not _65290_ (_13761_, _13760_);
  and _65291_ (_13762_, _13602_, _13549_);
  or _65292_ (_13763_, _13762_, \oc8051_golden_model_1.IRAM[7] [2]);
  and _65293_ (_13764_, _13763_, _13761_);
  not _65294_ (_13765_, _13762_);
  or _65295_ (_13766_, _13765_, _12595_);
  and _65296_ (_13767_, _13766_, _13764_);
  and _65297_ (_13768_, _13760_, _13497_);
  or _65298_ (_40724_, _13768_, _13767_);
  or _65299_ (_13769_, _13762_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _65300_ (_13770_, _13769_, _13761_);
  or _65301_ (_13771_, _13765_, _12797_);
  and _65302_ (_13772_, _13771_, _13770_);
  and _65303_ (_13773_, _13760_, _13503_);
  or _65304_ (_40725_, _13773_, _13772_);
  or _65305_ (_13774_, _13762_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _65306_ (_13775_, _13774_, _13761_);
  or _65307_ (_13776_, _13765_, _13006_);
  and _65308_ (_13777_, _13776_, _13775_);
  and _65309_ (_13778_, _13760_, _13509_);
  or _65310_ (_40727_, _13778_, _13777_);
  or _65311_ (_13779_, _13762_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _65312_ (_13780_, _13779_, _13761_);
  or _65313_ (_13781_, _13765_, _13514_);
  and _65314_ (_13782_, _13781_, _13780_);
  and _65315_ (_13783_, _13760_, _13517_);
  or _65316_ (_40728_, _13783_, _13782_);
  or _65317_ (_13784_, _13762_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _65318_ (_13785_, _13784_, _13761_);
  or _65319_ (_13786_, _13765_, _13405_);
  and _65320_ (_13787_, _13786_, _13785_);
  and _65321_ (_13788_, _13760_, _13523_);
  or _65322_ (_40729_, _13788_, _13787_);
  or _65323_ (_13789_, _13762_, \oc8051_golden_model_1.IRAM[7] [7]);
  and _65324_ (_13790_, _13789_, _13761_);
  or _65325_ (_13791_, _13765_, _13527_);
  and _65326_ (_13792_, _13791_, _13790_);
  and _65327_ (_13793_, _13760_, _13530_);
  or _65328_ (_40730_, _13793_, _13792_);
  and _65329_ (_13794_, _05123_, _04951_);
  and _65330_ (_13795_, _13794_, _11994_);
  not _65331_ (_13796_, _13795_);
  or _65332_ (_13797_, _13796_, _12171_);
  and _65333_ (_13798_, _05138_, _12192_);
  and _65334_ (_13799_, _13798_, _03499_);
  not _65335_ (_13800_, _13799_);
  or _65336_ (_13801_, _13795_, \oc8051_golden_model_1.IRAM[8] [0]);
  and _65337_ (_13802_, _13801_, _13800_);
  and _65338_ (_13803_, _13802_, _13797_);
  and _65339_ (_13804_, _13799_, _13480_);
  or _65340_ (_40735_, _13804_, _13803_);
  or _65341_ (_13805_, _13796_, _12388_);
  or _65342_ (_13806_, _13795_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _65343_ (_13807_, _13806_, _13800_);
  and _65344_ (_13808_, _13807_, _13805_);
  and _65345_ (_13809_, _13799_, _13486_);
  or _65346_ (_40736_, _13809_, _13808_);
  or _65347_ (_13810_, _13795_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _65348_ (_13811_, _13810_, _13800_);
  or _65349_ (_13812_, _13796_, _13436_);
  and _65350_ (_13813_, _13812_, _13811_);
  and _65351_ (_13814_, _12600_, _05137_);
  and _65352_ (_13815_, _13799_, _13814_);
  or _65353_ (_40737_, _13815_, _13813_);
  or _65354_ (_13816_, _13795_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _65355_ (_13817_, _13816_, _13800_);
  or _65356_ (_13818_, _13796_, _13443_);
  and _65357_ (_13819_, _13818_, _13817_);
  and _65358_ (_13820_, _12802_, _05137_);
  and _65359_ (_13821_, _13799_, _13820_);
  or _65360_ (_40738_, _13821_, _13819_);
  or _65361_ (_13822_, _13795_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _65362_ (_13823_, _13822_, _13800_);
  or _65363_ (_13824_, _13796_, _13450_);
  and _65364_ (_13825_, _13824_, _13823_);
  and _65365_ (_13826_, _13011_, _05137_);
  and _65366_ (_13827_, _13799_, _13826_);
  or _65367_ (_40739_, _13827_, _13825_);
  or _65368_ (_13828_, _13795_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _65369_ (_13829_, _13828_, _13800_);
  or _65370_ (_13830_, _13796_, _13202_);
  and _65371_ (_13831_, _13830_, _13829_);
  and _65372_ (_13832_, _13209_, _05137_);
  and _65373_ (_13833_, _13799_, _13832_);
  or _65374_ (_40741_, _13833_, _13831_);
  or _65375_ (_13834_, _13795_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _65376_ (_13835_, _13834_, _13800_);
  or _65377_ (_13836_, _13796_, _13462_);
  and _65378_ (_13837_, _13836_, _13835_);
  and _65379_ (_13838_, _13410_, _05137_);
  and _65380_ (_13839_, _13799_, _13838_);
  or _65381_ (_40742_, _13839_, _13837_);
  nor _65382_ (_13840_, _13795_, \oc8051_golden_model_1.IRAM[8] [7]);
  nor _65383_ (_13841_, _13796_, _06800_);
  or _65384_ (_13842_, _13841_, _13840_);
  nor _65385_ (_13843_, _13842_, _13799_);
  and _65386_ (_13844_, _13799_, _06824_);
  or _65387_ (_40743_, _13844_, _13843_);
  and _65388_ (_13845_, _13794_, _13417_);
  not _65389_ (_13846_, _13845_);
  or _65390_ (_13847_, _13846_, _12171_);
  or _65391_ (_13848_, _13845_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _65392_ (_13849_, _13798_, _04804_);
  not _65393_ (_13850_, _13849_);
  and _65394_ (_13851_, _13850_, _13848_);
  and _65395_ (_13852_, _13851_, _13847_);
  and _65396_ (_13853_, _13849_, _13480_);
  or _65397_ (_40747_, _13853_, _13852_);
  or _65398_ (_13854_, _13846_, _12388_);
  or _65399_ (_13855_, _13845_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _65400_ (_13856_, _13855_, _13850_);
  and _65401_ (_13857_, _13856_, _13854_);
  and _65402_ (_13858_, _13849_, _13486_);
  or _65403_ (_40748_, _13858_, _13857_);
  or _65404_ (_13859_, _13845_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _65405_ (_13860_, _13859_, _13850_);
  or _65406_ (_13861_, _13846_, _13436_);
  and _65407_ (_13862_, _13861_, _13860_);
  and _65408_ (_13863_, _13849_, _13814_);
  or _65409_ (_40749_, _13863_, _13862_);
  or _65410_ (_13864_, _13845_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _65411_ (_13865_, _13864_, _13850_);
  or _65412_ (_13866_, _13846_, _13443_);
  and _65413_ (_13867_, _13866_, _13865_);
  and _65414_ (_13868_, _13849_, _13820_);
  or _65415_ (_40750_, _13868_, _13867_);
  or _65416_ (_13869_, _13846_, _13450_);
  or _65417_ (_13870_, _13845_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _65418_ (_13871_, _13870_, _13850_);
  and _65419_ (_13872_, _13871_, _13869_);
  and _65420_ (_13873_, _13849_, _13826_);
  or _65421_ (_40751_, _13873_, _13872_);
  or _65422_ (_13874_, _13845_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _65423_ (_13875_, _13874_, _13850_);
  or _65424_ (_13876_, _13846_, _13202_);
  and _65425_ (_13877_, _13876_, _13875_);
  and _65426_ (_13878_, _13849_, _13832_);
  or _65427_ (_40753_, _13878_, _13877_);
  or _65428_ (_13879_, _13845_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _65429_ (_13880_, _13879_, _13850_);
  or _65430_ (_13881_, _13846_, _13462_);
  and _65431_ (_13882_, _13881_, _13880_);
  and _65432_ (_13883_, _13849_, _13838_);
  or _65433_ (_40754_, _13883_, _13882_);
  or _65434_ (_13884_, _13845_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _65435_ (_13885_, _13884_, _13850_);
  or _65436_ (_13886_, _13846_, _06800_);
  and _65437_ (_13887_, _13886_, _13885_);
  and _65438_ (_13888_, _13849_, _06824_);
  or _65439_ (_40755_, _13888_, _13887_);
  and _65440_ (_13889_, _13794_, _13471_);
  not _65441_ (_13890_, _13889_);
  or _65442_ (_13891_, _13890_, _12171_);
  or _65443_ (_13892_, _13889_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _65444_ (_13893_, _13798_, _05967_);
  not _65445_ (_13894_, _13893_);
  and _65446_ (_13895_, _13894_, _13892_);
  and _65447_ (_13896_, _13895_, _13891_);
  and _65448_ (_13897_, _13893_, _13480_);
  or _65449_ (_40759_, _13897_, _13896_);
  or _65450_ (_13898_, _13889_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _65451_ (_13899_, _13898_, _13894_);
  or _65452_ (_13900_, _13890_, _12388_);
  and _65453_ (_13901_, _13900_, _13899_);
  and _65454_ (_13902_, _13893_, _13486_);
  or _65455_ (_40760_, _13902_, _13901_);
  or _65456_ (_13903_, _13889_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _65457_ (_13904_, _13903_, _13894_);
  or _65458_ (_13905_, _13890_, _13436_);
  and _65459_ (_13906_, _13905_, _13904_);
  and _65460_ (_13907_, _13893_, _13814_);
  or _65461_ (_40761_, _13907_, _13906_);
  or _65462_ (_13908_, _13889_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _65463_ (_13909_, _13908_, _13894_);
  or _65464_ (_13910_, _13890_, _13443_);
  and _65465_ (_13911_, _13910_, _13909_);
  and _65466_ (_13912_, _13893_, _13820_);
  or _65467_ (_40762_, _13912_, _13911_);
  or _65468_ (_13913_, _13889_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _65469_ (_13914_, _13913_, _13894_);
  or _65470_ (_13915_, _13890_, _13450_);
  and _65471_ (_13916_, _13915_, _13914_);
  and _65472_ (_13917_, _13893_, _13826_);
  or _65473_ (_40764_, _13917_, _13916_);
  or _65474_ (_13918_, _13889_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _65475_ (_13919_, _13918_, _13894_);
  or _65476_ (_13920_, _13890_, _13202_);
  and _65477_ (_13921_, _13920_, _13919_);
  and _65478_ (_13922_, _13893_, _13832_);
  or _65479_ (_40765_, _13922_, _13921_);
  or _65480_ (_13923_, _13889_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _65481_ (_13924_, _13923_, _13894_);
  or _65482_ (_13925_, _13890_, _13462_);
  and _65483_ (_13926_, _13925_, _13924_);
  and _65484_ (_13927_, _13893_, _13838_);
  or _65485_ (_40766_, _13927_, _13926_);
  or _65486_ (_13928_, _13889_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _65487_ (_13929_, _13928_, _13894_);
  or _65488_ (_13930_, _13890_, _06800_);
  and _65489_ (_13931_, _13930_, _13929_);
  and _65490_ (_13932_, _13893_, _06824_);
  or _65491_ (_40767_, _13932_, _13931_);
  and _65492_ (_13933_, _13794_, _04799_);
  not _65493_ (_13934_, _13933_);
  or _65494_ (_13935_, _13934_, _12171_);
  and _65495_ (_13936_, _13798_, _03497_);
  not _65496_ (_13937_, _13936_);
  or _65497_ (_13938_, _13933_, \oc8051_golden_model_1.IRAM[11] [0]);
  and _65498_ (_13939_, _13938_, _13937_);
  and _65499_ (_13940_, _13939_, _13935_);
  and _65500_ (_13941_, _13936_, _13480_);
  or _65501_ (_40771_, _13941_, _13940_);
  or _65502_ (_13942_, _13934_, _12388_);
  or _65503_ (_13943_, _13933_, \oc8051_golden_model_1.IRAM[11] [1]);
  and _65504_ (_13944_, _13943_, _13937_);
  and _65505_ (_13945_, _13944_, _13942_);
  and _65506_ (_13946_, _13936_, _13486_);
  or _65507_ (_40772_, _13946_, _13945_);
  or _65508_ (_13947_, _13933_, \oc8051_golden_model_1.IRAM[11] [2]);
  and _65509_ (_13948_, _13947_, _13937_);
  or _65510_ (_13949_, _13934_, _13436_);
  and _65511_ (_13950_, _13949_, _13948_);
  and _65512_ (_13951_, _13936_, _13814_);
  or _65513_ (_40773_, _13951_, _13950_);
  or _65514_ (_13952_, _13934_, _13443_);
  or _65515_ (_13953_, _13933_, \oc8051_golden_model_1.IRAM[11] [3]);
  and _65516_ (_13954_, _13953_, _13937_);
  and _65517_ (_13955_, _13954_, _13952_);
  and _65518_ (_13956_, _13936_, _13820_);
  or _65519_ (_40774_, _13956_, _13955_);
  or _65520_ (_13957_, _13934_, _13450_);
  or _65521_ (_13958_, _13933_, \oc8051_golden_model_1.IRAM[11] [4]);
  and _65522_ (_13959_, _13958_, _13937_);
  and _65523_ (_13960_, _13959_, _13957_);
  and _65524_ (_13961_, _13936_, _13826_);
  or _65525_ (_40776_, _13961_, _13960_);
  or _65526_ (_13962_, _13934_, _13202_);
  or _65527_ (_13963_, _13933_, \oc8051_golden_model_1.IRAM[11] [5]);
  and _65528_ (_13964_, _13963_, _13937_);
  and _65529_ (_13965_, _13964_, _13962_);
  and _65530_ (_13966_, _13936_, _13832_);
  or _65531_ (_40777_, _13966_, _13965_);
  or _65532_ (_13967_, _13934_, _13462_);
  or _65533_ (_13968_, _13933_, \oc8051_golden_model_1.IRAM[11] [6]);
  and _65534_ (_13969_, _13968_, _13937_);
  and _65535_ (_13970_, _13969_, _13967_);
  and _65536_ (_13971_, _13936_, _13838_);
  or _65537_ (_40778_, _13971_, _13970_);
  or _65538_ (_13972_, _13934_, _06800_);
  or _65539_ (_13973_, _13933_, \oc8051_golden_model_1.IRAM[11] [7]);
  and _65540_ (_13974_, _13973_, _13937_);
  and _65541_ (_13975_, _13974_, _13972_);
  and _65542_ (_13976_, _13936_, _06824_);
  or _65543_ (_40779_, _13976_, _13975_);
  and _65544_ (_13977_, _11994_, _05124_);
  not _65545_ (_13978_, _13977_);
  or _65546_ (_13979_, _13978_, _12171_);
  and _65547_ (_13980_, _05139_, _03499_);
  not _65548_ (_13981_, _13980_);
  or _65549_ (_13982_, _13977_, \oc8051_golden_model_1.IRAM[12] [0]);
  and _65550_ (_13983_, _13982_, _13981_);
  and _65551_ (_13984_, _13983_, _13979_);
  and _65552_ (_13985_, _13980_, _13480_);
  or _65553_ (_40783_, _13985_, _13984_);
  or _65554_ (_13986_, _13977_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _65555_ (_13987_, _13986_, _13981_);
  or _65556_ (_13988_, _13978_, _12388_);
  and _65557_ (_13989_, _13988_, _13987_);
  and _65558_ (_13990_, _13980_, _13486_);
  or _65559_ (_40784_, _13990_, _13989_);
  or _65560_ (_13991_, _13977_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _65561_ (_13992_, _13991_, _13981_);
  or _65562_ (_13993_, _13978_, _13436_);
  and _65563_ (_13994_, _13993_, _13992_);
  and _65564_ (_13995_, _13980_, _13814_);
  or _65565_ (_40786_, _13995_, _13994_);
  or _65566_ (_13996_, _13977_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _65567_ (_13997_, _13996_, _13981_);
  or _65568_ (_13998_, _13978_, _13443_);
  and _65569_ (_13999_, _13998_, _13997_);
  and _65570_ (_14000_, _13980_, _13820_);
  or _65571_ (_40787_, _14000_, _13999_);
  or _65572_ (_14001_, _13977_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _65573_ (_14002_, _14001_, _13981_);
  or _65574_ (_14003_, _13978_, _13450_);
  and _65575_ (_14004_, _14003_, _14002_);
  and _65576_ (_14005_, _13980_, _13826_);
  or _65577_ (_40788_, _14005_, _14004_);
  or _65578_ (_14006_, _13977_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _65579_ (_14007_, _14006_, _13981_);
  or _65580_ (_14008_, _13978_, _13202_);
  and _65581_ (_14009_, _14008_, _14007_);
  and _65582_ (_14010_, _13980_, _13832_);
  or _65583_ (_40789_, _14010_, _14009_);
  or _65584_ (_14011_, _13977_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _65585_ (_14012_, _14011_, _13981_);
  or _65586_ (_14013_, _13978_, _13462_);
  and _65587_ (_14014_, _14013_, _14012_);
  and _65588_ (_14015_, _13980_, _13838_);
  or _65589_ (_40790_, _14015_, _14014_);
  or _65590_ (_14016_, _13977_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _65591_ (_14017_, _14016_, _13981_);
  or _65592_ (_14018_, _13978_, _06800_);
  and _65593_ (_14019_, _14018_, _14017_);
  and _65594_ (_14020_, _13980_, _06824_);
  or _65595_ (_40792_, _14020_, _14019_);
  and _65596_ (_14021_, _13417_, _05124_);
  not _65597_ (_14022_, _14021_);
  or _65598_ (_14023_, _14022_, _12171_);
  or _65599_ (_14024_, _14021_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _65600_ (_14025_, _05139_, _04804_);
  not _65601_ (_14026_, _14025_);
  and _65602_ (_14027_, _14026_, _14024_);
  and _65603_ (_14028_, _14027_, _14023_);
  and _65604_ (_14029_, _14025_, _13480_);
  or _65605_ (_40795_, _14029_, _14028_);
  or _65606_ (_14030_, _14021_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _65607_ (_14031_, _14030_, _14026_);
  or _65608_ (_14032_, _14022_, _12388_);
  and _65609_ (_14033_, _14032_, _14031_);
  and _65610_ (_14034_, _14025_, _13486_);
  or _65611_ (_40796_, _14034_, _14033_);
  or _65612_ (_14035_, _14021_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _65613_ (_14036_, _14035_, _14026_);
  or _65614_ (_14037_, _14022_, _13436_);
  and _65615_ (_14038_, _14037_, _14036_);
  and _65616_ (_14039_, _14025_, _13814_);
  or _65617_ (_40798_, _14039_, _14038_);
  or _65618_ (_14040_, _14021_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _65619_ (_14041_, _14040_, _14026_);
  or _65620_ (_14042_, _14022_, _13443_);
  and _65621_ (_14043_, _14042_, _14041_);
  and _65622_ (_14044_, _14025_, _13820_);
  or _65623_ (_40799_, _14044_, _14043_);
  or _65624_ (_14045_, _14021_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _65625_ (_14046_, _14045_, _14026_);
  or _65626_ (_14047_, _14022_, _13450_);
  and _65627_ (_14048_, _14047_, _14046_);
  and _65628_ (_14049_, _14025_, _13826_);
  or _65629_ (_40800_, _14049_, _14048_);
  or _65630_ (_14050_, _14021_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _65631_ (_14051_, _14050_, _14026_);
  or _65632_ (_14052_, _14022_, _13202_);
  and _65633_ (_14053_, _14052_, _14051_);
  and _65634_ (_14054_, _14025_, _13832_);
  or _65635_ (_40801_, _14054_, _14053_);
  or _65636_ (_14055_, _14021_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _65637_ (_14056_, _14055_, _14026_);
  or _65638_ (_14057_, _14022_, _13462_);
  and _65639_ (_14058_, _14057_, _14056_);
  and _65640_ (_14059_, _14025_, _13838_);
  or _65641_ (_40802_, _14059_, _14058_);
  nor _65642_ (_14060_, _14021_, \oc8051_golden_model_1.IRAM[13] [7]);
  nor _65643_ (_14061_, _14022_, _06800_);
  or _65644_ (_14062_, _14061_, _14060_);
  nand _65645_ (_14063_, _14062_, _14026_);
  or _65646_ (_14064_, _14026_, _06824_);
  and _65647_ (_40804_, _14064_, _14063_);
  and _65648_ (_14065_, _13471_, _05124_);
  not _65649_ (_14066_, _14065_);
  or _65650_ (_14067_, _14066_, _12171_);
  or _65651_ (_14068_, _14065_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _65652_ (_14069_, _05967_, _05139_);
  not _65653_ (_14070_, _14069_);
  and _65654_ (_14071_, _14070_, _14068_);
  and _65655_ (_14072_, _14071_, _14067_);
  and _65656_ (_14073_, _14069_, _13480_);
  or _65657_ (_40807_, _14073_, _14072_);
  or _65658_ (_14074_, _14066_, _12388_);
  or _65659_ (_14075_, _14065_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _65660_ (_14076_, _14075_, _14070_);
  and _65661_ (_14077_, _14076_, _14074_);
  and _65662_ (_14078_, _14069_, _13486_);
  or _65663_ (_40809_, _14078_, _14077_);
  or _65664_ (_14079_, _14065_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _65665_ (_14080_, _14079_, _14070_);
  or _65666_ (_14081_, _14066_, _13436_);
  and _65667_ (_14082_, _14081_, _14080_);
  and _65668_ (_14083_, _14069_, _13814_);
  or _65669_ (_40810_, _14083_, _14082_);
  or _65670_ (_14084_, _14065_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _65671_ (_14085_, _14084_, _14070_);
  or _65672_ (_14086_, _14066_, _13443_);
  and _65673_ (_14087_, _14086_, _14085_);
  and _65674_ (_14088_, _14069_, _13820_);
  or _65675_ (_40811_, _14088_, _14087_);
  or _65676_ (_14089_, _14065_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _65677_ (_14090_, _14089_, _14070_);
  or _65678_ (_14091_, _14066_, _13450_);
  and _65679_ (_14092_, _14091_, _14090_);
  and _65680_ (_14093_, _14069_, _13826_);
  or _65681_ (_40812_, _14093_, _14092_);
  or _65682_ (_14094_, _14065_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _65683_ (_14095_, _14094_, _14070_);
  or _65684_ (_14096_, _14066_, _13202_);
  and _65685_ (_14097_, _14096_, _14095_);
  and _65686_ (_14098_, _14069_, _13832_);
  or _65687_ (_40813_, _14098_, _14097_);
  or _65688_ (_14099_, _14065_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _65689_ (_14100_, _14099_, _14070_);
  or _65690_ (_14101_, _14066_, _13462_);
  and _65691_ (_14102_, _14101_, _14100_);
  and _65692_ (_14103_, _14069_, _13838_);
  or _65693_ (_40815_, _14103_, _14102_);
  or _65694_ (_14104_, _14065_, \oc8051_golden_model_1.IRAM[14] [7]);
  and _65695_ (_14105_, _14104_, _14070_);
  or _65696_ (_14106_, _14066_, _06800_);
  and _65697_ (_14107_, _14106_, _14105_);
  and _65698_ (_14108_, _14069_, _06824_);
  or _65699_ (_40816_, _14108_, _14107_);
  or _65700_ (_14109_, _12171_, _05143_);
  or _65701_ (_14110_, _05125_, \oc8051_golden_model_1.IRAM[15] [0]);
  and _65702_ (_14111_, _14110_, _05141_);
  and _65703_ (_14112_, _14111_, _14109_);
  and _65704_ (_14113_, _13480_, _05140_);
  or _65705_ (_40819_, _14113_, _14112_);
  or _65706_ (_14114_, _05125_, \oc8051_golden_model_1.IRAM[15] [1]);
  and _65707_ (_14115_, _14114_, _05141_);
  or _65708_ (_14116_, _12388_, _05143_);
  and _65709_ (_14117_, _14116_, _14115_);
  and _65710_ (_14118_, _13486_, _05140_);
  or _65711_ (_40821_, _14118_, _14117_);
  or _65712_ (_14119_, _05125_, \oc8051_golden_model_1.IRAM[15] [2]);
  and _65713_ (_14120_, _14119_, _05141_);
  or _65714_ (_14121_, _13436_, _05143_);
  and _65715_ (_14122_, _14121_, _14120_);
  and _65716_ (_14123_, _13814_, _05140_);
  or _65717_ (_40822_, _14123_, _14122_);
  or _65718_ (_14124_, _05125_, \oc8051_golden_model_1.IRAM[15] [3]);
  and _65719_ (_14125_, _14124_, _05141_);
  or _65720_ (_14126_, _13443_, _05143_);
  and _65721_ (_14127_, _14126_, _14125_);
  and _65722_ (_14128_, _13820_, _05140_);
  or _65723_ (_40823_, _14128_, _14127_);
  or _65724_ (_14129_, _05125_, \oc8051_golden_model_1.IRAM[15] [4]);
  and _65725_ (_14130_, _14129_, _05141_);
  or _65726_ (_14131_, _13450_, _05143_);
  and _65727_ (_14132_, _14131_, _14130_);
  and _65728_ (_14133_, _13826_, _05140_);
  or _65729_ (_40824_, _14133_, _14132_);
  or _65730_ (_14134_, _05125_, \oc8051_golden_model_1.IRAM[15] [5]);
  and _65731_ (_14135_, _14134_, _05141_);
  or _65732_ (_14136_, _13202_, _05143_);
  and _65733_ (_14137_, _14136_, _14135_);
  and _65734_ (_14138_, _13832_, _05140_);
  or _65735_ (_40825_, _14138_, _14137_);
  or _65736_ (_14139_, _05125_, \oc8051_golden_model_1.IRAM[15] [6]);
  and _65737_ (_14140_, _14139_, _05141_);
  or _65738_ (_14141_, _13462_, _05143_);
  and _65739_ (_14142_, _14141_, _14140_);
  and _65740_ (_14143_, _13838_, _05140_);
  or _65741_ (_40827_, _14143_, _14142_);
  nor _65742_ (_14144_, _43000_, _07418_);
  nor _65743_ (_14145_, _05248_, _07418_);
  and _65744_ (_14146_, _12128_, _05248_);
  or _65745_ (_14147_, _14146_, _14145_);
  and _65746_ (_14148_, _14147_, _03780_);
  nor _65747_ (_14149_, _05666_, _06830_);
  or _65748_ (_14150_, _14149_, _14145_);
  or _65749_ (_14151_, _14150_, _04081_);
  and _65750_ (_14152_, _05248_, \oc8051_golden_model_1.ACC [0]);
  or _65751_ (_14153_, _14152_, _14145_);
  and _65752_ (_14154_, _14153_, _04409_);
  nor _65753_ (_14155_, _04409_, _07418_);
  or _65754_ (_14156_, _14155_, _03610_);
  or _65755_ (_14157_, _14156_, _14154_);
  and _65756_ (_14158_, _14157_, _04055_);
  and _65757_ (_14159_, _14158_, _14151_);
  and _65758_ (_14160_, _12021_, _05910_);
  nor _65759_ (_14161_, _05910_, _07418_);
  or _65760_ (_14162_, _14161_, _14160_);
  and _65761_ (_14163_, _14162_, _03715_);
  or _65762_ (_14164_, _14163_, _14159_);
  and _65763_ (_14165_, _14164_, _03996_);
  and _65764_ (_14166_, _05248_, _04620_);
  or _65765_ (_14167_, _14166_, _14145_);
  and _65766_ (_14168_, _14167_, _03723_);
  or _65767_ (_14169_, _14168_, _03729_);
  or _65768_ (_14170_, _14169_, _14165_);
  or _65769_ (_14171_, _14153_, _03737_);
  and _65770_ (_14172_, _14171_, _03736_);
  and _65771_ (_14173_, _14172_, _14170_);
  and _65772_ (_14174_, _14145_, _03714_);
  or _65773_ (_14175_, _14174_, _03719_);
  or _65774_ (_14176_, _14175_, _14173_);
  or _65775_ (_14177_, _14150_, _06840_);
  and _65776_ (_14178_, _14177_, _14176_);
  or _65777_ (_14179_, _14178_, _06869_);
  nor _65778_ (_14180_, _07351_, _07349_);
  nor _65779_ (_14181_, _14180_, _07352_);
  or _65780_ (_14182_, _14181_, _06875_);
  and _65781_ (_14183_, _14182_, _03710_);
  and _65782_ (_14184_, _14183_, _14179_);
  nor _65783_ (_14185_, _12052_, _07391_);
  or _65784_ (_14186_, _14185_, _14161_);
  and _65785_ (_14187_, _14186_, _03505_);
  or _65786_ (_14188_, _14187_, _07390_);
  or _65787_ (_14189_, _14188_, _14184_);
  or _65788_ (_14190_, _14167_, _06838_);
  and _65789_ (_14191_, _14190_, _07400_);
  and _65790_ (_14192_, _14191_, _14189_);
  and _65791_ (_14193_, _06546_, _05248_);
  or _65792_ (_14194_, _14193_, _14145_);
  and _65793_ (_14195_, _14194_, _04481_);
  or _65794_ (_14196_, _14195_, _03222_);
  or _65795_ (_14197_, _14196_, _14192_);
  nor _65796_ (_14198_, _12109_, _06830_);
  or _65797_ (_14199_, _14145_, _03589_);
  or _65798_ (_14200_, _14199_, _14198_);
  and _65799_ (_14201_, _14200_, _07411_);
  and _65800_ (_14202_, _14201_, _14197_);
  nor _65801_ (_14203_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor _65802_ (_14204_, _14203_, _07330_);
  or _65803_ (_14205_, _07760_, _14204_);
  nand _65804_ (_14206_, _07760_, _03335_);
  and _65805_ (_14207_, _14206_, _07405_);
  and _65806_ (_14208_, _14207_, _14205_);
  or _65807_ (_14209_, _14208_, _08828_);
  or _65808_ (_14210_, _14209_, _14202_);
  and _65809_ (_14211_, _12124_, _05248_);
  or _65810_ (_14212_, _14145_, _07766_);
  or _65811_ (_14213_, _14212_, _14211_);
  and _65812_ (_14214_, _05248_, _06274_);
  or _65813_ (_14215_, _14214_, _14145_);
  or _65814_ (_14216_, _14215_, _05886_);
  and _65815_ (_14217_, _14216_, _07778_);
  and _65816_ (_14218_, _14217_, _14213_);
  and _65817_ (_14219_, _14218_, _14210_);
  or _65818_ (_14220_, _14219_, _14148_);
  and _65819_ (_14221_, _14220_, _07777_);
  nand _65820_ (_14222_, _14215_, _03622_);
  nor _65821_ (_14223_, _14222_, _14149_);
  or _65822_ (_14224_, _14223_, _14221_);
  and _65823_ (_14225_, _14224_, _06828_);
  or _65824_ (_14226_, _14145_, _05666_);
  and _65825_ (_14227_, _14153_, _03790_);
  and _65826_ (_14228_, _14227_, _14226_);
  or _65827_ (_14229_, _14228_, _03624_);
  or _65828_ (_14230_, _14229_, _14225_);
  nor _65829_ (_14231_, _12122_, _06830_);
  or _65830_ (_14232_, _14145_, _07795_);
  or _65831_ (_14233_, _14232_, _14231_);
  and _65832_ (_14234_, _14233_, _07793_);
  and _65833_ (_14235_, _14234_, _14230_);
  nor _65834_ (_14236_, _12003_, _06830_);
  or _65835_ (_14237_, _14236_, _14145_);
  and _65836_ (_14238_, _14237_, _03785_);
  or _65837_ (_14239_, _14238_, _03815_);
  or _65838_ (_14240_, _14239_, _14235_);
  or _65839_ (_14241_, _14150_, _04246_);
  and _65840_ (_14242_, _14241_, _03823_);
  and _65841_ (_14243_, _14242_, _14240_);
  and _65842_ (_14244_, _14145_, _03453_);
  or _65843_ (_14245_, _14244_, _03447_);
  or _65844_ (_14246_, _14245_, _14243_);
  or _65845_ (_14247_, _14150_, _03514_);
  and _65846_ (_14248_, _14247_, _43000_);
  and _65847_ (_14249_, _14248_, _14246_);
  or _65848_ (_14250_, _14249_, _14144_);
  and _65849_ (_43480_, _14250_, _41806_);
  nor _65850_ (_14251_, _43000_, _07412_);
  or _65851_ (_14252_, _05248_, \oc8051_golden_model_1.B [1]);
  and _65852_ (_14253_, _12213_, _05248_);
  not _65853_ (_14254_, _14253_);
  and _65854_ (_14255_, _14254_, _14252_);
  or _65855_ (_14256_, _14255_, _04081_);
  nand _65856_ (_14257_, _05248_, _03274_);
  and _65857_ (_14258_, _14257_, _14252_);
  and _65858_ (_14259_, _14258_, _04409_);
  nor _65859_ (_14260_, _04409_, _07412_);
  or _65860_ (_14261_, _14260_, _03610_);
  or _65861_ (_14262_, _14261_, _14259_);
  and _65862_ (_14263_, _14262_, _04055_);
  and _65863_ (_14264_, _14263_, _14256_);
  not _65864_ (_14265_, _03730_);
  and _65865_ (_14266_, _12224_, _05910_);
  nor _65866_ (_14267_, _05910_, _07412_);
  or _65867_ (_14268_, _14267_, _03723_);
  or _65868_ (_14269_, _14268_, _14266_);
  and _65869_ (_14270_, _14269_, _14265_);
  or _65870_ (_14271_, _14270_, _14264_);
  nor _65871_ (_14272_, _05248_, _07412_);
  and _65872_ (_14273_, _05248_, _06764_);
  or _65873_ (_14274_, _14273_, _14272_);
  or _65874_ (_14275_, _14274_, _03996_);
  and _65875_ (_14276_, _14275_, _14271_);
  or _65876_ (_14277_, _14276_, _03729_);
  or _65877_ (_14278_, _14258_, _03737_);
  and _65878_ (_14279_, _14278_, _03736_);
  and _65879_ (_14280_, _14279_, _14277_);
  and _65880_ (_14281_, _12211_, _05910_);
  or _65881_ (_14282_, _14281_, _14267_);
  and _65882_ (_14283_, _14282_, _03714_);
  or _65883_ (_14284_, _14283_, _14280_);
  and _65884_ (_14285_, _14284_, _06840_);
  and _65885_ (_14286_, _14266_, _12239_);
  or _65886_ (_14287_, _14286_, _14267_);
  and _65887_ (_14288_, _14287_, _03719_);
  or _65888_ (_14289_, _14288_, _06869_);
  or _65889_ (_14290_, _14289_, _14285_);
  or _65890_ (_14291_, _07296_, _07295_);
  nand _65891_ (_14292_, _14291_, _07353_);
  or _65892_ (_14293_, _14291_, _07353_);
  and _65893_ (_14294_, _14293_, _14292_);
  or _65894_ (_14295_, _14294_, _06875_);
  and _65895_ (_14296_, _14295_, _03710_);
  and _65896_ (_14297_, _14296_, _14290_);
  nor _65897_ (_14298_, _12256_, _07391_);
  or _65898_ (_14299_, _14298_, _14267_);
  and _65899_ (_14300_, _14299_, _03505_);
  or _65900_ (_14301_, _14300_, _07390_);
  or _65901_ (_14302_, _14301_, _14297_);
  or _65902_ (_14303_, _14274_, _06838_);
  and _65903_ (_14304_, _14303_, _14302_);
  or _65904_ (_14305_, _14304_, _04481_);
  and _65905_ (_14306_, _06501_, _05248_);
  or _65906_ (_14307_, _14272_, _07400_);
  or _65907_ (_14308_, _14307_, _14306_);
  and _65908_ (_14309_, _14308_, _03589_);
  and _65909_ (_14310_, _14309_, _14305_);
  nand _65910_ (_14311_, _12313_, _05248_);
  and _65911_ (_14312_, _14252_, _03222_);
  and _65912_ (_14313_, _14312_, _14311_);
  or _65913_ (_14314_, _14313_, _07405_);
  or _65914_ (_14315_, _14314_, _14310_);
  and _65915_ (_14316_, _07760_, _07707_);
  nor _65916_ (_14317_, _07755_, _07754_);
  or _65917_ (_14318_, _14317_, _07756_);
  nor _65918_ (_14319_, _14318_, _07760_);
  or _65919_ (_14320_, _14319_, _14316_);
  or _65920_ (_14321_, _14320_, _07411_);
  and _65921_ (_14322_, _14321_, _05886_);
  and _65922_ (_14323_, _14322_, _14315_);
  nand _65923_ (_14324_, _05248_, _04303_);
  and _65924_ (_14325_, _14324_, _03601_);
  and _65925_ (_14326_, _14325_, _14252_);
  or _65926_ (_14327_, _14326_, _14323_);
  and _65927_ (_14328_, _14327_, _07766_);
  or _65928_ (_14329_, _12327_, _06830_);
  and _65929_ (_14330_, _14252_, _03600_);
  and _65930_ (_14331_, _14330_, _14329_);
  or _65931_ (_14332_, _14331_, _14328_);
  and _65932_ (_14333_, _14332_, _07778_);
  or _65933_ (_14334_, _12333_, _06830_);
  and _65934_ (_14335_, _14252_, _03780_);
  and _65935_ (_14336_, _14335_, _14334_);
  or _65936_ (_14337_, _14336_, _14333_);
  and _65937_ (_14338_, _14337_, _07777_);
  or _65938_ (_14339_, _12207_, _06830_);
  and _65939_ (_14340_, _14252_, _03622_);
  and _65940_ (_14341_, _14340_, _14339_);
  or _65941_ (_14342_, _14341_, _14338_);
  and _65942_ (_14343_, _14342_, _06828_);
  or _65943_ (_14344_, _14272_, _05618_);
  and _65944_ (_14345_, _14258_, _03790_);
  and _65945_ (_14346_, _14345_, _14344_);
  or _65946_ (_14347_, _14346_, _14343_);
  and _65947_ (_14348_, _14347_, _03786_);
  or _65948_ (_14349_, _14324_, _05618_);
  and _65949_ (_14350_, _14252_, _03624_);
  and _65950_ (_14351_, _14350_, _14349_);
  or _65951_ (_14352_, _14257_, _05618_);
  and _65952_ (_14353_, _14252_, _03785_);
  and _65953_ (_14354_, _14353_, _14352_);
  or _65954_ (_14355_, _14354_, _03815_);
  or _65955_ (_14356_, _14355_, _14351_);
  or _65956_ (_14357_, _14356_, _14348_);
  or _65957_ (_14358_, _14255_, _04246_);
  and _65958_ (_14359_, _14358_, _03823_);
  and _65959_ (_14360_, _14359_, _14357_);
  and _65960_ (_14361_, _14282_, _03453_);
  or _65961_ (_14362_, _14361_, _03447_);
  or _65962_ (_14363_, _14362_, _14360_);
  or _65963_ (_14364_, _14272_, _03514_);
  or _65964_ (_14365_, _14364_, _14253_);
  and _65965_ (_14366_, _14365_, _43000_);
  and _65966_ (_14367_, _14366_, _14363_);
  or _65967_ (_14368_, _14367_, _14251_);
  and _65968_ (_43481_, _14368_, _41806_);
  nor _65969_ (_14369_, _43000_, _07426_);
  nor _65970_ (_14370_, _05248_, _07426_);
  nor _65971_ (_14371_, _06830_, _04875_);
  or _65972_ (_14372_, _14371_, _14370_);
  or _65973_ (_14373_, _14372_, _06838_);
  and _65974_ (_14374_, _12411_, _05910_);
  and _65975_ (_14375_, _14374_, _12443_);
  nor _65976_ (_14376_, _05910_, _07426_);
  or _65977_ (_14377_, _14376_, _06840_);
  or _65978_ (_14378_, _14377_, _14375_);
  or _65979_ (_14379_, _14372_, _03996_);
  nor _65980_ (_14380_, _12416_, _06830_);
  or _65981_ (_14381_, _14380_, _14370_);
  or _65982_ (_14382_, _14381_, _04081_);
  and _65983_ (_14383_, _05248_, \oc8051_golden_model_1.ACC [2]);
  or _65984_ (_14384_, _14383_, _14370_);
  and _65985_ (_14385_, _14384_, _04409_);
  nor _65986_ (_14386_, _04409_, _07426_);
  or _65987_ (_14387_, _14386_, _03610_);
  or _65988_ (_14388_, _14387_, _14385_);
  and _65989_ (_14389_, _14388_, _04055_);
  and _65990_ (_14390_, _14389_, _14382_);
  or _65991_ (_14391_, _14376_, _14374_);
  and _65992_ (_14392_, _14391_, _03715_);
  or _65993_ (_14393_, _14392_, _03723_);
  or _65994_ (_14394_, _14393_, _14390_);
  and _65995_ (_14395_, _14394_, _14379_);
  or _65996_ (_14396_, _14395_, _03729_);
  or _65997_ (_14397_, _14384_, _03737_);
  and _65998_ (_14398_, _14397_, _03736_);
  and _65999_ (_14399_, _14398_, _14396_);
  and _66000_ (_14400_, _12409_, _05910_);
  or _66001_ (_14401_, _14400_, _14376_);
  and _66002_ (_14402_, _14401_, _03714_);
  or _66003_ (_14403_, _14402_, _03719_);
  or _66004_ (_14404_, _14403_, _14399_);
  and _66005_ (_14405_, _14404_, _14378_);
  or _66006_ (_14406_, _14405_, _06869_);
  nor _66007_ (_14407_, _07355_, _07252_);
  nor _66008_ (_14408_, _14407_, _07356_);
  or _66009_ (_14409_, _14408_, _06875_);
  and _66010_ (_14410_, _14409_, _03710_);
  and _66011_ (_14411_, _14410_, _14406_);
  nor _66012_ (_14412_, _12461_, _07391_);
  or _66013_ (_14413_, _14412_, _14376_);
  and _66014_ (_14414_, _14413_, _03505_);
  or _66015_ (_14415_, _14414_, _07390_);
  or _66016_ (_14416_, _14415_, _14411_);
  and _66017_ (_14417_, _14416_, _14373_);
  or _66018_ (_14418_, _14417_, _04481_);
  and _66019_ (_14419_, _06637_, _05248_);
  or _66020_ (_14420_, _14370_, _07400_);
  or _66021_ (_14421_, _14420_, _14419_);
  and _66022_ (_14422_, _14421_, _14418_);
  or _66023_ (_14423_, _14422_, _03222_);
  nor _66024_ (_14424_, _12519_, _06830_);
  or _66025_ (_14425_, _14370_, _03589_);
  or _66026_ (_14426_, _14425_, _14424_);
  and _66027_ (_14427_, _14426_, _07411_);
  and _66028_ (_14428_, _14427_, _14423_);
  not _66029_ (_14429_, _07760_);
  or _66030_ (_14430_, _14429_, _07697_);
  nor _66031_ (_14431_, _07756_, _07708_);
  not _66032_ (_14432_, _14431_);
  and _66033_ (_14433_, _14432_, _07700_);
  nor _66034_ (_14434_, _14432_, _07700_);
  nor _66035_ (_14435_, _14434_, _14433_);
  or _66036_ (_14436_, _14435_, _07760_);
  and _66037_ (_14437_, _14436_, _07405_);
  and _66038_ (_14438_, _14437_, _14430_);
  or _66039_ (_14439_, _14438_, _08828_);
  or _66040_ (_14440_, _14439_, _14428_);
  and _66041_ (_14441_, _12533_, _05248_);
  or _66042_ (_14442_, _14370_, _07766_);
  or _66043_ (_14443_, _14442_, _14441_);
  and _66044_ (_14444_, _05248_, _06332_);
  or _66045_ (_14445_, _14444_, _14370_);
  or _66046_ (_14446_, _14445_, _05886_);
  and _66047_ (_14447_, _14446_, _07778_);
  and _66048_ (_14448_, _14447_, _14443_);
  and _66049_ (_14449_, _14448_, _14440_);
  and _66050_ (_14450_, _12539_, _05248_);
  or _66051_ (_14451_, _14450_, _14370_);
  and _66052_ (_14452_, _14451_, _03780_);
  or _66053_ (_14453_, _14452_, _14449_);
  and _66054_ (_14454_, _14453_, _07777_);
  or _66055_ (_14455_, _14370_, _05718_);
  and _66056_ (_14456_, _14445_, _03622_);
  and _66057_ (_14457_, _14456_, _14455_);
  or _66058_ (_14458_, _14457_, _14454_);
  and _66059_ (_14459_, _14458_, _06828_);
  and _66060_ (_14460_, _14384_, _03790_);
  and _66061_ (_14461_, _14460_, _14455_);
  or _66062_ (_14462_, _14461_, _03624_);
  or _66063_ (_14463_, _14462_, _14459_);
  nor _66064_ (_14464_, _12532_, _06830_);
  or _66065_ (_14465_, _14370_, _07795_);
  or _66066_ (_14466_, _14465_, _14464_);
  and _66067_ (_14467_, _14466_, _07793_);
  and _66068_ (_14468_, _14467_, _14463_);
  nor _66069_ (_14469_, _12538_, _06830_);
  or _66070_ (_14470_, _14469_, _14370_);
  and _66071_ (_14471_, _14470_, _03785_);
  or _66072_ (_14472_, _14471_, _03815_);
  or _66073_ (_14473_, _14472_, _14468_);
  or _66074_ (_14474_, _14381_, _04246_);
  and _66075_ (_14475_, _14474_, _03823_);
  and _66076_ (_14476_, _14475_, _14473_);
  and _66077_ (_14477_, _14401_, _03453_);
  or _66078_ (_14478_, _14477_, _03447_);
  or _66079_ (_14479_, _14478_, _14476_);
  and _66080_ (_14480_, _12592_, _05248_);
  or _66081_ (_14481_, _14370_, _03514_);
  or _66082_ (_14482_, _14481_, _14480_);
  and _66083_ (_14483_, _14482_, _43000_);
  and _66084_ (_14484_, _14483_, _14479_);
  or _66085_ (_14485_, _14484_, _14369_);
  and _66086_ (_43482_, _14485_, _41806_);
  nor _66087_ (_14486_, _43000_, _07427_);
  nor _66088_ (_14487_, _05248_, _07427_);
  nor _66089_ (_14488_, _12718_, _06830_);
  or _66090_ (_14489_, _14488_, _14487_);
  and _66091_ (_14490_, _14489_, _03222_);
  nor _66092_ (_14491_, _05910_, _07427_);
  and _66093_ (_14492_, _12631_, _05910_);
  or _66094_ (_14493_, _14492_, _14491_);
  or _66095_ (_14494_, _14491_, _12648_);
  and _66096_ (_14495_, _14494_, _14493_);
  or _66097_ (_14496_, _14495_, _06840_);
  nor _66098_ (_14497_, _12627_, _06830_);
  or _66099_ (_14498_, _14497_, _14487_);
  or _66100_ (_14499_, _14498_, _04081_);
  and _66101_ (_14500_, _05248_, \oc8051_golden_model_1.ACC [3]);
  or _66102_ (_14501_, _14500_, _14487_);
  and _66103_ (_14502_, _14501_, _04409_);
  nor _66104_ (_14503_, _04409_, _07427_);
  or _66105_ (_14504_, _14503_, _03610_);
  or _66106_ (_14505_, _14504_, _14502_);
  and _66107_ (_14506_, _14505_, _04055_);
  and _66108_ (_14507_, _14506_, _14499_);
  and _66109_ (_14508_, _14493_, _03715_);
  or _66110_ (_14509_, _14508_, _03723_);
  or _66111_ (_14510_, _14509_, _14507_);
  nor _66112_ (_14511_, _06830_, _05005_);
  or _66113_ (_14512_, _14511_, _14487_);
  or _66114_ (_14513_, _14512_, _03996_);
  and _66115_ (_14514_, _14513_, _14510_);
  or _66116_ (_14515_, _14514_, _03729_);
  or _66117_ (_14516_, _14501_, _03737_);
  and _66118_ (_14517_, _14516_, _03736_);
  and _66119_ (_14518_, _14517_, _14515_);
  and _66120_ (_14519_, _12641_, _05910_);
  or _66121_ (_14520_, _14519_, _14491_);
  and _66122_ (_14521_, _14520_, _03714_);
  or _66123_ (_14522_, _14521_, _03719_);
  or _66124_ (_14523_, _14522_, _14518_);
  and _66125_ (_14524_, _14523_, _14496_);
  or _66126_ (_14525_, _14524_, _06869_);
  nor _66127_ (_14526_, _07358_, _07194_);
  nor _66128_ (_14527_, _14526_, _07359_);
  or _66129_ (_14528_, _14527_, _06875_);
  and _66130_ (_14529_, _14528_, _03710_);
  and _66131_ (_14530_, _14529_, _14525_);
  nor _66132_ (_14531_, _12612_, _07391_);
  or _66133_ (_14532_, _14531_, _14491_);
  and _66134_ (_14533_, _14532_, _03505_);
  or _66135_ (_14534_, _14533_, _07390_);
  or _66136_ (_14535_, _14534_, _14530_);
  or _66137_ (_14536_, _14512_, _06838_);
  and _66138_ (_14537_, _14536_, _14535_);
  or _66139_ (_14538_, _14537_, _04481_);
  and _66140_ (_14539_, _06592_, _05248_);
  or _66141_ (_14540_, _14487_, _07400_);
  or _66142_ (_14541_, _14540_, _14539_);
  and _66143_ (_14542_, _14541_, _03589_);
  and _66144_ (_14543_, _14542_, _14538_);
  or _66145_ (_14544_, _14543_, _14490_);
  and _66146_ (_14545_, _14544_, _07411_);
  nand _66147_ (_14546_, _07760_, _07689_);
  nor _66148_ (_14547_, _14433_, _07699_);
  nor _66149_ (_14548_, _14547_, _07692_);
  and _66150_ (_14549_, _14547_, _07692_);
  or _66151_ (_14550_, _14549_, _14548_);
  or _66152_ (_14551_, _14550_, _07760_);
  and _66153_ (_14552_, _14551_, _07405_);
  and _66154_ (_14553_, _14552_, _14546_);
  or _66155_ (_14554_, _14553_, _08828_);
  or _66156_ (_14555_, _14554_, _14545_);
  and _66157_ (_14556_, _12733_, _05248_);
  or _66158_ (_14557_, _14487_, _07766_);
  or _66159_ (_14558_, _14557_, _14556_);
  and _66160_ (_14559_, _05248_, _06276_);
  or _66161_ (_14560_, _14559_, _14487_);
  or _66162_ (_14561_, _14560_, _05886_);
  and _66163_ (_14562_, _14561_, _07778_);
  and _66164_ (_14563_, _14562_, _14558_);
  and _66165_ (_14564_, _14563_, _14555_);
  and _66166_ (_14565_, _12739_, _05248_);
  or _66167_ (_14566_, _14565_, _14487_);
  and _66168_ (_14567_, _14566_, _03780_);
  or _66169_ (_14568_, _14567_, _14564_);
  and _66170_ (_14569_, _14568_, _07777_);
  or _66171_ (_14570_, _14487_, _05567_);
  and _66172_ (_14571_, _14560_, _03622_);
  and _66173_ (_14572_, _14571_, _14570_);
  or _66174_ (_14573_, _14572_, _14569_);
  and _66175_ (_14574_, _14573_, _06828_);
  and _66176_ (_14575_, _14501_, _03790_);
  and _66177_ (_14576_, _14575_, _14570_);
  or _66178_ (_14577_, _14576_, _03624_);
  or _66179_ (_14578_, _14577_, _14574_);
  nor _66180_ (_14579_, _12732_, _06830_);
  or _66181_ (_14580_, _14487_, _07795_);
  or _66182_ (_14581_, _14580_, _14579_);
  and _66183_ (_14582_, _14581_, _07793_);
  and _66184_ (_14583_, _14582_, _14578_);
  nor _66185_ (_14584_, _12738_, _06830_);
  or _66186_ (_14585_, _14584_, _14487_);
  and _66187_ (_14586_, _14585_, _03785_);
  or _66188_ (_14587_, _14586_, _03815_);
  or _66189_ (_14588_, _14587_, _14583_);
  or _66190_ (_14589_, _14498_, _04246_);
  and _66191_ (_14590_, _14589_, _03823_);
  and _66192_ (_14591_, _14590_, _14588_);
  and _66193_ (_14592_, _14520_, _03453_);
  or _66194_ (_14593_, _14592_, _03447_);
  or _66195_ (_14594_, _14593_, _14591_);
  and _66196_ (_14595_, _12794_, _05248_);
  or _66197_ (_14596_, _14487_, _03514_);
  or _66198_ (_14597_, _14596_, _14595_);
  and _66199_ (_14598_, _14597_, _43000_);
  and _66200_ (_14599_, _14598_, _14594_);
  or _66201_ (_14600_, _14599_, _14486_);
  and _66202_ (_43485_, _14600_, _41806_);
  nor _66203_ (_14601_, _43000_, _07550_);
  nor _66204_ (_14602_, _05248_, _07550_);
  nor _66205_ (_14603_, _12933_, _06830_);
  or _66206_ (_14604_, _14603_, _14602_);
  and _66207_ (_14605_, _14604_, _03222_);
  nor _66208_ (_14606_, _05777_, _06830_);
  or _66209_ (_14607_, _14606_, _14602_);
  or _66210_ (_14608_, _14607_, _06838_);
  nor _66211_ (_14609_, _05910_, _07550_);
  and _66212_ (_14610_, _12827_, _05910_);
  or _66213_ (_14611_, _14610_, _14609_);
  and _66214_ (_14612_, _14611_, _03714_);
  nor _66215_ (_14613_, _12841_, _06830_);
  or _66216_ (_14614_, _14613_, _14602_);
  or _66217_ (_14615_, _14614_, _04081_);
  and _66218_ (_14616_, _05248_, \oc8051_golden_model_1.ACC [4]);
  or _66219_ (_14617_, _14616_, _14602_);
  and _66220_ (_14618_, _14617_, _04409_);
  nor _66221_ (_14619_, _04409_, _07550_);
  or _66222_ (_14620_, _14619_, _03610_);
  or _66223_ (_14621_, _14620_, _14618_);
  and _66224_ (_14622_, _14621_, _04055_);
  and _66225_ (_14623_, _14622_, _14615_);
  and _66226_ (_14624_, _12845_, _05910_);
  or _66227_ (_14625_, _14624_, _14609_);
  and _66228_ (_14626_, _14625_, _03715_);
  or _66229_ (_14627_, _14626_, _03723_);
  or _66230_ (_14628_, _14627_, _14623_);
  or _66231_ (_14629_, _14607_, _03996_);
  and _66232_ (_14630_, _14629_, _14628_);
  or _66233_ (_14631_, _14630_, _03729_);
  or _66234_ (_14632_, _14617_, _03737_);
  and _66235_ (_14633_, _14632_, _03736_);
  and _66236_ (_14634_, _14633_, _14631_);
  or _66237_ (_14635_, _14634_, _14612_);
  and _66238_ (_14636_, _14635_, _06840_);
  or _66239_ (_14637_, _14609_, _12860_);
  and _66240_ (_14638_, _14637_, _03719_);
  and _66241_ (_14639_, _14638_, _14625_);
  or _66242_ (_14640_, _14639_, _06869_);
  or _66243_ (_14641_, _14640_, _14636_);
  nor _66244_ (_14642_, _07363_, _07361_);
  nor _66245_ (_14643_, _14642_, _07364_);
  or _66246_ (_14644_, _14643_, _06875_);
  and _66247_ (_14645_, _14644_, _03710_);
  and _66248_ (_14646_, _14645_, _14641_);
  nor _66249_ (_14647_, _12825_, _07391_);
  or _66250_ (_14648_, _14647_, _14609_);
  and _66251_ (_14649_, _14648_, _03505_);
  or _66252_ (_14650_, _14649_, _07390_);
  or _66253_ (_14651_, _14650_, _14646_);
  and _66254_ (_14652_, _14651_, _14608_);
  or _66255_ (_14653_, _14652_, _04481_);
  and _66256_ (_14654_, _06730_, _05248_);
  or _66257_ (_14655_, _14602_, _07400_);
  or _66258_ (_14656_, _14655_, _14654_);
  and _66259_ (_14657_, _14656_, _03589_);
  and _66260_ (_14658_, _14657_, _14653_);
  or _66261_ (_14659_, _14658_, _14605_);
  and _66262_ (_14660_, _14659_, _07411_);
  or _66263_ (_14661_, _14429_, _07727_);
  nor _66264_ (_14662_, _14547_, _07691_);
  or _66265_ (_14663_, _14662_, _07690_);
  nand _66266_ (_14664_, _14663_, _07730_);
  or _66267_ (_14665_, _14663_, _07730_);
  and _66268_ (_14666_, _14665_, _14664_);
  or _66269_ (_14667_, _14666_, _07760_);
  and _66270_ (_14668_, _14667_, _07405_);
  and _66271_ (_14669_, _14668_, _14661_);
  or _66272_ (_14670_, _14669_, _08828_);
  or _66273_ (_14671_, _14670_, _14660_);
  and _66274_ (_14672_, _12821_, _05248_);
  or _66275_ (_14673_, _14602_, _07766_);
  or _66276_ (_14674_, _14673_, _14672_);
  and _66277_ (_14675_, _06298_, _05248_);
  or _66278_ (_14676_, _14675_, _14602_);
  or _66279_ (_14677_, _14676_, _05886_);
  and _66280_ (_14678_, _14677_, _07778_);
  and _66281_ (_14679_, _14678_, _14674_);
  and _66282_ (_14680_, _14679_, _14671_);
  and _66283_ (_14681_, _12817_, _05248_);
  or _66284_ (_14682_, _14681_, _14602_);
  and _66285_ (_14683_, _14682_, _03780_);
  or _66286_ (_14684_, _14683_, _14680_);
  and _66287_ (_14685_, _14684_, _07777_);
  or _66288_ (_14686_, _14602_, _05825_);
  and _66289_ (_14687_, _14676_, _03622_);
  and _66290_ (_14688_, _14687_, _14686_);
  or _66291_ (_14689_, _14688_, _14685_);
  and _66292_ (_14690_, _14689_, _06828_);
  and _66293_ (_14691_, _14617_, _03790_);
  and _66294_ (_14692_, _14691_, _14686_);
  or _66295_ (_14693_, _14692_, _03624_);
  or _66296_ (_14694_, _14693_, _14690_);
  nor _66297_ (_14695_, _12819_, _06830_);
  or _66298_ (_14696_, _14602_, _07795_);
  or _66299_ (_14697_, _14696_, _14695_);
  and _66300_ (_14698_, _14697_, _07793_);
  and _66301_ (_14699_, _14698_, _14694_);
  nor _66302_ (_14700_, _12816_, _06830_);
  or _66303_ (_14701_, _14700_, _14602_);
  and _66304_ (_14702_, _14701_, _03785_);
  or _66305_ (_14703_, _14702_, _03815_);
  or _66306_ (_14704_, _14703_, _14699_);
  or _66307_ (_14705_, _14614_, _04246_);
  and _66308_ (_14706_, _14705_, _03823_);
  and _66309_ (_14707_, _14706_, _14704_);
  and _66310_ (_14708_, _14611_, _03453_);
  or _66311_ (_14709_, _14708_, _03447_);
  or _66312_ (_14710_, _14709_, _14707_);
  and _66313_ (_14711_, _13003_, _05248_);
  or _66314_ (_14712_, _14602_, _03514_);
  or _66315_ (_14713_, _14712_, _14711_);
  and _66316_ (_14714_, _14713_, _43000_);
  and _66317_ (_14715_, _14714_, _14710_);
  or _66318_ (_14716_, _14715_, _14601_);
  and _66319_ (_43486_, _14716_, _41806_);
  nor _66320_ (_14717_, _43000_, _07541_);
  nor _66321_ (_14718_, _05248_, _07541_);
  nor _66322_ (_14719_, _13127_, _06830_);
  or _66323_ (_14720_, _14719_, _14718_);
  and _66324_ (_14721_, _14720_, _03222_);
  nor _66325_ (_14722_, _05469_, _06830_);
  or _66326_ (_14723_, _14722_, _14718_);
  or _66327_ (_14724_, _14723_, _06838_);
  nor _66328_ (_14725_, _05910_, _07541_);
  and _66329_ (_14726_, _13047_, _05910_);
  or _66330_ (_14727_, _14726_, _14725_);
  and _66331_ (_14728_, _14727_, _03714_);
  nor _66332_ (_14729_, _13014_, _06830_);
  or _66333_ (_14730_, _14729_, _14718_);
  and _66334_ (_14731_, _14730_, _03610_);
  nor _66335_ (_14732_, _04409_, _07541_);
  and _66336_ (_14733_, _05248_, \oc8051_golden_model_1.ACC [5]);
  or _66337_ (_14734_, _14733_, _14718_);
  and _66338_ (_14735_, _14734_, _04409_);
  or _66339_ (_14736_, _14735_, _14732_);
  and _66340_ (_14737_, _14736_, _04081_);
  or _66341_ (_14738_, _14737_, _14265_);
  or _66342_ (_14739_, _14738_, _14731_);
  and _66343_ (_14740_, _13037_, _05910_);
  or _66344_ (_14741_, _14740_, _14725_);
  or _66345_ (_14742_, _14741_, _04055_);
  or _66346_ (_14743_, _14723_, _03996_);
  and _66347_ (_14744_, _14743_, _14742_);
  and _66348_ (_14745_, _14744_, _14739_);
  or _66349_ (_14746_, _14745_, _03729_);
  or _66350_ (_14747_, _14734_, _03737_);
  and _66351_ (_14748_, _14747_, _03736_);
  and _66352_ (_14749_, _14748_, _14746_);
  or _66353_ (_14750_, _14749_, _14728_);
  and _66354_ (_14751_, _14750_, _06840_);
  or _66355_ (_14752_, _14725_, _13054_);
  and _66356_ (_14753_, _14752_, _03719_);
  and _66357_ (_14754_, _14753_, _14741_);
  or _66358_ (_14755_, _14754_, _06869_);
  or _66359_ (_14756_, _14755_, _14751_);
  nor _66360_ (_14757_, _07366_, _07068_);
  nor _66361_ (_14758_, _14757_, _07367_);
  or _66362_ (_14759_, _14758_, _06875_);
  and _66363_ (_14760_, _14759_, _03710_);
  and _66364_ (_14761_, _14760_, _14756_);
  nor _66365_ (_14762_, _13020_, _07391_);
  or _66366_ (_14763_, _14762_, _14725_);
  and _66367_ (_14764_, _14763_, _03505_);
  or _66368_ (_14765_, _14764_, _07390_);
  or _66369_ (_14766_, _14765_, _14761_);
  and _66370_ (_14767_, _14766_, _14724_);
  or _66371_ (_14768_, _14767_, _04481_);
  and _66372_ (_14769_, _06684_, _05248_);
  or _66373_ (_14770_, _14718_, _07400_);
  or _66374_ (_14771_, _14770_, _14769_);
  and _66375_ (_14772_, _14771_, _03589_);
  and _66376_ (_14773_, _14772_, _14768_);
  or _66377_ (_14774_, _14773_, _14721_);
  and _66378_ (_14775_, _14774_, _07411_);
  nand _66379_ (_14776_, _07760_, _07737_);
  not _66380_ (_14777_, _07729_);
  and _66381_ (_14778_, _14664_, _14777_);
  and _66382_ (_14779_, _14778_, _07740_);
  nor _66383_ (_14780_, _14778_, _07740_);
  or _66384_ (_14781_, _14780_, _14779_);
  or _66385_ (_14782_, _14781_, _07760_);
  and _66386_ (_14783_, _14782_, _07405_);
  and _66387_ (_14784_, _14783_, _14776_);
  or _66388_ (_14785_, _14784_, _08828_);
  or _66389_ (_14786_, _14785_, _14775_);
  and _66390_ (_14787_, _13141_, _05248_);
  or _66391_ (_14788_, _14718_, _07766_);
  or _66392_ (_14789_, _14788_, _14787_);
  and _66393_ (_14790_, _06306_, _05248_);
  or _66394_ (_14791_, _14790_, _14718_);
  or _66395_ (_14792_, _14791_, _05886_);
  and _66396_ (_14793_, _14792_, _07778_);
  and _66397_ (_14794_, _14793_, _14789_);
  and _66398_ (_14795_, _14794_, _14786_);
  and _66399_ (_14796_, _13147_, _05248_);
  or _66400_ (_14797_, _14796_, _14718_);
  and _66401_ (_14798_, _14797_, _03780_);
  or _66402_ (_14799_, _14798_, _14795_);
  and _66403_ (_14800_, _14799_, _07777_);
  or _66404_ (_14801_, _14718_, _05518_);
  and _66405_ (_14802_, _14791_, _03622_);
  and _66406_ (_14803_, _14802_, _14801_);
  or _66407_ (_14804_, _14803_, _14800_);
  and _66408_ (_14805_, _14804_, _06828_);
  and _66409_ (_14806_, _14734_, _03790_);
  and _66410_ (_14807_, _14806_, _14801_);
  or _66411_ (_14808_, _14807_, _03624_);
  or _66412_ (_14809_, _14808_, _14805_);
  nor _66413_ (_14810_, _13140_, _06830_);
  or _66414_ (_14811_, _14718_, _07795_);
  or _66415_ (_14812_, _14811_, _14810_);
  and _66416_ (_14813_, _14812_, _07793_);
  and _66417_ (_14814_, _14813_, _14809_);
  nor _66418_ (_14815_, _13146_, _06830_);
  or _66419_ (_14816_, _14815_, _14718_);
  and _66420_ (_14817_, _14816_, _03785_);
  or _66421_ (_14818_, _14817_, _03815_);
  or _66422_ (_14819_, _14818_, _14814_);
  or _66423_ (_14820_, _14730_, _04246_);
  and _66424_ (_14821_, _14820_, _03823_);
  and _66425_ (_14822_, _14821_, _14819_);
  and _66426_ (_14823_, _14727_, _03453_);
  or _66427_ (_14824_, _14823_, _03447_);
  or _66428_ (_14825_, _14824_, _14822_);
  and _66429_ (_14826_, _13199_, _05248_);
  or _66430_ (_14827_, _14718_, _03514_);
  or _66431_ (_14828_, _14827_, _14826_);
  and _66432_ (_14829_, _14828_, _43000_);
  and _66433_ (_14830_, _14829_, _14825_);
  or _66434_ (_14831_, _14830_, _14717_);
  and _66435_ (_43487_, _14831_, _41806_);
  nor _66436_ (_14832_, _43000_, _07673_);
  nor _66437_ (_14833_, _05248_, _07673_);
  nor _66438_ (_14834_, _13332_, _06830_);
  or _66439_ (_14835_, _14834_, _14833_);
  and _66440_ (_14836_, _14835_, _03222_);
  nor _66441_ (_14837_, _05363_, _06830_);
  or _66442_ (_14838_, _14837_, _14833_);
  or _66443_ (_14839_, _14838_, _06838_);
  nor _66444_ (_14840_, _05910_, _07673_);
  and _66445_ (_14841_, _13253_, _05910_);
  or _66446_ (_14842_, _14841_, _14840_);
  and _66447_ (_14843_, _14842_, _03714_);
  nor _66448_ (_14844_, _13242_, _06830_);
  or _66449_ (_14845_, _14844_, _14833_);
  or _66450_ (_14846_, _14845_, _04081_);
  and _66451_ (_14847_, _05248_, \oc8051_golden_model_1.ACC [6]);
  or _66452_ (_14848_, _14847_, _14833_);
  and _66453_ (_14849_, _14848_, _04409_);
  nor _66454_ (_14850_, _04409_, _07673_);
  or _66455_ (_14851_, _14850_, _03610_);
  or _66456_ (_14852_, _14851_, _14849_);
  and _66457_ (_14853_, _14852_, _04055_);
  and _66458_ (_14854_, _14853_, _14846_);
  and _66459_ (_14855_, _13229_, _05910_);
  or _66460_ (_14856_, _14855_, _14840_);
  and _66461_ (_14857_, _14856_, _03715_);
  or _66462_ (_14858_, _14857_, _03723_);
  or _66463_ (_14859_, _14858_, _14854_);
  or _66464_ (_14860_, _14838_, _03996_);
  and _66465_ (_14861_, _14860_, _14859_);
  or _66466_ (_14862_, _14861_, _03729_);
  or _66467_ (_14863_, _14848_, _03737_);
  and _66468_ (_14864_, _14863_, _03736_);
  and _66469_ (_14865_, _14864_, _14862_);
  or _66470_ (_14866_, _14865_, _14843_);
  and _66471_ (_14867_, _14866_, _06840_);
  or _66472_ (_14868_, _14840_, _13260_);
  and _66473_ (_14869_, _14868_, _03719_);
  and _66474_ (_14870_, _14869_, _14856_);
  or _66475_ (_14871_, _14870_, _06869_);
  or _66476_ (_14872_, _14871_, _14867_);
  nor _66477_ (_14873_, _07382_, _07369_);
  nor _66478_ (_14874_, _14873_, _07383_);
  or _66479_ (_14875_, _14874_, _06875_);
  and _66480_ (_14876_, _14875_, _03710_);
  and _66481_ (_14877_, _14876_, _14872_);
  nor _66482_ (_14878_, _13226_, _07391_);
  or _66483_ (_14879_, _14878_, _14840_);
  and _66484_ (_14880_, _14879_, _03505_);
  or _66485_ (_14881_, _14880_, _07390_);
  or _66486_ (_14882_, _14881_, _14877_);
  and _66487_ (_14883_, _14882_, _14839_);
  or _66488_ (_14884_, _14883_, _04481_);
  and _66489_ (_14885_, _06455_, _05248_);
  or _66490_ (_14886_, _14833_, _07400_);
  or _66491_ (_14887_, _14886_, _14885_);
  and _66492_ (_14888_, _14887_, _03589_);
  and _66493_ (_14889_, _14888_, _14884_);
  or _66494_ (_14890_, _14889_, _14836_);
  and _66495_ (_14891_, _14890_, _07411_);
  nor _66496_ (_14892_, _14778_, _07738_);
  or _66497_ (_14893_, _14892_, _07739_);
  and _66498_ (_14894_, _14893_, _07721_);
  nor _66499_ (_14895_, _14893_, _07721_);
  or _66500_ (_14896_, _14895_, _14894_);
  or _66501_ (_14897_, _14896_, _07760_);
  or _66502_ (_14898_, _14429_, _07679_);
  and _66503_ (_14899_, _14898_, _07405_);
  and _66504_ (_14900_, _14899_, _14897_);
  or _66505_ (_14901_, _14900_, _08828_);
  or _66506_ (_14902_, _14901_, _14891_);
  and _66507_ (_14903_, _13347_, _05248_);
  or _66508_ (_14904_, _14833_, _07766_);
  or _66509_ (_14905_, _14904_, _14903_);
  and _66510_ (_14906_, _13339_, _05248_);
  or _66511_ (_14907_, _14906_, _14833_);
  or _66512_ (_14908_, _14907_, _05886_);
  and _66513_ (_14909_, _14908_, _07778_);
  and _66514_ (_14910_, _14909_, _14905_);
  and _66515_ (_14911_, _14910_, _14902_);
  and _66516_ (_14912_, _13353_, _05248_);
  or _66517_ (_14913_, _14912_, _14833_);
  and _66518_ (_14914_, _14913_, _03780_);
  or _66519_ (_14915_, _14914_, _14911_);
  and _66520_ (_14916_, _14915_, _07777_);
  or _66521_ (_14917_, _14833_, _05412_);
  and _66522_ (_14918_, _14907_, _03622_);
  and _66523_ (_14919_, _14918_, _14917_);
  or _66524_ (_14920_, _14919_, _14916_);
  and _66525_ (_14921_, _14920_, _06828_);
  and _66526_ (_14922_, _14848_, _03790_);
  and _66527_ (_14923_, _14922_, _14917_);
  or _66528_ (_14924_, _14923_, _03624_);
  or _66529_ (_14925_, _14924_, _14921_);
  nor _66530_ (_14926_, _13346_, _06830_);
  or _66531_ (_14927_, _14833_, _07795_);
  or _66532_ (_14928_, _14927_, _14926_);
  and _66533_ (_14929_, _14928_, _07793_);
  and _66534_ (_14930_, _14929_, _14925_);
  nor _66535_ (_14931_, _13352_, _06830_);
  or _66536_ (_14932_, _14931_, _14833_);
  and _66537_ (_14933_, _14932_, _03785_);
  or _66538_ (_14934_, _14933_, _03815_);
  or _66539_ (_14935_, _14934_, _14930_);
  or _66540_ (_14936_, _14845_, _04246_);
  and _66541_ (_14937_, _14936_, _03823_);
  and _66542_ (_14938_, _14937_, _14935_);
  and _66543_ (_14939_, _14842_, _03453_);
  or _66544_ (_14940_, _14939_, _03447_);
  or _66545_ (_14941_, _14940_, _14938_);
  and _66546_ (_14942_, _13402_, _05248_);
  or _66547_ (_14943_, _14833_, _03514_);
  or _66548_ (_14944_, _14943_, _14942_);
  and _66549_ (_14945_, _14944_, _43000_);
  and _66550_ (_14946_, _14945_, _14941_);
  or _66551_ (_14947_, _14946_, _14832_);
  and _66552_ (_43488_, _14947_, _41806_);
  nor _66553_ (_14948_, _43000_, _03335_);
  and _66554_ (_14949_, _08780_, \oc8051_golden_model_1.ACC [1]);
  nand _66555_ (_14950_, _08732_, _06075_);
  nand _66556_ (_14951_, _08318_, _03517_);
  and _66557_ (_14952_, _14951_, _08734_);
  and _66558_ (_14953_, _03605_, _03202_);
  and _66559_ (_14954_, _03616_, _03202_);
  nand _66560_ (_14955_, _08458_, _10057_);
  nor _66561_ (_14956_, _05666_, _07908_);
  nor _66562_ (_14957_, _05254_, _03335_);
  and _66563_ (_14958_, _05254_, _06274_);
  nor _66564_ (_14959_, _14958_, _14957_);
  nor _66565_ (_14960_, _14959_, _14956_);
  and _66566_ (_14961_, _14960_, _03622_);
  nor _66567_ (_14962_, _04198_, _04197_);
  or _66568_ (_14963_, _14962_, _08681_);
  and _66569_ (_14964_, _12124_, _05254_);
  nor _66570_ (_14965_, _14964_, _14957_);
  nand _66571_ (_14966_, _14965_, _03600_);
  or _66572_ (_14967_, _12128_, _03779_);
  and _66573_ (_14968_, _14967_, _07905_);
  nand _66574_ (_14969_, _04048_, _03216_);
  and _66575_ (_14970_, _05254_, _04620_);
  nor _66576_ (_14971_, _14970_, _14957_);
  nand _66577_ (_14972_, _14971_, _07390_);
  nand _66578_ (_14973_, _07974_, _07913_);
  or _66579_ (_14974_, _08063_, _04620_);
  nor _66580_ (_14975_, _08066_, _04422_);
  or _66581_ (_14976_, _14975_, _06546_);
  and _66582_ (_14977_, _08079_, _04620_);
  or _66583_ (_14978_, _04064_, \oc8051_golden_model_1.ACC [0]);
  nand _66584_ (_14979_, _04064_, \oc8051_golden_model_1.ACC [0]);
  and _66585_ (_14980_, _14979_, _14978_);
  and _66586_ (_14981_, _14980_, _08078_);
  or _66587_ (_14982_, _14981_, _08066_);
  or _66588_ (_14983_, _14982_, _14977_);
  and _66589_ (_14984_, _14983_, _03235_);
  or _66590_ (_14985_, _14984_, _04422_);
  and _66591_ (_14986_, _14985_, _04081_);
  and _66592_ (_14987_, _14986_, _14976_);
  nor _66593_ (_14988_, _14957_, _14956_);
  nor _66594_ (_14989_, _14988_, _04081_);
  or _66595_ (_14990_, _14989_, _03715_);
  or _66596_ (_14991_, _14990_, _14987_);
  nor _66597_ (_14992_, _05903_, _03335_);
  and _66598_ (_14993_, _12021_, _05903_);
  nor _66599_ (_14994_, _14993_, _14992_);
  nand _66600_ (_14995_, _14994_, _03715_);
  and _66601_ (_14996_, _14995_, _03996_);
  and _66602_ (_14997_, _14996_, _14991_);
  nor _66603_ (_14998_, _14971_, _03996_);
  or _66604_ (_14999_, _14998_, _08064_);
  or _66605_ (_15000_, _14999_, _14997_);
  and _66606_ (_15001_, _15000_, _14974_);
  or _66607_ (_15002_, _15001_, _04443_);
  or _66608_ (_15003_, _06546_, _08128_);
  and _66609_ (_15004_, _15003_, _03737_);
  and _66610_ (_15005_, _15004_, _15002_);
  nor _66611_ (_15006_, _08285_, _03737_);
  or _66612_ (_15007_, _15006_, _08132_);
  or _66613_ (_15008_, _15007_, _15005_);
  nand _66614_ (_15009_, _08132_, _07484_);
  and _66615_ (_15010_, _15009_, _15008_);
  or _66616_ (_15011_, _15010_, _03714_);
  or _66617_ (_15012_, _14957_, _03736_);
  and _66618_ (_15013_, _15012_, _06840_);
  and _66619_ (_15014_, _15013_, _15011_);
  nor _66620_ (_15015_, _14988_, _06840_);
  or _66621_ (_15016_, _15015_, _06869_);
  or _66622_ (_15017_, _15016_, _15014_);
  nand _66623_ (_15018_, _03494_, _03223_);
  or _66624_ (_15019_, _15018_, _12559_);
  not _66625_ (_15020_, _07330_);
  nand _66626_ (_15021_, _15020_, _06869_);
  and _66627_ (_15022_, _15021_, _15019_);
  and _66628_ (_15023_, _15022_, _08058_);
  and _66629_ (_15024_, _15023_, _15017_);
  nor _66630_ (_15025_, _08170_, _08059_);
  or _66631_ (_15026_, _15025_, _08051_);
  or _66632_ (_15027_, _15026_, _15024_);
  nor _66633_ (_15028_, _08035_, _03335_);
  nor _66634_ (_15029_, _15028_, _08036_);
  nand _66635_ (_15030_, _08051_, _15029_);
  and _66636_ (_15031_, _15030_, _03766_);
  and _66637_ (_15032_, _15031_, _15027_);
  nor _66638_ (_15033_, _08566_, _03335_);
  nor _66639_ (_15034_, _15033_, _10217_);
  nand _66640_ (_15035_, _15034_, _07914_);
  and _66641_ (_15036_, _15035_, _08187_);
  or _66642_ (_15037_, _15036_, _15032_);
  and _66643_ (_15038_, _15037_, _14973_);
  or _66644_ (_15039_, _15038_, _07912_);
  nand _66645_ (_15040_, _04048_, _07912_);
  and _66646_ (_15041_, _15040_, _03710_);
  and _66647_ (_15042_, _15041_, _15039_);
  nor _66648_ (_15043_, _12052_, _08339_);
  nor _66649_ (_15044_, _15043_, _14992_);
  nor _66650_ (_15045_, _15044_, _03710_);
  or _66651_ (_15046_, _15045_, _07390_);
  or _66652_ (_15047_, _15046_, _15042_);
  and _66653_ (_15048_, _15047_, _14972_);
  or _66654_ (_15049_, _15048_, _04481_);
  and _66655_ (_15050_, _06546_, _05254_);
  nor _66656_ (_15051_, _15050_, _14957_);
  nand _66657_ (_15052_, _15051_, _04481_);
  and _66658_ (_15053_, _15052_, _03589_);
  and _66659_ (_15054_, _15053_, _15049_);
  nor _66660_ (_15055_, _12109_, _07908_);
  nor _66661_ (_15056_, _15055_, _14957_);
  nor _66662_ (_15057_, _15056_, _03589_);
  or _66663_ (_15058_, _15057_, _07405_);
  or _66664_ (_15059_, _15058_, _15054_);
  nand _66665_ (_15060_, _07760_, _07405_);
  and _66666_ (_15061_, _15060_, _15059_);
  or _66667_ (_15062_, _15061_, _03216_);
  and _66668_ (_15063_, _15062_, _14969_);
  or _66669_ (_15064_, _15063_, _03601_);
  nand _66670_ (_15065_, _14959_, _03601_);
  and _66671_ (_15066_, _15065_, _08364_);
  and _66672_ (_15067_, _15066_, _15064_);
  nor _66673_ (_15068_, _08364_, _04048_);
  or _66674_ (_15069_, _15068_, _08371_);
  or _66675_ (_15070_, _15069_, _15067_);
  and _66676_ (_15071_, _04634_, _03335_);
  nor _66677_ (_15072_, _15071_, _08681_);
  or _66678_ (_15073_, _08377_, _15072_);
  and _66679_ (_15074_, _15073_, _08383_);
  and _66680_ (_15075_, _15074_, _15070_);
  or _66681_ (_15076_, _08386_, _15072_);
  and _66682_ (_15077_, _15076_, _08388_);
  or _66683_ (_15078_, _15077_, _15075_);
  or _66684_ (_15079_, _08394_, _15072_);
  and _66685_ (_15080_, _15079_, _08393_);
  and _66686_ (_15081_, _15080_, _15078_);
  nor _66687_ (_15082_, _06546_, \oc8051_golden_model_1.ACC [0]);
  nor _66688_ (_15083_, _15082_, _08645_);
  and _66689_ (_15084_, _08392_, _15083_);
  or _66690_ (_15085_, _15084_, _03778_);
  or _66691_ (_15086_, _15085_, _15081_);
  and _66692_ (_15087_, _15086_, _14968_);
  and _66693_ (_15088_, _10058_, _07904_);
  or _66694_ (_15089_, _15088_, _03600_);
  or _66695_ (_15090_, _15089_, _15087_);
  and _66696_ (_15091_, _15090_, _14966_);
  or _66697_ (_15092_, _15091_, _03780_);
  not _66698_ (_15093_, _03592_);
  and _66699_ (_15094_, _08070_, _15093_);
  nor _66700_ (_15095_, _15094_, _04193_);
  nor _66701_ (_15096_, _15095_, _03982_);
  or _66702_ (_15097_, _14957_, _07778_);
  and _66703_ (_15098_, _15097_, _15096_);
  and _66704_ (_15099_, _15098_, _15092_);
  nor _66705_ (_15100_, _10321_, _04193_);
  not _66706_ (_15101_, _15100_);
  and _66707_ (_15102_, _15096_, _15101_);
  not _66708_ (_15103_, _15102_);
  or _66709_ (_15104_, _15100_, _08681_);
  and _66710_ (_15105_, _15104_, _15103_);
  or _66711_ (_15106_, _15105_, _04199_);
  or _66712_ (_15107_, _15106_, _15099_);
  and _66713_ (_15108_, _15107_, _14963_);
  or _66714_ (_15109_, _15108_, _08420_);
  or _66715_ (_15110_, _08425_, _08645_);
  and _66716_ (_15111_, _15110_, _03789_);
  and _66717_ (_15112_, _15111_, _15109_);
  or _66718_ (_15113_, _12005_, _08429_);
  and _66719_ (_15114_, _15113_, _08431_);
  or _66720_ (_15115_, _15114_, _15112_);
  or _66721_ (_15116_, _08435_, _08751_);
  and _66722_ (_15117_, _15116_, _07777_);
  and _66723_ (_15118_, _15117_, _15115_);
  or _66724_ (_15119_, _15118_, _14961_);
  nor _66725_ (_15120_, _07895_, _04190_);
  not _66726_ (_15121_, _15120_);
  and _66727_ (_15122_, _15121_, _15119_);
  nor _66728_ (_15123_, _10321_, _04190_);
  nor _66729_ (_15124_, _15121_, _15071_);
  or _66730_ (_15125_, _15124_, _15123_);
  or _66731_ (_15126_, _15125_, _15122_);
  and _66732_ (_15127_, _04058_, _03200_);
  not _66733_ (_15128_, _15127_);
  nand _66734_ (_15129_, _15123_, _15071_);
  and _66735_ (_15130_, _15129_, _15128_);
  and _66736_ (_15131_, _15130_, _15126_);
  nor _66737_ (_15132_, _15071_, _15128_);
  or _66738_ (_15133_, _15132_, _08450_);
  or _66739_ (_15134_, _15133_, _15131_);
  nand _66740_ (_15135_, _08450_, _15082_);
  and _66741_ (_15136_, _15135_, _03784_);
  and _66742_ (_15137_, _15136_, _15134_);
  nand _66743_ (_15138_, _12003_, _08461_);
  and _66744_ (_15139_, _15138_, _08460_);
  or _66745_ (_15140_, _15139_, _15137_);
  and _66746_ (_15141_, _15140_, _14955_);
  or _66747_ (_15142_, _15141_, _03624_);
  nor _66748_ (_15143_, _12122_, _07908_);
  nor _66749_ (_15144_, _15143_, _14957_);
  nand _66750_ (_15145_, _15144_, _03624_);
  and _66751_ (_15146_, _15145_, _07898_);
  and _66752_ (_15147_, _15146_, _15142_);
  nor _66753_ (_15148_, _08170_, _07898_);
  or _66754_ (_15149_, _15148_, _08475_);
  or _66755_ (_15150_, _15149_, _15147_);
  nand _66756_ (_15151_, _08475_, _15029_);
  and _66757_ (_15152_, _15151_, _15150_);
  or _66758_ (_15153_, _15152_, _03776_);
  nand _66759_ (_15154_, _15034_, _03776_);
  and _66760_ (_15155_, _15154_, _08589_);
  and _66761_ (_15156_, _15155_, _15153_);
  nor _66762_ (_15157_, _08589_, _07974_);
  or _66763_ (_15158_, _15157_, _08587_);
  or _66764_ (_15159_, _15158_, _15156_);
  nand _66765_ (_15160_, _08587_, _07871_);
  and _66766_ (_15161_, _15160_, _08617_);
  and _66767_ (_15162_, _15161_, _15159_);
  and _66768_ (_15163_, _08618_, _15072_);
  nor _66769_ (_15164_, _15163_, _15162_);
  or _66770_ (_15165_, _15164_, _14954_);
  nand _66771_ (_15166_, _14954_, _15083_);
  and _66772_ (_15167_, _15166_, _15165_);
  nor _66773_ (_15168_, _15167_, _14953_);
  and _66774_ (_15169_, _15083_, _14953_);
  or _66775_ (_15170_, _15169_, _03517_);
  or _66776_ (_15171_, _15170_, _15168_);
  and _66777_ (_15172_, _15171_, _14952_);
  and _66778_ (_15173_, _08701_, _10058_);
  or _66779_ (_15174_, _15173_, _08732_);
  or _66780_ (_15175_, _15174_, _15172_);
  and _66781_ (_15176_, _15175_, _14950_);
  or _66782_ (_15177_, _15176_, _03815_);
  nand _66783_ (_15178_, _14988_, _03815_);
  and _66784_ (_15179_, _15178_, _08776_);
  and _66785_ (_15180_, _15179_, _15177_);
  and _66786_ (_15181_, _08775_, _03335_);
  or _66787_ (_15182_, _15181_, _15180_);
  and _66788_ (_15183_, _15182_, _10359_);
  or _66789_ (_15184_, _15183_, _14949_);
  and _66790_ (_15185_, _15184_, _03823_);
  and _66791_ (_15186_, _14957_, _03453_);
  or _66792_ (_15187_, _15186_, _03447_);
  or _66793_ (_15188_, _15187_, _15185_);
  nand _66794_ (_15189_, _14988_, _03447_);
  and _66795_ (_15190_, _15189_, _08799_);
  and _66796_ (_15191_, _15190_, _15188_);
  and _66797_ (_15192_, _08798_, _03335_);
  or _66798_ (_15193_, _15192_, _08805_);
  or _66799_ (_15194_, _15193_, _15191_);
  nand _66800_ (_15195_, _08805_, _03274_);
  and _66801_ (_15196_, _15195_, _43000_);
  and _66802_ (_15197_, _15196_, _15194_);
  or _66803_ (_15198_, _15197_, _14948_);
  and _66804_ (_43491_, _15198_, _41806_);
  nor _66805_ (_15199_, _43000_, _03274_);
  nand _66806_ (_15200_, _08732_, _03335_);
  nor _66807_ (_15201_, _08645_, _08644_);
  nor _66808_ (_15202_, _15201_, _08646_);
  or _66809_ (_15203_, _15202_, _08624_);
  nor _66810_ (_15204_, _05254_, _03274_);
  and _66811_ (_15205_, _12207_, _05254_);
  nor _66812_ (_15206_, _15205_, _15204_);
  nor _66813_ (_15207_, _15206_, _07777_);
  and _66814_ (_15208_, _12327_, _05254_);
  nor _66815_ (_15209_, _15208_, _15204_);
  and _66816_ (_15210_, _15209_, _03600_);
  nand _66817_ (_15211_, _03414_, _03216_);
  and _66818_ (_15212_, _05254_, _06764_);
  nor _66819_ (_15213_, _15212_, _15204_);
  nand _66820_ (_15214_, _15213_, _07390_);
  or _66821_ (_15215_, _08063_, _06764_);
  or _66822_ (_15216_, _08078_, _06764_);
  nor _66823_ (_15217_, _04064_, _03274_);
  and _66824_ (_15218_, _04064_, _03274_);
  nor _66825_ (_15219_, _15218_, _15217_);
  nand _66826_ (_15220_, _15219_, _08078_);
  and _66827_ (_15221_, _15220_, _08067_);
  and _66828_ (_15222_, _15221_, _15216_);
  or _66829_ (_15223_, _15222_, _08066_);
  and _66830_ (_15224_, _15223_, _03235_);
  or _66831_ (_15225_, _15224_, _04422_);
  and _66832_ (_15226_, _15222_, _05966_);
  or _66833_ (_15227_, _15226_, _06501_);
  and _66834_ (_15228_, _15227_, _15225_);
  or _66835_ (_15229_, _15228_, _03610_);
  nor _66836_ (_15230_, _05254_, \oc8051_golden_model_1.ACC [1]);
  and _66837_ (_15231_, _12213_, _05254_);
  nor _66838_ (_15232_, _15231_, _15230_);
  or _66839_ (_15233_, _15232_, _04081_);
  and _66840_ (_15234_, _15233_, _15229_);
  or _66841_ (_15235_, _15234_, _08089_);
  nor _66842_ (_15236_, _08096_, \oc8051_golden_model_1.PSW [6]);
  nor _66843_ (_15237_, _15236_, \oc8051_golden_model_1.ACC [1]);
  and _66844_ (_15238_, _15236_, \oc8051_golden_model_1.ACC [1]);
  nor _66845_ (_15239_, _15238_, _15237_);
  nand _66846_ (_15240_, _15239_, _08089_);
  and _66847_ (_15241_, _15240_, _03730_);
  and _66848_ (_15242_, _15241_, _15235_);
  nor _66849_ (_15243_, _05903_, _03274_);
  and _66850_ (_15244_, _12224_, _05903_);
  nor _66851_ (_15245_, _15244_, _15243_);
  nor _66852_ (_15246_, _15245_, _04055_);
  nor _66853_ (_15247_, _15213_, _03996_);
  or _66854_ (_15248_, _15247_, _08064_);
  or _66855_ (_15249_, _15248_, _15246_);
  or _66856_ (_15250_, _15249_, _15242_);
  and _66857_ (_15251_, _15250_, _15215_);
  or _66858_ (_15252_, _15251_, _04443_);
  or _66859_ (_15253_, _06501_, _08128_);
  and _66860_ (_15254_, _15253_, _03737_);
  and _66861_ (_15255_, _15254_, _15252_);
  nor _66862_ (_15256_, _08271_, _03737_);
  or _66863_ (_15257_, _15256_, _08132_);
  or _66864_ (_15258_, _15257_, _15255_);
  nand _66865_ (_15259_, _08132_, _07478_);
  and _66866_ (_15260_, _15259_, _15258_);
  or _66867_ (_15261_, _15260_, _03714_);
  and _66868_ (_15262_, _12211_, _05903_);
  nor _66869_ (_15263_, _15262_, _15243_);
  nand _66870_ (_15264_, _15263_, _03714_);
  and _66871_ (_15265_, _15264_, _06840_);
  and _66872_ (_15266_, _15265_, _15261_);
  and _66873_ (_15267_, _15244_, _12239_);
  nor _66874_ (_15268_, _15267_, _15243_);
  nor _66875_ (_15269_, _15268_, _06840_);
  or _66876_ (_15270_, _15269_, _06869_);
  or _66877_ (_15271_, _15270_, _15266_);
  and _66878_ (_15272_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor _66879_ (_15273_, _15272_, _07703_);
  nor _66880_ (_15274_, _15273_, _07331_);
  or _66881_ (_15275_, _15274_, _06875_);
  and _66882_ (_15276_, _15275_, _08059_);
  and _66883_ (_15277_, _15276_, _15271_);
  and _66884_ (_15278_, \oc8051_golden_model_1.PSW [7], _03335_);
  and _66885_ (_15279_, _07871_, \oc8051_golden_model_1.ACC [0]);
  not _66886_ (_15280_, _15279_);
  and _66887_ (_15281_, _15280_, _04620_);
  nor _66888_ (_15282_, _15281_, _15278_);
  and _66889_ (_15283_, _15282_, _08680_);
  nor _66890_ (_15284_, _15282_, _08680_);
  or _66891_ (_15285_, _15284_, _15283_);
  nor _66892_ (_15286_, _15285_, _08051_);
  nor _66893_ (_15287_, _15286_, _11350_);
  or _66894_ (_15288_, _15287_, _15277_);
  and _66895_ (_15289_, _15280_, _06546_);
  nor _66896_ (_15290_, _15289_, _15278_);
  and _66897_ (_15291_, _15290_, _08644_);
  nor _66898_ (_15292_, _15290_, _08644_);
  or _66899_ (_15293_, _15292_, _15291_);
  or _66900_ (_15294_, _10201_, _15293_);
  and _66901_ (_15295_, _15294_, _15288_);
  or _66902_ (_15296_, _15295_, _03761_);
  nor _66903_ (_15297_, _08285_, _15279_);
  nor _66904_ (_15298_, _15297_, _15278_);
  and _66905_ (_15299_, _15298_, _08316_);
  nor _66906_ (_15300_, _15298_, _08316_);
  or _66907_ (_15301_, _15300_, _15299_);
  nand _66908_ (_15302_, _15301_, _03761_);
  and _66909_ (_15303_, _15302_, _07914_);
  and _66910_ (_15304_, _15303_, _15296_);
  nor _66911_ (_15305_, _15279_, _04048_);
  nor _66912_ (_15306_, _15305_, _15278_);
  and _66913_ (_15307_, _15306_, _08753_);
  nor _66914_ (_15308_, _15306_, _08753_);
  or _66915_ (_15309_, _15308_, _15307_);
  and _66916_ (_15310_, _15309_, _07913_);
  or _66917_ (_15311_, _15310_, _07912_);
  or _66918_ (_15312_, _15311_, _15304_);
  nand _66919_ (_15313_, _03414_, _07912_);
  and _66920_ (_15314_, _15313_, _03710_);
  and _66921_ (_15315_, _15314_, _15312_);
  nor _66922_ (_15316_, _12256_, _08339_);
  nor _66923_ (_15317_, _15316_, _15243_);
  nor _66924_ (_15318_, _15317_, _03710_);
  or _66925_ (_15319_, _15318_, _07390_);
  or _66926_ (_15320_, _15319_, _15315_);
  and _66927_ (_15321_, _15320_, _15214_);
  or _66928_ (_15322_, _15321_, _04481_);
  and _66929_ (_15323_, _06501_, _05254_);
  nor _66930_ (_15324_, _15323_, _15204_);
  nand _66931_ (_15325_, _15324_, _04481_);
  and _66932_ (_15326_, _15325_, _03589_);
  and _66933_ (_15327_, _15326_, _15322_);
  nor _66934_ (_15328_, _12313_, _07908_);
  nor _66935_ (_15329_, _15328_, _15204_);
  nor _66936_ (_15330_, _15329_, _03589_);
  or _66937_ (_15331_, _15330_, _07405_);
  or _66938_ (_15332_, _15331_, _15327_);
  or _66939_ (_15333_, _07668_, _07411_);
  and _66940_ (_15334_, _15333_, _15332_);
  or _66941_ (_15335_, _15334_, _03216_);
  and _66942_ (_15336_, _15335_, _15211_);
  or _66943_ (_15337_, _15336_, _03601_);
  and _66944_ (_15338_, _05254_, _04303_);
  nor _66945_ (_15339_, _15338_, _15230_);
  or _66946_ (_15340_, _15339_, _05886_);
  and _66947_ (_15341_, _15340_, _08364_);
  and _66948_ (_15342_, _15341_, _15337_);
  nor _66949_ (_15343_, _08364_, _03414_);
  or _66950_ (_15344_, _15343_, _11344_);
  or _66951_ (_15345_, _15344_, _15342_);
  or _66952_ (_15346_, _11343_, _08680_);
  and _66953_ (_15347_, _15346_, _08393_);
  and _66954_ (_15348_, _15347_, _15345_);
  and _66955_ (_15349_, _08392_, _08644_);
  or _66956_ (_15350_, _15349_, _03778_);
  or _66957_ (_15351_, _15350_, _15348_);
  or _66958_ (_15352_, _12333_, _03779_);
  and _66959_ (_15353_, _15352_, _07905_);
  nand _66960_ (_15354_, _15353_, _15351_);
  nand _66961_ (_15355_, _08753_, _07904_);
  and _66962_ (_15356_, _15355_, _07766_);
  and _66963_ (_15357_, _15356_, _15354_);
  or _66964_ (_15358_, _15357_, _15210_);
  and _66965_ (_15359_, _15358_, _07778_);
  nor _66966_ (_15360_, _15204_, _07778_);
  or _66967_ (_15361_, _15360_, _15103_);
  nor _66968_ (_15362_, _15361_, _15359_);
  or _66969_ (_15363_, _08678_, _04199_);
  and _66970_ (_15364_, _15363_, _08421_);
  or _66971_ (_15365_, _15364_, _15362_);
  and _66972_ (_15366_, _04058_, _03191_);
  not _66973_ (_15367_, _15366_);
  or _66974_ (_15368_, _08678_, _15367_);
  and _66975_ (_15369_, _15368_, _15365_);
  or _66976_ (_15370_, _15369_, _08420_);
  or _66977_ (_15371_, _08425_, _08642_);
  and _66978_ (_15372_, _15371_, _03789_);
  and _66979_ (_15373_, _15372_, _15370_);
  or _66980_ (_15374_, _12331_, _08429_);
  and _66981_ (_15375_, _15374_, _08431_);
  or _66982_ (_15376_, _15375_, _15373_);
  or _66983_ (_15377_, _08435_, _08750_);
  and _66984_ (_15378_, _15377_, _07777_);
  and _66985_ (_15379_, _15378_, _15376_);
  or _66986_ (_15380_, _15379_, _15207_);
  and _66987_ (_15381_, _15380_, _15121_);
  nor _66988_ (_15382_, _15121_, _08679_);
  or _66989_ (_15383_, _15382_, _15123_);
  or _66990_ (_15384_, _15383_, _15381_);
  nand _66991_ (_15385_, _15123_, _08679_);
  and _66992_ (_15386_, _15385_, _15128_);
  and _66993_ (_15387_, _15386_, _15384_);
  nor _66994_ (_15388_, _08679_, _15128_);
  or _66995_ (_15389_, _15388_, _08450_);
  or _66996_ (_15390_, _15389_, _15387_);
  nand _66997_ (_15391_, _08450_, _08643_);
  and _66998_ (_15392_, _15391_, _03784_);
  and _66999_ (_15393_, _15392_, _15390_);
  nor _67000_ (_15394_, _12332_, _03784_);
  or _67001_ (_15395_, _15394_, _08458_);
  or _67002_ (_15396_, _15395_, _15393_);
  nand _67003_ (_15397_, _08458_, _08752_);
  and _67004_ (_15398_, _15397_, _15396_);
  or _67005_ (_15399_, _15398_, _03624_);
  nor _67006_ (_15400_, _12326_, _07908_);
  or _67007_ (_15401_, _15400_, _15204_);
  or _67008_ (_15402_, _15401_, _07795_);
  and _67009_ (_15403_, _15402_, _07898_);
  and _67010_ (_15404_, _15403_, _15399_);
  and _67011_ (_15405_, _07875_, _07870_);
  nor _67012_ (_15406_, _15405_, _07876_);
  and _67013_ (_15407_, _15406_, _08468_);
  or _67014_ (_15408_, _15407_, _08475_);
  or _67015_ (_15409_, _15408_, _15404_);
  and _67016_ (_15410_, _08487_, _08485_);
  nor _67017_ (_15411_, _15410_, _08488_);
  or _67018_ (_15412_, _15411_, _08477_);
  and _67019_ (_15413_, _15412_, _03777_);
  and _67020_ (_15414_, _15413_, _15409_);
  and _67021_ (_15415_, _08568_, _08564_);
  nor _67022_ (_15416_, _15415_, _08569_);
  and _67023_ (_15417_, _15416_, _03776_);
  or _67024_ (_15418_, _15417_, _15414_);
  and _67025_ (_15419_, _15418_, _08589_);
  and _67026_ (_15420_, _08598_, _07972_);
  nor _67027_ (_15421_, _15420_, _08599_);
  and _67028_ (_15422_, _15421_, _08506_);
  or _67029_ (_15423_, _15422_, _08587_);
  or _67030_ (_15424_, _15423_, _15419_);
  nand _67031_ (_15425_, _08587_, _03335_);
  and _67032_ (_15426_, _15425_, _08617_);
  and _67033_ (_15427_, _15426_, _15424_);
  nor _67034_ (_15428_, _08681_, _08680_);
  nor _67035_ (_15429_, _15428_, _08682_);
  and _67036_ (_15430_, _15429_, _08618_);
  or _67037_ (_15431_, _15430_, _08620_);
  or _67038_ (_15432_, _15431_, _15427_);
  and _67039_ (_15433_, _15432_, _15203_);
  or _67040_ (_15434_, _15433_, _03517_);
  and _67041_ (_15435_, _08711_, _08316_);
  nor _67042_ (_15436_, _15435_, _08712_);
  or _67043_ (_15437_, _15436_, _03518_);
  and _67044_ (_15438_, _15437_, _08734_);
  and _67045_ (_15439_, _15438_, _15434_);
  nor _67046_ (_15440_, _08753_, _08751_);
  nor _67047_ (_15441_, _15440_, _08754_);
  and _67048_ (_15442_, _15441_, _08701_);
  or _67049_ (_15443_, _15442_, _08732_);
  or _67050_ (_15444_, _15443_, _15439_);
  and _67051_ (_15445_, _15444_, _15200_);
  or _67052_ (_15446_, _15445_, _03815_);
  or _67053_ (_15447_, _15232_, _04246_);
  and _67054_ (_15448_, _15447_, _08776_);
  and _67055_ (_15449_, _15448_, _15446_);
  nor _67056_ (_15450_, _08806_, _08781_);
  nor _67057_ (_15451_, _15450_, _08776_);
  or _67058_ (_15452_, _15451_, _08780_);
  or _67059_ (_15453_, _15452_, _15449_);
  nand _67060_ (_15454_, _08780_, _07584_);
  and _67061_ (_15455_, _15454_, _03823_);
  and _67062_ (_15456_, _15455_, _15453_);
  nor _67063_ (_15457_, _15263_, _03823_);
  or _67064_ (_15458_, _15457_, _03447_);
  or _67065_ (_15459_, _15458_, _15456_);
  nor _67066_ (_15460_, _15231_, _15204_);
  nand _67067_ (_15461_, _15460_, _03447_);
  and _67068_ (_15462_, _15461_, _08799_);
  and _67069_ (_15463_, _15462_, _15459_);
  and _67070_ (_15464_, _15450_, _08798_);
  or _67071_ (_15465_, _15464_, _08805_);
  or _67072_ (_15466_, _15465_, _15463_);
  nand _67073_ (_15467_, _08805_, _07584_);
  and _67074_ (_15468_, _15467_, _43000_);
  and _67075_ (_15469_, _15468_, _15466_);
  or _67076_ (_15470_, _15469_, _15199_);
  and _67077_ (_43492_, _15470_, _41806_);
  nor _67078_ (_15471_, _43000_, _07584_);
  nor _67079_ (_15472_, _05254_, _07584_);
  and _67080_ (_15473_, _12533_, _05254_);
  nor _67081_ (_15474_, _15473_, _15472_);
  nand _67082_ (_15475_, _15474_, _03600_);
  not _67083_ (_15476_, _04182_);
  or _67084_ (_15477_, _08640_, _15476_);
  and _67085_ (_15478_, _04058_, _03181_);
  nand _67086_ (_15479_, _03904_, _03216_);
  nor _67087_ (_15480_, _07908_, _04875_);
  nor _67088_ (_15481_, _15480_, _15472_);
  nand _67089_ (_15482_, _15481_, _07390_);
  nand _67090_ (_15483_, _08064_, _04875_);
  or _67091_ (_15484_, _14975_, _06637_);
  nor _67092_ (_15485_, _08078_, _04875_);
  nor _67093_ (_15486_, _04064_, _07584_);
  and _67094_ (_15487_, _04064_, _07584_);
  or _67095_ (_15488_, _15487_, _15486_);
  and _67096_ (_15489_, _15488_, _08078_);
  or _67097_ (_15490_, _15489_, _08066_);
  or _67098_ (_15491_, _15490_, _15485_);
  and _67099_ (_15492_, _15491_, _03235_);
  or _67100_ (_15493_, _15492_, _04422_);
  and _67101_ (_15494_, _15493_, _15484_);
  and _67102_ (_15495_, _15494_, _04081_);
  nor _67103_ (_15496_, _12416_, _07908_);
  nor _67104_ (_15497_, _15496_, _15472_);
  nor _67105_ (_15498_, _15497_, _04081_);
  or _67106_ (_15499_, _15498_, _08089_);
  or _67107_ (_15500_, _15499_, _15495_);
  nand _67108_ (_15501_, _15236_, \oc8051_golden_model_1.ACC [2]);
  and _67109_ (_15502_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor _67110_ (_15503_, _15502_, _08095_);
  or _67111_ (_15504_, _15503_, _15236_);
  and _67112_ (_15505_, _15504_, _15501_);
  nand _67113_ (_15506_, _15505_, _08089_);
  and _67114_ (_15507_, _15506_, _03730_);
  and _67115_ (_15508_, _15507_, _15500_);
  nor _67116_ (_15509_, _05903_, _07584_);
  and _67117_ (_15510_, _12411_, _05903_);
  nor _67118_ (_15511_, _15510_, _15509_);
  nor _67119_ (_15512_, _15511_, _04055_);
  nor _67120_ (_15513_, _15481_, _03996_);
  or _67121_ (_15514_, _15513_, _08064_);
  or _67122_ (_15515_, _15514_, _15512_);
  or _67123_ (_15516_, _15515_, _15508_);
  and _67124_ (_15517_, _15516_, _15483_);
  or _67125_ (_15518_, _15517_, _04443_);
  or _67126_ (_15519_, _06637_, _08128_);
  and _67127_ (_15520_, _15519_, _03737_);
  and _67128_ (_15521_, _15520_, _15518_);
  nor _67129_ (_15522_, _08260_, _03737_);
  or _67130_ (_15523_, _15522_, _08132_);
  or _67131_ (_15524_, _15523_, _15521_);
  nand _67132_ (_15525_, _08132_, _07433_);
  and _67133_ (_15526_, _15525_, _15524_);
  or _67134_ (_15527_, _15526_, _03714_);
  and _67135_ (_15528_, _12409_, _05903_);
  nor _67136_ (_15529_, _15528_, _15509_);
  nand _67137_ (_15530_, _15529_, _03714_);
  and _67138_ (_15531_, _15530_, _06840_);
  and _67139_ (_15532_, _15531_, _15527_);
  and _67140_ (_15533_, _15510_, _12443_);
  nor _67141_ (_15534_, _15533_, _15509_);
  nor _67142_ (_15535_, _15534_, _06840_);
  or _67143_ (_15536_, _15535_, _06869_);
  or _67144_ (_15537_, _15536_, _15532_);
  nor _67145_ (_15538_, _07333_, _07331_);
  nor _67146_ (_15539_, _15538_, _07334_);
  or _67147_ (_15540_, _15539_, _06875_);
  and _67148_ (_15541_, _15540_, _15537_);
  or _67149_ (_15542_, _15541_, _08060_);
  and _67150_ (_15543_, _04406_, \oc8051_golden_model_1.ACC [1]);
  and _67151_ (_15544_, _04620_, _03335_);
  nor _67152_ (_15545_, _15544_, _08680_);
  nor _67153_ (_15546_, _15545_, _15543_);
  nor _67154_ (_15547_, _08676_, _15546_);
  and _67155_ (_15548_, _08676_, _15546_);
  nor _67156_ (_15549_, _15548_, _15547_);
  nor _67157_ (_15550_, _15072_, _08680_);
  not _67158_ (_15551_, _15550_);
  or _67159_ (_15552_, _15551_, _15549_);
  and _67160_ (_15553_, _15552_, \oc8051_golden_model_1.PSW [7]);
  nor _67161_ (_15554_, _15549_, \oc8051_golden_model_1.PSW [7]);
  or _67162_ (_15555_, _15554_, _15553_);
  nand _67163_ (_15556_, _15551_, _15549_);
  and _67164_ (_15557_, _15556_, _15555_);
  nor _67165_ (_15558_, _15557_, _08051_);
  or _67166_ (_15559_, _15558_, _11350_);
  and _67167_ (_15560_, _15559_, _15542_);
  nor _67168_ (_15561_, _06501_, _03274_);
  and _67169_ (_15562_, _06546_, _03335_);
  nor _67170_ (_15563_, _15562_, _08644_);
  nor _67171_ (_15564_, _15563_, _15561_);
  nor _67172_ (_15565_, _08640_, _15564_);
  and _67173_ (_15566_, _08640_, _15564_);
  nor _67174_ (_15567_, _15566_, _15565_);
  nor _67175_ (_15568_, _15083_, _08644_);
  and _67176_ (_15569_, _15568_, \oc8051_golden_model_1.PSW [7]);
  not _67177_ (_15570_, _15569_);
  nor _67178_ (_15571_, _15570_, _15567_);
  and _67179_ (_15572_, _15570_, _15567_);
  nor _67180_ (_15573_, _15572_, _15571_);
  nor _67181_ (_15574_, _15573_, _10201_);
  or _67182_ (_15575_, _15574_, _03761_);
  or _67183_ (_15576_, _15575_, _15560_);
  nor _67184_ (_15577_, _08290_, _08288_);
  nor _67185_ (_15578_, _15577_, _08291_);
  and _67186_ (_15579_, _08319_, \oc8051_golden_model_1.PSW [7]);
  not _67187_ (_15580_, _15579_);
  nor _67188_ (_15581_, _15580_, _15578_);
  and _67189_ (_15582_, _15580_, _15578_);
  nor _67190_ (_15583_, _15582_, _15581_);
  nand _67191_ (_15584_, _15583_, _03761_);
  and _67192_ (_15585_, _15584_, _07914_);
  and _67193_ (_15586_, _15585_, _15576_);
  nor _67194_ (_15587_, _04048_, \oc8051_golden_model_1.ACC [0]);
  nor _67195_ (_15588_, _08753_, _15587_);
  nor _67196_ (_15589_, _15588_, _10033_);
  nor _67197_ (_15590_, _08748_, _15589_);
  and _67198_ (_15591_, _08748_, _15589_);
  nor _67199_ (_15592_, _15591_, _15590_);
  not _67200_ (_15593_, _10059_);
  or _67201_ (_15594_, _15593_, _15592_);
  and _67202_ (_15595_, _15594_, \oc8051_golden_model_1.PSW [7]);
  nor _67203_ (_15596_, _15592_, \oc8051_golden_model_1.PSW [7]);
  or _67204_ (_15597_, _15596_, _15595_);
  nand _67205_ (_15598_, _15593_, _15592_);
  and _67206_ (_15599_, _15598_, _15597_);
  nor _67207_ (_15600_, _15599_, _07914_);
  or _67208_ (_15601_, _15600_, _07912_);
  or _67209_ (_15602_, _15601_, _15586_);
  nand _67210_ (_15603_, _03904_, _07912_);
  and _67211_ (_15604_, _15603_, _03710_);
  and _67212_ (_15605_, _15604_, _15602_);
  nor _67213_ (_15606_, _12461_, _08339_);
  nor _67214_ (_15607_, _15606_, _15509_);
  nor _67215_ (_15608_, _15607_, _03710_);
  or _67216_ (_15609_, _15608_, _07390_);
  or _67217_ (_15610_, _15609_, _15605_);
  and _67218_ (_15611_, _15610_, _15482_);
  or _67219_ (_15612_, _15611_, _04481_);
  and _67220_ (_15613_, _06637_, _05254_);
  nor _67221_ (_15614_, _15613_, _15472_);
  nand _67222_ (_15615_, _15614_, _04481_);
  and _67223_ (_15616_, _15615_, _03589_);
  and _67224_ (_15617_, _15616_, _15612_);
  nor _67225_ (_15618_, _12519_, _07908_);
  nor _67226_ (_15619_, _15618_, _15472_);
  nor _67227_ (_15620_, _15619_, _03589_);
  or _67228_ (_15621_, _15620_, _07405_);
  or _67229_ (_15622_, _15621_, _15617_);
  or _67230_ (_15623_, _07604_, _07411_);
  and _67231_ (_15624_, _15623_, _15622_);
  or _67232_ (_15626_, _15624_, _03216_);
  and _67233_ (_15627_, _15626_, _15479_);
  or _67234_ (_15628_, _15627_, _03601_);
  and _67235_ (_15629_, _05254_, _06332_);
  nor _67236_ (_15630_, _15629_, _15472_);
  nand _67237_ (_15631_, _15630_, _03601_);
  and _67238_ (_15632_, _15631_, _08364_);
  and _67239_ (_15633_, _15632_, _15628_);
  nor _67240_ (_15634_, _08364_, _03904_);
  or _67241_ (_15635_, _15634_, _08371_);
  or _67242_ (_15637_, _15635_, _15633_);
  or _67243_ (_15638_, _08377_, _08676_);
  and _67244_ (_15639_, _15638_, _08383_);
  and _67245_ (_15640_, _15639_, _15637_);
  and _67246_ (_15641_, _04488_, _03181_);
  nor _67247_ (_15642_, _08383_, _08677_);
  or _67248_ (_15643_, _15642_, _15641_);
  or _67249_ (_15644_, _15643_, _15640_);
  nand _67250_ (_15645_, _15641_, _08677_);
  and _67251_ (_15646_, _15645_, _15644_);
  or _67252_ (_15648_, _15646_, _15478_);
  and _67253_ (_15649_, _03616_, _03181_);
  not _67254_ (_15650_, _15649_);
  not _67255_ (_15651_, _15478_);
  or _67256_ (_15652_, _08676_, _15651_);
  and _67257_ (_15653_, _15652_, _15650_);
  and _67258_ (_15654_, _15653_, _15648_);
  or _67259_ (_15655_, _08640_, _04182_);
  and _67260_ (_15656_, _15655_, _08392_);
  or _67261_ (_15657_, _15656_, _15654_);
  and _67262_ (_15659_, _15657_, _15477_);
  or _67263_ (_15660_, _15659_, _03778_);
  or _67264_ (_15661_, _12539_, _03779_);
  and _67265_ (_15662_, _15661_, _07905_);
  and _67266_ (_15663_, _15662_, _15660_);
  and _67267_ (_15664_, _08748_, _07904_);
  or _67268_ (_15665_, _15664_, _03600_);
  or _67269_ (_15666_, _15665_, _15663_);
  and _67270_ (_15667_, _15666_, _15475_);
  or _67271_ (_15668_, _15667_, _03780_);
  or _67272_ (_15670_, _15472_, _07778_);
  and _67273_ (_15671_, _15670_, _08417_);
  and _67274_ (_15672_, _15671_, _15668_);
  and _67275_ (_15673_, _08421_, _08674_);
  or _67276_ (_15674_, _15673_, _08420_);
  or _67277_ (_15675_, _15674_, _15672_);
  or _67278_ (_15676_, _08425_, _08638_);
  and _67279_ (_15677_, _15676_, _03789_);
  and _67280_ (_15678_, _15677_, _15675_);
  and _67281_ (_15679_, _12537_, _03788_);
  or _67282_ (_15681_, _15679_, _08429_);
  or _67283_ (_15682_, _15681_, _15678_);
  or _67284_ (_15683_, _08435_, _08746_);
  and _67285_ (_15684_, _15683_, _07777_);
  and _67286_ (_15685_, _15684_, _15682_);
  not _67287_ (_15686_, _11332_);
  or _67288_ (_15687_, _15630_, _12538_);
  nor _67289_ (_15688_, _15687_, _07777_);
  or _67290_ (_15689_, _15688_, _15686_);
  or _67291_ (_15690_, _15689_, _15685_);
  nor _67292_ (_15692_, _08675_, _11333_);
  or _67293_ (_15693_, _15692_, _08447_);
  and _67294_ (_15694_, _15693_, _15690_);
  not _67295_ (_15695_, _11333_);
  nor _67296_ (_15696_, _08675_, _15695_);
  or _67297_ (_15697_, _15696_, _08450_);
  or _67298_ (_15698_, _15697_, _15694_);
  nand _67299_ (_15699_, _08450_, _08639_);
  and _67300_ (_15700_, _15699_, _03784_);
  and _67301_ (_15701_, _15700_, _15698_);
  nor _67302_ (_15703_, _12538_, _03784_);
  or _67303_ (_15704_, _15703_, _08458_);
  or _67304_ (_15705_, _15704_, _15701_);
  nand _67305_ (_15706_, _08458_, _08747_);
  and _67306_ (_15707_, _15706_, _15705_);
  or _67307_ (_15708_, _15707_, _03624_);
  nor _67308_ (_15709_, _12532_, _07908_);
  nor _67309_ (_15710_, _15709_, _15472_);
  nand _67310_ (_15711_, _15710_, _03624_);
  and _67311_ (_15712_, _15711_, _07898_);
  and _67312_ (_15714_, _15712_, _15708_);
  and _67313_ (_15715_, _07877_, _07863_);
  nor _67314_ (_15716_, _15715_, _07878_);
  and _67315_ (_15717_, _15716_, _08468_);
  or _67316_ (_15718_, _15717_, _15714_);
  and _67317_ (_15719_, _15718_, _08477_);
  and _67318_ (_15720_, _08489_, _08027_);
  nor _67319_ (_15721_, _15720_, _08490_);
  and _67320_ (_15722_, _15721_, _08475_);
  or _67321_ (_15723_, _15722_, _03776_);
  or _67322_ (_15725_, _15723_, _15719_);
  and _67323_ (_15726_, _08570_, _08558_);
  nor _67324_ (_15727_, _15726_, _08571_);
  or _67325_ (_15728_, _15727_, _03777_);
  and _67326_ (_15729_, _15728_, _08589_);
  and _67327_ (_15730_, _15729_, _15725_);
  and _67328_ (_15731_, _08600_, _07953_);
  nor _67329_ (_15732_, _15731_, _08601_);
  and _67330_ (_15733_, _15732_, _08506_);
  or _67331_ (_15734_, _15733_, _08587_);
  or _67332_ (_15736_, _15734_, _15730_);
  nand _67333_ (_15737_, _08587_, _03274_);
  and _67334_ (_15738_, _15737_, _08617_);
  and _67335_ (_15739_, _15738_, _15736_);
  and _67336_ (_15740_, _08683_, _08677_);
  nor _67337_ (_15741_, _15740_, _08684_);
  and _67338_ (_15742_, _15741_, _08618_);
  or _67339_ (_15743_, _15742_, _08620_);
  or _67340_ (_15744_, _15743_, _15739_);
  and _67341_ (_15745_, _08647_, _08641_);
  nor _67342_ (_15747_, _15745_, _08648_);
  or _67343_ (_15748_, _15747_, _08624_);
  and _67344_ (_15749_, _15748_, _03518_);
  and _67345_ (_15750_, _15749_, _15744_);
  and _67346_ (_15751_, _08713_, _08290_);
  nor _67347_ (_15752_, _15751_, _08714_);
  or _67348_ (_15753_, _15752_, _08701_);
  and _67349_ (_15754_, _15753_, _08703_);
  or _67350_ (_15755_, _15754_, _15750_);
  and _67351_ (_15756_, _08755_, _08749_);
  nor _67352_ (_15758_, _15756_, _08756_);
  or _67353_ (_15759_, _15758_, _08734_);
  and _67354_ (_15760_, _15759_, _08733_);
  and _67355_ (_15761_, _15760_, _15755_);
  and _67356_ (_15762_, _08732_, \oc8051_golden_model_1.ACC [1]);
  or _67357_ (_15763_, _15762_, _03815_);
  or _67358_ (_15764_, _15763_, _15761_);
  nand _67359_ (_15765_, _15497_, _03815_);
  and _67360_ (_15766_, _15765_, _08776_);
  and _67361_ (_15767_, _15766_, _15764_);
  and _67362_ (_15769_, _08095_, _03335_);
  nor _67363_ (_15770_, _08781_, _07584_);
  or _67364_ (_15771_, _15770_, _15769_);
  and _67365_ (_15772_, _15771_, _08775_);
  or _67366_ (_15773_, _15772_, _08780_);
  or _67367_ (_15774_, _15773_, _15767_);
  nand _67368_ (_15775_, _08780_, _07578_);
  and _67369_ (_15776_, _15775_, _03823_);
  and _67370_ (_15777_, _15776_, _15774_);
  nor _67371_ (_15778_, _15529_, _03823_);
  or _67372_ (_15780_, _15778_, _03447_);
  or _67373_ (_15781_, _15780_, _15777_);
  and _67374_ (_15782_, _12592_, _05254_);
  nor _67375_ (_15783_, _15782_, _15472_);
  nand _67376_ (_15784_, _15783_, _03447_);
  and _67377_ (_15785_, _15784_, _08799_);
  and _67378_ (_15786_, _15785_, _15781_);
  and _67379_ (_15787_, _08806_, \oc8051_golden_model_1.ACC [2]);
  nor _67380_ (_15788_, _08806_, \oc8051_golden_model_1.ACC [2]);
  nor _67381_ (_15789_, _15788_, _15787_);
  nor _67382_ (_15791_, _15789_, _08805_);
  nor _67383_ (_15792_, _15791_, _11964_);
  or _67384_ (_15793_, _15792_, _15786_);
  nand _67385_ (_15794_, _08805_, _07578_);
  and _67386_ (_15795_, _15794_, _43000_);
  and _67387_ (_15796_, _15795_, _15793_);
  or _67388_ (_15797_, _15796_, _15471_);
  and _67389_ (_43493_, _15797_, _41806_);
  nor _67390_ (_15798_, _43000_, _07578_);
  nor _67391_ (_15799_, _08673_, _08671_);
  nor _67392_ (_15800_, _08685_, _15799_);
  and _67393_ (_15801_, _08685_, _15799_);
  nor _67394_ (_15802_, _15801_, _15800_);
  nand _67395_ (_15803_, _15802_, _08618_);
  and _67396_ (_15804_, _07879_, _07857_);
  nor _67397_ (_15805_, _15804_, _07880_);
  or _67398_ (_15806_, _15805_, _07898_);
  nand _67399_ (_15807_, _15686_, _08673_);
  and _67400_ (_15808_, _15807_, _15695_);
  or _67401_ (_15809_, _14962_, _08671_);
  nor _67402_ (_15811_, _05254_, _07578_);
  and _67403_ (_15812_, _12733_, _05254_);
  nor _67404_ (_15813_, _15812_, _15811_);
  nand _67405_ (_15814_, _15813_, _03600_);
  nor _67406_ (_15815_, _08364_, _03581_);
  nand _67407_ (_15816_, _03581_, _03216_);
  nor _67408_ (_15817_, _07908_, _05005_);
  nor _67409_ (_15818_, _15817_, _15811_);
  nand _67410_ (_15819_, _15818_, _07390_);
  and _67411_ (_15820_, _03904_, \oc8051_golden_model_1.ACC [2]);
  nor _67412_ (_15822_, _15590_, _15820_);
  nor _67413_ (_15823_, _10030_, _15822_);
  and _67414_ (_15824_, _10030_, _15822_);
  nor _67415_ (_15825_, _15824_, _15823_);
  and _67416_ (_15826_, _15825_, \oc8051_golden_model_1.PSW [7]);
  nor _67417_ (_15827_, _15825_, \oc8051_golden_model_1.PSW [7]);
  nor _67418_ (_15828_, _15827_, _15826_);
  and _67419_ (_15829_, _15828_, _15595_);
  nor _67420_ (_15830_, _15828_, _15595_);
  or _67421_ (_15831_, _15830_, _15829_);
  nand _67422_ (_15833_, _15831_, _07913_);
  nor _67423_ (_15834_, _05903_, _07578_);
  and _67424_ (_15835_, _12631_, _05903_);
  and _67425_ (_15836_, _15835_, _12648_);
  nor _67426_ (_15837_, _15836_, _15834_);
  nor _67427_ (_15838_, _15837_, _06840_);
  nand _67428_ (_15839_, _08064_, _05005_);
  or _67429_ (_15840_, _14975_, _06592_);
  nand _67430_ (_15841_, _08079_, _05005_);
  nor _67431_ (_15842_, _04064_, _07578_);
  and _67432_ (_15844_, _04064_, _07578_);
  nor _67433_ (_15845_, _15844_, _15842_);
  nand _67434_ (_15846_, _15845_, _08078_);
  and _67435_ (_15847_, _15846_, _15841_);
  or _67436_ (_15848_, _15847_, _08066_);
  and _67437_ (_15849_, _15848_, _03235_);
  or _67438_ (_15850_, _15849_, _04422_);
  and _67439_ (_15851_, _15850_, _04081_);
  and _67440_ (_15852_, _15851_, _15840_);
  nor _67441_ (_15853_, _12627_, _07908_);
  nor _67442_ (_15855_, _15853_, _15811_);
  nor _67443_ (_15856_, _15855_, _04081_);
  or _67444_ (_15857_, _15856_, _08089_);
  or _67445_ (_15858_, _15857_, _15852_);
  not _67446_ (_15859_, \oc8051_golden_model_1.PSW [6]);
  nor _67447_ (_15860_, _08095_, _15859_);
  nor _67448_ (_15861_, _15860_, \oc8051_golden_model_1.ACC [3]);
  or _67449_ (_15862_, _15861_, _08096_);
  nand _67450_ (_15863_, _15862_, _08089_);
  and _67451_ (_15864_, _15863_, _15858_);
  or _67452_ (_15866_, _15864_, _03715_);
  nor _67453_ (_15867_, _15835_, _15834_);
  nand _67454_ (_15868_, _15867_, _03715_);
  and _67455_ (_15869_, _15868_, _03996_);
  and _67456_ (_15870_, _15869_, _15866_);
  nor _67457_ (_15871_, _15818_, _03996_);
  or _67458_ (_15872_, _15871_, _08064_);
  or _67459_ (_15873_, _15872_, _15870_);
  and _67460_ (_15874_, _15873_, _15839_);
  or _67461_ (_15875_, _15874_, _04443_);
  or _67462_ (_15877_, _06592_, _08128_);
  and _67463_ (_15878_, _15877_, _03737_);
  and _67464_ (_15879_, _15878_, _15875_);
  nor _67465_ (_15880_, _08248_, _03737_);
  or _67466_ (_15881_, _15880_, _08132_);
  or _67467_ (_15882_, _15881_, _15879_);
  nand _67468_ (_15883_, _08132_, _06075_);
  and _67469_ (_15884_, _15883_, _15882_);
  or _67470_ (_15885_, _15884_, _03714_);
  and _67471_ (_15886_, _12641_, _05903_);
  nor _67472_ (_15888_, _15886_, _15834_);
  nand _67473_ (_15889_, _15888_, _03714_);
  and _67474_ (_15890_, _15889_, _06840_);
  and _67475_ (_15891_, _15890_, _15885_);
  or _67476_ (_15892_, _15891_, _15838_);
  and _67477_ (_15893_, _15892_, _06875_);
  nor _67478_ (_15894_, _07336_, _07334_);
  nor _67479_ (_15895_, _15894_, _07337_);
  nand _67480_ (_15896_, _15895_, _06869_);
  nand _67481_ (_15897_, _15896_, _08059_);
  or _67482_ (_15899_, _15897_, _15893_);
  and _67483_ (_15900_, _04875_, \oc8051_golden_model_1.ACC [2]);
  nor _67484_ (_15901_, _15547_, _15900_);
  nor _67485_ (_15902_, _15799_, _15901_);
  and _67486_ (_15903_, _15799_, _15901_);
  nor _67487_ (_15904_, _15903_, _15902_);
  and _67488_ (_15905_, _15904_, \oc8051_golden_model_1.PSW [7]);
  nor _67489_ (_15906_, _15904_, \oc8051_golden_model_1.PSW [7]);
  nor _67490_ (_15907_, _15906_, _15905_);
  and _67491_ (_15908_, _15907_, _15553_);
  nor _67492_ (_15910_, _15907_, _15553_);
  or _67493_ (_15911_, _15910_, _15908_);
  nand _67494_ (_15912_, _15911_, _08060_);
  and _67495_ (_15913_, _15912_, _15899_);
  or _67496_ (_15914_, _15913_, _08051_);
  not _67497_ (_15915_, _15568_);
  or _67498_ (_15916_, _15915_, _15567_);
  and _67499_ (_15917_, _15916_, \oc8051_golden_model_1.PSW [7]);
  nor _67500_ (_15918_, _06637_, _07584_);
  nor _67501_ (_15919_, _15565_, _15918_);
  nor _67502_ (_15921_, _08637_, _08635_);
  nor _67503_ (_15922_, _15921_, _15919_);
  and _67504_ (_15923_, _15921_, _15919_);
  nor _67505_ (_15924_, _15923_, _15922_);
  and _67506_ (_15925_, _15924_, \oc8051_golden_model_1.PSW [7]);
  nor _67507_ (_15926_, _15924_, \oc8051_golden_model_1.PSW [7]);
  nor _67508_ (_15927_, _15926_, _15925_);
  and _67509_ (_15928_, _15927_, _15917_);
  nor _67510_ (_15929_, _15927_, _15917_);
  or _67511_ (_15930_, _15929_, _15928_);
  nand _67512_ (_15932_, _15930_, _08051_);
  and _67513_ (_15933_, _15932_, _03766_);
  and _67514_ (_15934_, _15933_, _15914_);
  nor _67515_ (_15935_, _08314_, _08292_);
  and _67516_ (_15936_, _08314_, _08292_);
  or _67517_ (_15937_, _15936_, _15935_);
  not _67518_ (_15938_, _15581_);
  and _67519_ (_15939_, _15938_, _15937_);
  nor _67520_ (_15940_, _15939_, _08321_);
  nand _67521_ (_15941_, _15940_, _07914_);
  and _67522_ (_15943_, _15941_, _08187_);
  or _67523_ (_15944_, _15943_, _15934_);
  and _67524_ (_15945_, _15944_, _15833_);
  or _67525_ (_15946_, _15945_, _07912_);
  nand _67526_ (_15947_, _03581_, _07912_);
  and _67527_ (_15948_, _15947_, _03710_);
  and _67528_ (_15949_, _15948_, _15946_);
  nor _67529_ (_15950_, _12612_, _08339_);
  nor _67530_ (_15951_, _15950_, _15834_);
  nor _67531_ (_15952_, _15951_, _03710_);
  or _67532_ (_15954_, _15952_, _07390_);
  or _67533_ (_15955_, _15954_, _15949_);
  and _67534_ (_15956_, _15955_, _15819_);
  or _67535_ (_15957_, _15956_, _04481_);
  and _67536_ (_15958_, _06592_, _05254_);
  nor _67537_ (_15959_, _15958_, _15811_);
  nand _67538_ (_15960_, _15959_, _04481_);
  and _67539_ (_15961_, _15960_, _03589_);
  and _67540_ (_15962_, _15961_, _15957_);
  nor _67541_ (_15963_, _12718_, _07908_);
  nor _67542_ (_15965_, _15963_, _15811_);
  nor _67543_ (_15966_, _15965_, _03589_);
  or _67544_ (_15967_, _15966_, _07405_);
  or _67545_ (_15968_, _15967_, _15962_);
  or _67546_ (_15969_, _07547_, _07411_);
  and _67547_ (_15970_, _15969_, _15968_);
  or _67548_ (_15971_, _15970_, _03216_);
  and _67549_ (_15972_, _15971_, _15816_);
  or _67550_ (_15973_, _15972_, _03601_);
  and _67551_ (_15974_, _05254_, _06276_);
  nor _67552_ (_15976_, _15974_, _15811_);
  nand _67553_ (_15977_, _15976_, _03601_);
  and _67554_ (_15978_, _15977_, _08364_);
  and _67555_ (_15979_, _15978_, _15973_);
  or _67556_ (_15980_, _15979_, _15815_);
  and _67557_ (_15981_, _15980_, _11343_);
  and _67558_ (_15982_, _11344_, _15799_);
  or _67559_ (_15983_, _15982_, _15981_);
  and _67560_ (_15984_, _15983_, _08393_);
  and _67561_ (_15985_, _08392_, _15921_);
  or _67562_ (_15987_, _15985_, _03778_);
  or _67563_ (_15988_, _15987_, _15984_);
  or _67564_ (_15989_, _12739_, _03779_);
  and _67565_ (_15990_, _15989_, _07905_);
  and _67566_ (_15991_, _15990_, _15988_);
  and _67567_ (_15992_, _10030_, _07904_);
  or _67568_ (_15993_, _15992_, _03600_);
  or _67569_ (_15994_, _15993_, _15991_);
  and _67570_ (_15995_, _15994_, _15814_);
  or _67571_ (_15996_, _15995_, _03780_);
  or _67572_ (_15998_, _15811_, _07778_);
  and _67573_ (_15999_, _15998_, _15096_);
  and _67574_ (_16000_, _15999_, _15996_);
  or _67575_ (_16001_, _15100_, _08671_);
  and _67576_ (_16002_, _16001_, _15103_);
  or _67577_ (_16003_, _16002_, _04199_);
  or _67578_ (_16004_, _16003_, _16000_);
  and _67579_ (_16005_, _16004_, _15809_);
  or _67580_ (_16006_, _16005_, _08420_);
  or _67581_ (_16007_, _08425_, _08635_);
  and _67582_ (_16009_, _16007_, _03789_);
  and _67583_ (_16010_, _16009_, _16006_);
  or _67584_ (_16011_, _12737_, _08429_);
  and _67585_ (_16012_, _16011_, _08431_);
  or _67586_ (_16013_, _16012_, _16010_);
  or _67587_ (_16014_, _08435_, _08744_);
  and _67588_ (_16015_, _16014_, _07777_);
  and _67589_ (_16016_, _16015_, _16013_);
  or _67590_ (_16017_, _15976_, _12738_);
  nor _67591_ (_16018_, _16017_, _07777_);
  or _67592_ (_16020_, _16018_, _15686_);
  or _67593_ (_16021_, _16020_, _16016_);
  and _67594_ (_16022_, _16021_, _15808_);
  nor _67595_ (_16023_, _08673_, _15695_);
  or _67596_ (_16024_, _16023_, _08450_);
  or _67597_ (_16025_, _16024_, _16022_);
  nand _67598_ (_16026_, _08450_, _08637_);
  and _67599_ (_16027_, _16026_, _03784_);
  and _67600_ (_16028_, _16027_, _16025_);
  nand _67601_ (_16029_, _12738_, _08461_);
  and _67602_ (_16031_, _16029_, _08460_);
  or _67603_ (_16032_, _16031_, _16028_);
  nand _67604_ (_16033_, _08458_, _08745_);
  and _67605_ (_16034_, _16033_, _07795_);
  and _67606_ (_16035_, _16034_, _16032_);
  nor _67607_ (_16036_, _12732_, _07908_);
  nor _67608_ (_16037_, _16036_, _15811_);
  nor _67609_ (_16038_, _16037_, _07795_);
  or _67610_ (_16039_, _16038_, _08468_);
  or _67611_ (_16040_, _16039_, _16035_);
  and _67612_ (_16042_, _16040_, _15806_);
  or _67613_ (_16043_, _16042_, _08475_);
  and _67614_ (_16044_, _08491_, _08022_);
  nor _67615_ (_16045_, _16044_, _08492_);
  or _67616_ (_16046_, _16045_, _08477_);
  and _67617_ (_16047_, _16046_, _03777_);
  and _67618_ (_16048_, _16047_, _16043_);
  and _67619_ (_16049_, _08572_, _08552_);
  nor _67620_ (_16050_, _16049_, _08573_);
  and _67621_ (_16051_, _16050_, _03776_);
  or _67622_ (_16053_, _16051_, _08506_);
  or _67623_ (_16054_, _16053_, _16048_);
  and _67624_ (_16055_, _08602_, _07948_);
  nor _67625_ (_16056_, _16055_, _08603_);
  or _67626_ (_16057_, _16056_, _08589_);
  and _67627_ (_16058_, _16057_, _08588_);
  and _67628_ (_16059_, _16058_, _16054_);
  and _67629_ (_16060_, _08587_, \oc8051_golden_model_1.ACC [2]);
  or _67630_ (_16061_, _16060_, _08618_);
  or _67631_ (_16062_, _16061_, _16059_);
  and _67632_ (_16064_, _16062_, _15803_);
  or _67633_ (_16065_, _16064_, _08620_);
  nor _67634_ (_16066_, _08649_, _15921_);
  and _67635_ (_16067_, _08649_, _15921_);
  nor _67636_ (_16068_, _16067_, _16066_);
  nand _67637_ (_16069_, _16068_, _08620_);
  and _67638_ (_16070_, _16069_, _03518_);
  and _67639_ (_16071_, _16070_, _16065_);
  nor _67640_ (_16072_, _08715_, _08314_);
  and _67641_ (_16073_, _08715_, _08314_);
  nor _67642_ (_16075_, _16073_, _16072_);
  and _67643_ (_16076_, _16075_, _03517_);
  or _67644_ (_16077_, _16076_, _08701_);
  or _67645_ (_16078_, _16077_, _16071_);
  nor _67646_ (_16079_, _08757_, _10030_);
  and _67647_ (_16080_, _08757_, _10030_);
  nor _67648_ (_16081_, _16080_, _16079_);
  nand _67649_ (_16082_, _16081_, _08701_);
  and _67650_ (_16083_, _16082_, _08733_);
  and _67651_ (_16084_, _16083_, _16078_);
  and _67652_ (_16086_, _08732_, \oc8051_golden_model_1.ACC [2]);
  or _67653_ (_16087_, _16086_, _03815_);
  or _67654_ (_16088_, _16087_, _16084_);
  nand _67655_ (_16089_, _15855_, _03815_);
  and _67656_ (_16090_, _16089_, _08776_);
  and _67657_ (_16091_, _16090_, _16088_);
  nor _67658_ (_16092_, _15769_, _07578_);
  or _67659_ (_16093_, _16092_, _08782_);
  and _67660_ (_16094_, _16093_, _08775_);
  or _67661_ (_16095_, _16094_, _08780_);
  or _67662_ (_16097_, _16095_, _16091_);
  nand _67663_ (_16098_, _08780_, _07484_);
  and _67664_ (_16099_, _16098_, _03823_);
  and _67665_ (_16100_, _16099_, _16097_);
  nor _67666_ (_16101_, _15888_, _03823_);
  or _67667_ (_16102_, _16101_, _03447_);
  or _67668_ (_16103_, _16102_, _16100_);
  and _67669_ (_16104_, _12794_, _05254_);
  nor _67670_ (_16105_, _16104_, _15811_);
  nand _67671_ (_16106_, _16105_, _03447_);
  and _67672_ (_16108_, _16106_, _08799_);
  and _67673_ (_16109_, _16108_, _16103_);
  or _67674_ (_16110_, _15787_, \oc8051_golden_model_1.ACC [3]);
  and _67675_ (_16111_, _16110_, _08807_);
  and _67676_ (_16112_, _16111_, _08798_);
  or _67677_ (_16113_, _16112_, _08805_);
  or _67678_ (_16114_, _16113_, _16109_);
  nand _67679_ (_16115_, _08805_, _07484_);
  and _67680_ (_16116_, _16115_, _43000_);
  and _67681_ (_16117_, _16116_, _16114_);
  or _67682_ (_16119_, _16117_, _15798_);
  and _67683_ (_43494_, _16119_, _41806_);
  nor _67684_ (_16120_, _43000_, _07484_);
  nand _67685_ (_16121_, _08732_, _07578_);
  nor _67686_ (_16122_, _05254_, _07484_);
  and _67687_ (_16123_, _12821_, _05254_);
  nor _67688_ (_16124_, _16123_, _16122_);
  nand _67689_ (_16125_, _16124_, _03600_);
  and _67690_ (_16126_, _08669_, _08381_);
  nor _67691_ (_16127_, _08364_, _03486_);
  nand _67692_ (_16129_, _03486_, _03216_);
  nor _67693_ (_16130_, _05777_, _07908_);
  nor _67694_ (_16131_, _16130_, _16122_);
  nand _67695_ (_16132_, _16131_, _07390_);
  and _67696_ (_16133_, _08322_, _08313_);
  nor _67697_ (_16134_, _16133_, _08323_);
  nand _67698_ (_16135_, _16134_, _03761_);
  and _67699_ (_16136_, _16135_, _07914_);
  or _67700_ (_16137_, _15928_, _15925_);
  and _67701_ (_16138_, _06592_, _07578_);
  or _67702_ (_16140_, _06592_, _07578_);
  and _67703_ (_16141_, _16140_, _15919_);
  or _67704_ (_16142_, _16141_, _16138_);
  nor _67705_ (_16143_, _08634_, _16142_);
  and _67706_ (_16144_, _08634_, _16142_);
  nor _67707_ (_16145_, _16144_, _16143_);
  and _67708_ (_16146_, _16145_, \oc8051_golden_model_1.PSW [7]);
  nor _67709_ (_16147_, _16145_, \oc8051_golden_model_1.PSW [7]);
  nor _67710_ (_16148_, _16147_, _16146_);
  and _67711_ (_16149_, _16148_, _16137_);
  nor _67712_ (_16151_, _16148_, _16137_);
  nor _67713_ (_16152_, _16151_, _16149_);
  and _67714_ (_16153_, _16152_, _08051_);
  nand _67715_ (_16154_, _08064_, _05777_);
  or _67716_ (_16155_, _08067_, _06730_);
  nor _67717_ (_16156_, _08078_, _05777_);
  or _67718_ (_16157_, _04064_, \oc8051_golden_model_1.ACC [4]);
  nand _67719_ (_16158_, _04064_, \oc8051_golden_model_1.ACC [4]);
  and _67720_ (_16159_, _16158_, _16157_);
  and _67721_ (_16160_, _16159_, _08078_);
  or _67722_ (_16162_, _16160_, _08066_);
  or _67723_ (_16163_, _16162_, _16156_);
  and _67724_ (_16164_, _16163_, _08069_);
  and _67725_ (_16165_, _16164_, _16155_);
  nor _67726_ (_16166_, _12841_, _07908_);
  nor _67727_ (_16167_, _16166_, _16122_);
  nor _67728_ (_16168_, _16167_, _04081_);
  or _67729_ (_16169_, _16168_, _08089_);
  or _67730_ (_16170_, _16169_, _16165_);
  nor _67731_ (_16171_, _08096_, \oc8051_golden_model_1.ACC [4]);
  or _67732_ (_16173_, _16171_, _08102_);
  nand _67733_ (_16174_, _16173_, _08089_);
  and _67734_ (_16175_, _16174_, _03730_);
  and _67735_ (_16176_, _16175_, _16170_);
  nor _67736_ (_16177_, _05903_, _07484_);
  and _67737_ (_16178_, _12845_, _05903_);
  nor _67738_ (_16179_, _16178_, _16177_);
  nor _67739_ (_16180_, _16179_, _04055_);
  nor _67740_ (_16181_, _16131_, _03996_);
  or _67741_ (_16182_, _16181_, _08064_);
  or _67742_ (_16184_, _16182_, _16180_);
  or _67743_ (_16185_, _16184_, _16176_);
  and _67744_ (_16186_, _16185_, _16154_);
  or _67745_ (_16187_, _16186_, _04443_);
  or _67746_ (_16188_, _06730_, _08128_);
  and _67747_ (_16189_, _16188_, _03737_);
  and _67748_ (_16190_, _16189_, _16187_);
  nor _67749_ (_16191_, _08235_, _03737_);
  or _67750_ (_16192_, _16191_, _08132_);
  or _67751_ (_16193_, _16192_, _16190_);
  nand _67752_ (_16195_, _08132_, _03335_);
  and _67753_ (_16196_, _16195_, _16193_);
  or _67754_ (_16197_, _16196_, _03714_);
  and _67755_ (_16198_, _12827_, _05903_);
  nor _67756_ (_16199_, _16198_, _16177_);
  nand _67757_ (_16200_, _16199_, _03714_);
  and _67758_ (_16201_, _16200_, _06840_);
  and _67759_ (_16202_, _16201_, _16197_);
  and _67760_ (_16203_, _16178_, _12860_);
  nor _67761_ (_16204_, _16203_, _16177_);
  nor _67762_ (_16206_, _16204_, _06840_);
  or _67763_ (_16207_, _16206_, _06869_);
  or _67764_ (_16208_, _16207_, _16202_);
  nor _67765_ (_16209_, _07339_, _07337_);
  nor _67766_ (_16210_, _16209_, _07340_);
  or _67767_ (_16211_, _16210_, _06875_);
  and _67768_ (_16212_, _16211_, _16208_);
  or _67769_ (_16213_, _16212_, _08060_);
  or _67770_ (_16214_, _15908_, _15905_);
  nor _67771_ (_16215_, _05005_, \oc8051_golden_model_1.ACC [3]);
  nand _67772_ (_16217_, _05005_, \oc8051_golden_model_1.ACC [3]);
  and _67773_ (_16218_, _16217_, _15901_);
  or _67774_ (_16219_, _16218_, _16215_);
  nor _67775_ (_16220_, _08669_, _16219_);
  and _67776_ (_16221_, _08669_, _16219_);
  nor _67777_ (_16222_, _16221_, _16220_);
  and _67778_ (_16223_, _16222_, \oc8051_golden_model_1.PSW [7]);
  nor _67779_ (_16224_, _16222_, \oc8051_golden_model_1.PSW [7]);
  nor _67780_ (_16225_, _16224_, _16223_);
  and _67781_ (_16226_, _16225_, _16214_);
  nor _67782_ (_16228_, _16225_, _16214_);
  nor _67783_ (_16229_, _16228_, _16226_);
  or _67784_ (_16230_, _16229_, _08059_);
  and _67785_ (_16231_, _16230_, _10201_);
  and _67786_ (_16232_, _16231_, _16213_);
  or _67787_ (_16233_, _16232_, _03761_);
  or _67788_ (_16234_, _16233_, _16153_);
  and _67789_ (_16235_, _16234_, _16136_);
  or _67790_ (_16236_, _15829_, _15826_);
  or _67791_ (_16237_, _15822_, _10039_);
  and _67792_ (_16239_, _16237_, _10038_);
  nor _67793_ (_16240_, _08743_, _16239_);
  and _67794_ (_16241_, _08743_, _16239_);
  nor _67795_ (_16242_, _16241_, _16240_);
  and _67796_ (_16243_, _16242_, \oc8051_golden_model_1.PSW [7]);
  nor _67797_ (_16244_, _16242_, \oc8051_golden_model_1.PSW [7]);
  nor _67798_ (_16245_, _16244_, _16243_);
  and _67799_ (_16246_, _16245_, _16236_);
  nor _67800_ (_16247_, _16245_, _16236_);
  nor _67801_ (_16248_, _16247_, _16246_);
  and _67802_ (_16250_, _16248_, _07913_);
  or _67803_ (_16251_, _16250_, _07912_);
  or _67804_ (_16252_, _16251_, _16235_);
  nand _67805_ (_16253_, _03486_, _07912_);
  and _67806_ (_16254_, _16253_, _03710_);
  and _67807_ (_16255_, _16254_, _16252_);
  nor _67808_ (_16256_, _12825_, _08339_);
  nor _67809_ (_16257_, _16256_, _16177_);
  nor _67810_ (_16258_, _16257_, _03710_);
  or _67811_ (_16259_, _16258_, _07390_);
  or _67812_ (_16261_, _16259_, _16255_);
  and _67813_ (_16262_, _16261_, _16132_);
  or _67814_ (_16263_, _16262_, _04481_);
  and _67815_ (_16264_, _06730_, _05254_);
  nor _67816_ (_16265_, _16264_, _16122_);
  nand _67817_ (_16266_, _16265_, _04481_);
  and _67818_ (_16267_, _16266_, _03589_);
  and _67819_ (_16268_, _16267_, _16263_);
  nor _67820_ (_16269_, _12933_, _07908_);
  nor _67821_ (_16270_, _16269_, _16122_);
  nor _67822_ (_16272_, _16270_, _03589_);
  or _67823_ (_16273_, _16272_, _07405_);
  or _67824_ (_16274_, _16273_, _16268_);
  or _67825_ (_16275_, _07493_, _07411_);
  and _67826_ (_16276_, _16275_, _16274_);
  or _67827_ (_16277_, _16276_, _03216_);
  and _67828_ (_16278_, _16277_, _16129_);
  or _67829_ (_16279_, _16278_, _03601_);
  and _67830_ (_16280_, _06298_, _05254_);
  nor _67831_ (_16281_, _16280_, _16122_);
  nand _67832_ (_16283_, _16281_, _03601_);
  and _67833_ (_16284_, _16283_, _08364_);
  and _67834_ (_16285_, _16284_, _16279_);
  or _67835_ (_16286_, _16285_, _16127_);
  and _67836_ (_16287_, _16286_, _08377_);
  and _67837_ (_16288_, _08371_, _08669_);
  or _67838_ (_16289_, _16288_, _08380_);
  or _67839_ (_16290_, _16289_, _16287_);
  not _67840_ (_16291_, _08381_);
  and _67841_ (_16292_, _08669_, _16291_);
  or _67842_ (_16294_, _16292_, _08382_);
  and _67843_ (_16295_, _16294_, _16290_);
  or _67844_ (_16296_, _16295_, _16126_);
  and _67845_ (_16297_, _16296_, _08387_);
  nor _67846_ (_16298_, _08387_, _08670_);
  or _67847_ (_16299_, _16298_, _15649_);
  or _67848_ (_16300_, _16299_, _16297_);
  or _67849_ (_16301_, _15650_, _08634_);
  and _67850_ (_16302_, _16301_, _15476_);
  and _67851_ (_16303_, _16302_, _16300_);
  and _67852_ (_16305_, _08634_, _04182_);
  or _67853_ (_16306_, _16305_, _03778_);
  or _67854_ (_16307_, _16306_, _16303_);
  or _67855_ (_16308_, _12817_, _03779_);
  and _67856_ (_16309_, _16308_, _07905_);
  and _67857_ (_16310_, _16309_, _16307_);
  and _67858_ (_16311_, _08743_, _07904_);
  or _67859_ (_16312_, _16311_, _03600_);
  or _67860_ (_16313_, _16312_, _16310_);
  and _67861_ (_16314_, _16313_, _16125_);
  or _67862_ (_16316_, _16314_, _03780_);
  or _67863_ (_16317_, _16122_, _07778_);
  and _67864_ (_16318_, _16317_, _08417_);
  and _67865_ (_16319_, _16318_, _16316_);
  and _67866_ (_16320_, _08421_, _08667_);
  or _67867_ (_16321_, _16320_, _08420_);
  or _67868_ (_16322_, _16321_, _16319_);
  or _67869_ (_16323_, _08425_, _08632_);
  and _67870_ (_16324_, _16323_, _03789_);
  and _67871_ (_16325_, _16324_, _16322_);
  or _67872_ (_16327_, _12815_, _08429_);
  and _67873_ (_16328_, _16327_, _08431_);
  or _67874_ (_16329_, _16328_, _16325_);
  or _67875_ (_16330_, _08435_, _08741_);
  and _67876_ (_16331_, _16330_, _07777_);
  and _67877_ (_16332_, _16331_, _16329_);
  or _67878_ (_16333_, _16281_, _12816_);
  nor _67879_ (_16334_, _16333_, _07777_);
  or _67880_ (_16335_, _16334_, _08446_);
  or _67881_ (_16336_, _16335_, _16332_);
  nand _67882_ (_16338_, _08446_, _08668_);
  and _67883_ (_16339_, _16338_, _16336_);
  or _67884_ (_16340_, _16339_, _08450_);
  nand _67885_ (_16341_, _08450_, _08633_);
  and _67886_ (_16342_, _16341_, _03784_);
  and _67887_ (_16343_, _16342_, _16340_);
  nor _67888_ (_16344_, _12816_, _03784_);
  or _67889_ (_16345_, _16344_, _08458_);
  or _67890_ (_16346_, _16345_, _16343_);
  nand _67891_ (_16347_, _08458_, _08742_);
  and _67892_ (_16349_, _16347_, _16346_);
  or _67893_ (_16350_, _16349_, _03624_);
  nor _67894_ (_16351_, _12819_, _07908_);
  nor _67895_ (_16352_, _16351_, _16122_);
  nand _67896_ (_16353_, _16352_, _03624_);
  and _67897_ (_16354_, _16353_, _07898_);
  and _67898_ (_16355_, _16354_, _16350_);
  and _67899_ (_16356_, _07881_, _07847_);
  nor _67900_ (_16357_, _16356_, _07882_);
  and _67901_ (_16358_, _16357_, _08468_);
  or _67902_ (_16360_, _16358_, _08475_);
  or _67903_ (_16361_, _16360_, _16355_);
  and _67904_ (_16362_, _08493_, _08014_);
  nor _67905_ (_16363_, _16362_, _08494_);
  or _67906_ (_16364_, _16363_, _08477_);
  and _67907_ (_16365_, _16364_, _16361_);
  or _67908_ (_16366_, _16365_, _03776_);
  and _67909_ (_16367_, _08574_, _08546_);
  nor _67910_ (_16368_, _16367_, _08575_);
  or _67911_ (_16369_, _16368_, _03777_);
  and _67912_ (_16371_, _16369_, _08589_);
  and _67913_ (_16372_, _16371_, _16366_);
  and _67914_ (_16373_, _08604_, _07941_);
  nor _67915_ (_16374_, _16373_, _08605_);
  and _67916_ (_16375_, _16374_, _08506_);
  or _67917_ (_16376_, _16375_, _08587_);
  or _67918_ (_16377_, _16376_, _16372_);
  nand _67919_ (_16378_, _08587_, _07578_);
  and _67920_ (_16379_, _16378_, _08617_);
  and _67921_ (_16380_, _16379_, _16377_);
  and _67922_ (_16382_, _08687_, _08670_);
  nor _67923_ (_16383_, _16382_, _08688_);
  and _67924_ (_16384_, _16383_, _08618_);
  or _67925_ (_16385_, _16384_, _16380_);
  and _67926_ (_16386_, _16385_, _08624_);
  nor _67927_ (_16387_, _08651_, _08634_);
  nor _67928_ (_16388_, _16387_, _08652_);
  and _67929_ (_16389_, _16388_, _08620_);
  or _67930_ (_16390_, _16389_, _03517_);
  or _67931_ (_16391_, _16390_, _16386_);
  nor _67932_ (_16393_, _08719_, _08707_);
  nor _67933_ (_16394_, _16393_, _08720_);
  or _67934_ (_16395_, _16394_, _03518_);
  and _67935_ (_16396_, _16395_, _08734_);
  and _67936_ (_16397_, _16396_, _16391_);
  nor _67937_ (_16398_, _08759_, _08743_);
  nor _67938_ (_16399_, _16398_, _08760_);
  and _67939_ (_16400_, _16399_, _08701_);
  or _67940_ (_16401_, _16400_, _08732_);
  or _67941_ (_16402_, _16401_, _16397_);
  and _67942_ (_16404_, _16402_, _16121_);
  or _67943_ (_16405_, _16404_, _03815_);
  nand _67944_ (_16406_, _16167_, _03815_);
  and _67945_ (_16407_, _16406_, _08776_);
  and _67946_ (_16408_, _16407_, _16405_);
  and _67947_ (_16409_, _08782_, _07484_);
  nor _67948_ (_16410_, _08782_, _07484_);
  nor _67949_ (_16411_, _16410_, _16409_);
  not _67950_ (_16412_, _16411_);
  and _67951_ (_16413_, _16412_, _08775_);
  or _67952_ (_16415_, _16413_, _08780_);
  or _67953_ (_16416_, _16415_, _16408_);
  nand _67954_ (_16417_, _08780_, _07478_);
  and _67955_ (_16418_, _16417_, _03823_);
  and _67956_ (_16419_, _16418_, _16416_);
  nor _67957_ (_16420_, _16199_, _03823_);
  or _67958_ (_16421_, _16420_, _03447_);
  or _67959_ (_16422_, _16421_, _16419_);
  and _67960_ (_16423_, _13003_, _05254_);
  nor _67961_ (_16424_, _16423_, _16122_);
  nand _67962_ (_16426_, _16424_, _03447_);
  and _67963_ (_16427_, _16426_, _08799_);
  and _67964_ (_16428_, _16427_, _16422_);
  and _67965_ (_16429_, _08807_, _07484_);
  nor _67966_ (_16430_, _16429_, _08808_);
  and _67967_ (_16431_, _16430_, _08798_);
  or _67968_ (_16432_, _16431_, _08805_);
  or _67969_ (_16433_, _16432_, _16428_);
  nand _67970_ (_16434_, _08805_, _07478_);
  and _67971_ (_16435_, _16434_, _43000_);
  and _67972_ (_16437_, _16435_, _16433_);
  or _67973_ (_16438_, _16437_, _16120_);
  and _67974_ (_43495_, _16438_, _41806_);
  nor _67975_ (_16439_, _43000_, _07478_);
  nor _67976_ (_16440_, _05254_, _07478_);
  nor _67977_ (_16441_, _13140_, _07908_);
  nor _67978_ (_16442_, _16441_, _16440_);
  nor _67979_ (_16443_, _16442_, _07795_);
  and _67980_ (_16444_, _06306_, _05254_);
  nor _67981_ (_16445_, _16444_, _16440_);
  or _67982_ (_16447_, _16445_, _13146_);
  nor _67983_ (_16448_, _16447_, _07777_);
  and _67984_ (_16449_, _13141_, _05254_);
  nor _67985_ (_16450_, _16449_, _16440_);
  nand _67986_ (_16451_, _16450_, _03600_);
  or _67987_ (_16452_, _08630_, _15476_);
  nor _67988_ (_16453_, _08665_, _08666_);
  nor _67989_ (_16454_, _15641_, _04181_);
  and _67990_ (_16455_, _16454_, _08382_);
  and _67991_ (_16456_, _16455_, _08377_);
  or _67992_ (_16458_, _16456_, _16453_);
  nand _67993_ (_16459_, _03860_, _03216_);
  nor _67994_ (_16460_, _05469_, _07908_);
  nor _67995_ (_16461_, _16460_, _16440_);
  nand _67996_ (_16462_, _16461_, _07390_);
  and _67997_ (_16463_, _03486_, \oc8051_golden_model_1.ACC [4]);
  nor _67998_ (_16464_, _16240_, _16463_);
  nor _67999_ (_16465_, _10026_, _16464_);
  and _68000_ (_16466_, _10026_, _16464_);
  nor _68001_ (_16467_, _16466_, _16465_);
  and _68002_ (_16469_, _16467_, \oc8051_golden_model_1.PSW [7]);
  nor _68003_ (_16470_, _16467_, \oc8051_golden_model_1.PSW [7]);
  nor _68004_ (_16471_, _16470_, _16469_);
  nor _68005_ (_16472_, _16246_, _16243_);
  not _68006_ (_16473_, _16472_);
  and _68007_ (_16474_, _16473_, _16471_);
  nor _68008_ (_16475_, _16473_, _16471_);
  nor _68009_ (_16476_, _16475_, _16474_);
  or _68010_ (_16477_, _16476_, _07914_);
  nor _68011_ (_16478_, _05903_, _07478_);
  and _68012_ (_16480_, _13037_, _05903_);
  and _68013_ (_16481_, _16480_, _13054_);
  nor _68014_ (_16482_, _16481_, _16478_);
  nor _68015_ (_16483_, _16482_, _06840_);
  nand _68016_ (_16484_, _08064_, _05469_);
  or _68017_ (_16485_, _08067_, _06684_);
  nor _68018_ (_16486_, _08078_, _05469_);
  and _68019_ (_16487_, _04064_, _07478_);
  nor _68020_ (_16488_, _04064_, _07478_);
  or _68021_ (_16489_, _16488_, _16487_);
  and _68022_ (_16491_, _16489_, _08078_);
  or _68023_ (_16492_, _16491_, _08066_);
  or _68024_ (_16493_, _16492_, _16486_);
  and _68025_ (_16494_, _16493_, _08069_);
  and _68026_ (_16495_, _16494_, _16485_);
  nor _68027_ (_16496_, _13014_, _07908_);
  nor _68028_ (_16497_, _16496_, _16440_);
  nor _68029_ (_16498_, _16497_, _04081_);
  or _68030_ (_16499_, _16498_, _08089_);
  or _68031_ (_16500_, _16499_, _16495_);
  and _68032_ (_16502_, _09893_, _08104_);
  nor _68033_ (_16503_, _09893_, _08104_);
  nor _68034_ (_16504_, _16503_, _16502_);
  nand _68035_ (_16505_, _16504_, _08089_);
  and _68036_ (_16506_, _16505_, _16500_);
  or _68037_ (_16507_, _16506_, _03715_);
  nor _68038_ (_16508_, _16480_, _16478_);
  nand _68039_ (_16509_, _16508_, _03715_);
  and _68040_ (_16510_, _16509_, _03996_);
  and _68041_ (_16511_, _16510_, _16507_);
  nor _68042_ (_16513_, _16461_, _03996_);
  or _68043_ (_16514_, _16513_, _08064_);
  or _68044_ (_16515_, _16514_, _16511_);
  and _68045_ (_16516_, _16515_, _16484_);
  or _68046_ (_16517_, _16516_, _04443_);
  or _68047_ (_16518_, _06684_, _08128_);
  and _68048_ (_16519_, _16518_, _03737_);
  and _68049_ (_16520_, _16519_, _16517_);
  nor _68050_ (_16521_, _08218_, _03737_);
  or _68051_ (_16522_, _16521_, _08132_);
  or _68052_ (_16524_, _16522_, _16520_);
  nand _68053_ (_16525_, _08132_, _03274_);
  and _68054_ (_16526_, _16525_, _16524_);
  or _68055_ (_16527_, _16526_, _03714_);
  and _68056_ (_16528_, _13047_, _05903_);
  nor _68057_ (_16529_, _16528_, _16478_);
  nand _68058_ (_16530_, _16529_, _03714_);
  and _68059_ (_16531_, _16530_, _06840_);
  and _68060_ (_16532_, _16531_, _16527_);
  or _68061_ (_16533_, _16532_, _16483_);
  and _68062_ (_16535_, _16533_, _06875_);
  nor _68063_ (_16536_, _07342_, _07340_);
  nor _68064_ (_16537_, _16536_, _07343_);
  and _68065_ (_16538_, _16537_, _06869_);
  or _68066_ (_16539_, _16538_, _10170_);
  or _68067_ (_16540_, _16539_, _16535_);
  and _68068_ (_16541_, _05777_, \oc8051_golden_model_1.ACC [4]);
  nor _68069_ (_16542_, _16220_, _16541_);
  nor _68070_ (_16543_, _16453_, _16542_);
  and _68071_ (_16544_, _16453_, _16542_);
  nor _68072_ (_16546_, _16544_, _16543_);
  and _68073_ (_16547_, _16546_, \oc8051_golden_model_1.PSW [7]);
  nor _68074_ (_16548_, _16546_, \oc8051_golden_model_1.PSW [7]);
  nor _68075_ (_16549_, _16548_, _16547_);
  nor _68076_ (_16550_, _16226_, _16223_);
  not _68077_ (_16551_, _16550_);
  and _68078_ (_16552_, _16551_, _16549_);
  nor _68079_ (_16553_, _16551_, _16549_);
  nor _68080_ (_16554_, _16553_, _16552_);
  or _68081_ (_16555_, _16554_, _08058_);
  and _68082_ (_16558_, _16555_, _08054_);
  and _68083_ (_16559_, _16558_, _16540_);
  and _68084_ (_16560_, _16554_, _08053_);
  or _68085_ (_16561_, _16560_, _08051_);
  or _68086_ (_16562_, _16561_, _16559_);
  nor _68087_ (_16563_, _06730_, _07484_);
  nor _68088_ (_16564_, _16143_, _16563_);
  nor _68089_ (_16565_, _08630_, _16564_);
  and _68090_ (_16566_, _08630_, _16564_);
  nor _68091_ (_16567_, _16566_, _16565_);
  and _68092_ (_16569_, _16567_, \oc8051_golden_model_1.PSW [7]);
  nor _68093_ (_16570_, _16567_, \oc8051_golden_model_1.PSW [7]);
  nor _68094_ (_16571_, _16570_, _16569_);
  nor _68095_ (_16572_, _16149_, _16146_);
  not _68096_ (_16573_, _16572_);
  and _68097_ (_16574_, _16573_, _16571_);
  nor _68098_ (_16575_, _16573_, _16571_);
  nor _68099_ (_16576_, _16575_, _16574_);
  or _68100_ (_16577_, _16576_, _10201_);
  and _68101_ (_16578_, _16577_, _03766_);
  and _68102_ (_16580_, _16578_, _16562_);
  and _68103_ (_16581_, _08324_, _08311_);
  nor _68104_ (_16582_, _16581_, _08325_);
  nor _68105_ (_16583_, _16582_, _03766_);
  or _68106_ (_16584_, _16583_, _07913_);
  or _68107_ (_16585_, _16584_, _16580_);
  and _68108_ (_16586_, _16585_, _16477_);
  or _68109_ (_16587_, _16586_, _07912_);
  nand _68110_ (_16588_, _03860_, _07912_);
  and _68111_ (_16589_, _16588_, _03710_);
  and _68112_ (_16591_, _16589_, _16587_);
  nor _68113_ (_16592_, _13020_, _08339_);
  nor _68114_ (_16593_, _16592_, _16478_);
  nor _68115_ (_16594_, _16593_, _03710_);
  or _68116_ (_16595_, _16594_, _07390_);
  or _68117_ (_16596_, _16595_, _16591_);
  and _68118_ (_16597_, _16596_, _16462_);
  or _68119_ (_16598_, _16597_, _04481_);
  and _68120_ (_16599_, _06684_, _05254_);
  nor _68121_ (_16600_, _16599_, _16440_);
  nand _68122_ (_16602_, _16600_, _04481_);
  and _68123_ (_16603_, _16602_, _03589_);
  and _68124_ (_16604_, _16603_, _16598_);
  nor _68125_ (_16605_, _13127_, _07908_);
  nor _68126_ (_16606_, _16605_, _16440_);
  nor _68127_ (_16607_, _16606_, _03589_);
  or _68128_ (_16608_, _16607_, _07405_);
  or _68129_ (_16609_, _16608_, _16604_);
  or _68130_ (_16610_, _07463_, _07411_);
  and _68131_ (_16611_, _16610_, _16609_);
  or _68132_ (_16613_, _16611_, _03216_);
  and _68133_ (_16614_, _16613_, _16459_);
  or _68134_ (_16615_, _16614_, _03601_);
  nand _68135_ (_16616_, _16445_, _03601_);
  and _68136_ (_16617_, _16616_, _08364_);
  and _68137_ (_16618_, _16617_, _16615_);
  or _68138_ (_16619_, _08364_, _03860_);
  nand _68139_ (_16620_, _16619_, _16456_);
  or _68140_ (_16621_, _16620_, _16618_);
  and _68141_ (_16622_, _16621_, _16458_);
  or _68142_ (_16624_, _16622_, _15478_);
  or _68143_ (_16625_, _16453_, _15651_);
  and _68144_ (_16626_, _16625_, _15650_);
  and _68145_ (_16627_, _16626_, _16624_);
  or _68146_ (_16628_, _08630_, _04182_);
  and _68147_ (_16629_, _16628_, _08392_);
  or _68148_ (_16630_, _16629_, _16627_);
  and _68149_ (_16631_, _16630_, _16452_);
  or _68150_ (_16632_, _16631_, _03778_);
  or _68151_ (_16633_, _13147_, _03779_);
  and _68152_ (_16635_, _16633_, _07905_);
  and _68153_ (_16636_, _16635_, _16632_);
  and _68154_ (_16637_, _10026_, _07904_);
  or _68155_ (_16638_, _16637_, _03600_);
  or _68156_ (_16639_, _16638_, _16636_);
  and _68157_ (_16640_, _16639_, _16451_);
  or _68158_ (_16641_, _16640_, _03780_);
  or _68159_ (_16642_, _16440_, _07778_);
  and _68160_ (_16643_, _16642_, _08417_);
  and _68161_ (_16644_, _16643_, _16641_);
  and _68162_ (_16646_, _08421_, _08665_);
  or _68163_ (_16647_, _16646_, _08420_);
  or _68164_ (_16648_, _16647_, _16644_);
  or _68165_ (_16649_, _08425_, _08628_);
  and _68166_ (_16650_, _16649_, _03789_);
  and _68167_ (_16651_, _16650_, _16648_);
  or _68168_ (_16652_, _13145_, _08429_);
  and _68169_ (_16653_, _16652_, _08431_);
  or _68170_ (_16654_, _16653_, _16651_);
  or _68171_ (_16655_, _08435_, _08739_);
  and _68172_ (_16657_, _16655_, _07777_);
  and _68173_ (_16658_, _16657_, _16654_);
  or _68174_ (_16659_, _16658_, _16448_);
  and _68175_ (_16660_, _16659_, _15121_);
  nor _68176_ (_16661_, _15121_, _08666_);
  or _68177_ (_16662_, _16661_, _15123_);
  or _68178_ (_16663_, _16662_, _16660_);
  nand _68179_ (_16664_, _15123_, _08666_);
  and _68180_ (_16665_, _16664_, _15128_);
  and _68181_ (_16666_, _16665_, _16663_);
  nor _68182_ (_16668_, _08666_, _15128_);
  or _68183_ (_16669_, _16668_, _08450_);
  or _68184_ (_16670_, _16669_, _16666_);
  nand _68185_ (_16671_, _08450_, _08629_);
  and _68186_ (_16672_, _16671_, _03784_);
  and _68187_ (_16673_, _16672_, _16670_);
  nor _68188_ (_16674_, _13146_, _03784_);
  or _68189_ (_16675_, _16674_, _08458_);
  or _68190_ (_16676_, _16675_, _16673_);
  nand _68191_ (_16677_, _08458_, _08740_);
  and _68192_ (_16679_, _16677_, _07795_);
  and _68193_ (_16680_, _16679_, _16676_);
  or _68194_ (_16681_, _16680_, _16443_);
  and _68195_ (_16682_, _16681_, _07898_);
  and _68196_ (_16683_, _07883_, _07841_);
  nor _68197_ (_16684_, _16683_, _07884_);
  and _68198_ (_16685_, _16684_, _08468_);
  or _68199_ (_16686_, _16685_, _08475_);
  or _68200_ (_16687_, _16686_, _16682_);
  and _68201_ (_16688_, _08495_, _08012_);
  nor _68202_ (_16690_, _16688_, _08496_);
  or _68203_ (_16691_, _16690_, _08477_);
  and _68204_ (_16692_, _16691_, _03777_);
  and _68205_ (_16693_, _16692_, _16687_);
  and _68206_ (_16694_, _08576_, _08540_);
  nor _68207_ (_16695_, _16694_, _08577_);
  or _68208_ (_16696_, _16695_, _08506_);
  and _68209_ (_16697_, _16696_, _08508_);
  or _68210_ (_16698_, _16697_, _16693_);
  and _68211_ (_16699_, _08606_, _07939_);
  nor _68212_ (_16701_, _16699_, _08607_);
  or _68213_ (_16702_, _16701_, _08589_);
  and _68214_ (_16703_, _16702_, _08588_);
  and _68215_ (_16704_, _16703_, _16698_);
  not _68216_ (_16705_, _04226_);
  and _68217_ (_16706_, _10320_, _16705_);
  nand _68218_ (_16707_, _08587_, \oc8051_golden_model_1.ACC [4]);
  nand _68219_ (_16708_, _16707_, _16706_);
  or _68220_ (_16709_, _16708_, _16704_);
  and _68221_ (_16710_, _03494_, _03202_);
  not _68222_ (_16712_, _16710_);
  nor _68223_ (_16713_, _08689_, _16453_);
  and _68224_ (_16714_, _08689_, _16453_);
  or _68225_ (_16715_, _16714_, _16713_);
  or _68226_ (_16716_, _16715_, _16706_);
  and _68227_ (_16717_, _16716_, _16712_);
  and _68228_ (_16718_, _16717_, _16709_);
  and _68229_ (_16719_, _16715_, _16710_);
  or _68230_ (_16720_, _16719_, _08620_);
  or _68231_ (_16721_, _16720_, _16718_);
  and _68232_ (_16723_, _08653_, _08631_);
  nor _68233_ (_16724_, _16723_, _08654_);
  or _68234_ (_16725_, _16724_, _08624_);
  and _68235_ (_16726_, _16725_, _03518_);
  and _68236_ (_16727_, _16726_, _16721_);
  and _68237_ (_16728_, _08721_, _08308_);
  nor _68238_ (_16729_, _16728_, _08722_);
  or _68239_ (_16730_, _16729_, _08701_);
  and _68240_ (_16731_, _16730_, _08703_);
  or _68241_ (_16732_, _16731_, _16727_);
  not _68242_ (_16734_, _10026_);
  nor _68243_ (_16735_, _08761_, _16734_);
  and _68244_ (_16736_, _08761_, _16734_);
  nor _68245_ (_16737_, _16736_, _16735_);
  or _68246_ (_16738_, _16737_, _08734_);
  and _68247_ (_16739_, _16738_, _08733_);
  and _68248_ (_16740_, _16739_, _16732_);
  and _68249_ (_16741_, _08732_, \oc8051_golden_model_1.ACC [4]);
  or _68250_ (_16742_, _16741_, _03815_);
  or _68251_ (_16743_, _16742_, _16740_);
  nand _68252_ (_16745_, _16497_, _03815_);
  and _68253_ (_16746_, _16745_, _08776_);
  and _68254_ (_16747_, _16746_, _16743_);
  nor _68255_ (_16748_, _16409_, _07478_);
  or _68256_ (_16749_, _16748_, _08783_);
  and _68257_ (_16750_, _16749_, _08775_);
  or _68258_ (_16751_, _16750_, _08780_);
  or _68259_ (_16752_, _16751_, _16747_);
  nand _68260_ (_16753_, _08780_, _07433_);
  and _68261_ (_16754_, _16753_, _03823_);
  and _68262_ (_16756_, _16754_, _16752_);
  nor _68263_ (_16757_, _16529_, _03823_);
  or _68264_ (_16758_, _16757_, _03447_);
  or _68265_ (_16759_, _16758_, _16756_);
  and _68266_ (_16760_, _13199_, _05254_);
  nor _68267_ (_16761_, _16760_, _16440_);
  nand _68268_ (_16762_, _16761_, _03447_);
  and _68269_ (_16763_, _16762_, _08799_);
  and _68270_ (_16764_, _16763_, _16759_);
  nor _68271_ (_16765_, _08808_, \oc8051_golden_model_1.ACC [5]);
  nor _68272_ (_16767_, _16765_, _08809_);
  nor _68273_ (_16768_, _16767_, _08805_);
  nor _68274_ (_16769_, _16768_, _11964_);
  or _68275_ (_16770_, _16769_, _16764_);
  nand _68276_ (_16771_, _08805_, _07433_);
  and _68277_ (_16772_, _16771_, _43000_);
  and _68278_ (_16773_, _16772_, _16770_);
  or _68279_ (_16774_, _16773_, _16439_);
  and _68280_ (_43496_, _16774_, _41806_);
  nor _68281_ (_16775_, _43000_, _07433_);
  nand _68282_ (_16777_, _08732_, _07478_);
  nor _68283_ (_16778_, _05254_, _07433_);
  and _68284_ (_16779_, _13339_, _05254_);
  nor _68285_ (_16780_, _16779_, _16778_);
  or _68286_ (_16781_, _16780_, _13352_);
  nor _68287_ (_16782_, _16781_, _07777_);
  and _68288_ (_16783_, _13347_, _05254_);
  nor _68289_ (_16784_, _16783_, _16778_);
  nand _68290_ (_16785_, _16784_, _03600_);
  and _68291_ (_16786_, _08387_, _16291_);
  not _68292_ (_16788_, _16786_);
  and _68293_ (_16789_, _16788_, _08664_);
  or _68294_ (_16790_, _08377_, _08664_);
  nand _68295_ (_16791_, _03549_, _03216_);
  nor _68296_ (_16792_, _05363_, _07908_);
  nor _68297_ (_16793_, _16792_, _16778_);
  nand _68298_ (_16794_, _16793_, _07390_);
  and _68299_ (_16795_, _08326_, _08307_);
  nor _68300_ (_16796_, _16795_, _08327_);
  nand _68301_ (_16797_, _16796_, _03761_);
  and _68302_ (_16799_, _16797_, _07914_);
  or _68303_ (_16800_, _06684_, _07478_);
  and _68304_ (_16801_, _06684_, _07478_);
  or _68305_ (_16802_, _16564_, _16801_);
  and _68306_ (_16803_, _16802_, _16800_);
  nor _68307_ (_16804_, _16803_, _08627_);
  and _68308_ (_16805_, _16803_, _08627_);
  nor _68309_ (_16806_, _16805_, _16804_);
  nor _68310_ (_16807_, _16574_, _16569_);
  and _68311_ (_16808_, _16807_, \oc8051_golden_model_1.PSW [7]);
  nor _68312_ (_16810_, _16808_, _16806_);
  and _68313_ (_16811_, _16808_, _16806_);
  nor _68314_ (_16812_, _16811_, _16810_);
  and _68315_ (_16813_, _16812_, _08051_);
  nand _68316_ (_16814_, _08064_, _05363_);
  nor _68317_ (_16815_, _13242_, _07908_);
  nor _68318_ (_16816_, _16815_, _16778_);
  nor _68319_ (_16817_, _16816_, _04081_);
  or _68320_ (_16818_, _08067_, _06455_);
  nor _68321_ (_16819_, _08078_, _05363_);
  and _68322_ (_16821_, _04064_, _07433_);
  nor _68323_ (_16822_, _04064_, _07433_);
  or _68324_ (_16823_, _16822_, _16821_);
  and _68325_ (_16824_, _16823_, _08078_);
  or _68326_ (_16825_, _16824_, _08066_);
  or _68327_ (_16826_, _16825_, _16819_);
  and _68328_ (_16827_, _16826_, _08069_);
  and _68329_ (_16828_, _16827_, _16818_);
  or _68330_ (_16829_, _16828_, _16817_);
  and _68331_ (_16830_, _16829_, _09882_);
  not _68332_ (_16832_, _08106_);
  nor _68333_ (_16833_, _16503_, _16832_);
  and _68334_ (_16834_, _09892_, _08107_);
  nor _68335_ (_16835_, _16834_, _16833_);
  nor _68336_ (_16836_, _16835_, _09882_);
  or _68337_ (_16837_, _16836_, _03715_);
  or _68338_ (_16838_, _16837_, _16830_);
  nor _68339_ (_16839_, _05903_, _07433_);
  and _68340_ (_16840_, _13229_, _05903_);
  nor _68341_ (_16841_, _16840_, _16839_);
  nand _68342_ (_16843_, _16841_, _03715_);
  and _68343_ (_16844_, _16843_, _03996_);
  and _68344_ (_16845_, _16844_, _16838_);
  nor _68345_ (_16846_, _16793_, _03996_);
  or _68346_ (_16847_, _16846_, _08064_);
  or _68347_ (_16848_, _16847_, _16845_);
  and _68348_ (_16849_, _16848_, _16814_);
  or _68349_ (_16850_, _16849_, _04443_);
  or _68350_ (_16851_, _06455_, _08128_);
  and _68351_ (_16852_, _16851_, _03737_);
  and _68352_ (_16854_, _16852_, _16850_);
  nor _68353_ (_16855_, _08203_, _03737_);
  or _68354_ (_16856_, _16855_, _08132_);
  or _68355_ (_16857_, _16856_, _16854_);
  nand _68356_ (_16858_, _08132_, _07584_);
  and _68357_ (_16859_, _16858_, _16857_);
  or _68358_ (_16860_, _16859_, _03714_);
  and _68359_ (_16861_, _13253_, _05903_);
  nor _68360_ (_16862_, _16861_, _16839_);
  nand _68361_ (_16863_, _16862_, _03714_);
  and _68362_ (_16865_, _16863_, _06840_);
  and _68363_ (_16866_, _16865_, _16860_);
  and _68364_ (_16867_, _16840_, _13260_);
  nor _68365_ (_16868_, _16867_, _16839_);
  nor _68366_ (_16869_, _16868_, _06840_);
  or _68367_ (_16870_, _16869_, _06869_);
  or _68368_ (_16871_, _16870_, _16866_);
  nor _68369_ (_16872_, _07345_, _07343_);
  nor _68370_ (_16873_, _16872_, _07346_);
  or _68371_ (_16874_, _16873_, _06875_);
  and _68372_ (_16876_, _16874_, _16871_);
  or _68373_ (_16877_, _16876_, _08060_);
  nand _68374_ (_16878_, _05469_, \oc8051_golden_model_1.ACC [5]);
  nor _68375_ (_16879_, _05469_, \oc8051_golden_model_1.ACC [5]);
  or _68376_ (_16880_, _16542_, _16879_);
  and _68377_ (_16881_, _16880_, _16878_);
  nor _68378_ (_16882_, _16881_, _08664_);
  and _68379_ (_16883_, _16881_, _08664_);
  nor _68380_ (_16884_, _16883_, _16882_);
  nor _68381_ (_16885_, _16552_, _16547_);
  and _68382_ (_16887_, _16885_, \oc8051_golden_model_1.PSW [7]);
  or _68383_ (_16888_, _16887_, _16884_);
  nand _68384_ (_16889_, _16887_, _16884_);
  and _68385_ (_16890_, _16889_, _16888_);
  and _68386_ (_16891_, _16890_, _10201_);
  or _68387_ (_16892_, _16891_, _11350_);
  and _68388_ (_16893_, _16892_, _16877_);
  or _68389_ (_16894_, _16893_, _03761_);
  or _68390_ (_16895_, _16894_, _16813_);
  and _68391_ (_16896_, _16895_, _16799_);
  or _68392_ (_16898_, _16464_, _10046_);
  and _68393_ (_16899_, _16898_, _10045_);
  nor _68394_ (_16900_, _16899_, _08738_);
  and _68395_ (_16901_, _16899_, _08738_);
  nor _68396_ (_16902_, _16901_, _16900_);
  nor _68397_ (_16903_, _16474_, _16469_);
  and _68398_ (_16904_, _16903_, \oc8051_golden_model_1.PSW [7]);
  or _68399_ (_16905_, _16904_, _16902_);
  nand _68400_ (_16906_, _16904_, _16902_);
  and _68401_ (_16907_, _16906_, _16905_);
  and _68402_ (_16909_, _16907_, _07913_);
  or _68403_ (_16910_, _16909_, _07912_);
  or _68404_ (_16911_, _16910_, _16896_);
  nand _68405_ (_16912_, _03549_, _07912_);
  and _68406_ (_16913_, _16912_, _03710_);
  and _68407_ (_16914_, _16913_, _16911_);
  nor _68408_ (_16915_, _13226_, _08339_);
  nor _68409_ (_16916_, _16915_, _16839_);
  nor _68410_ (_16917_, _16916_, _03710_);
  or _68411_ (_16918_, _16917_, _07390_);
  or _68412_ (_16920_, _16918_, _16914_);
  and _68413_ (_16921_, _16920_, _16794_);
  or _68414_ (_16922_, _16921_, _04481_);
  and _68415_ (_16923_, _06455_, _05254_);
  nor _68416_ (_16924_, _16923_, _16778_);
  nand _68417_ (_16925_, _16924_, _04481_);
  and _68418_ (_16926_, _16925_, _03589_);
  and _68419_ (_16927_, _16926_, _16922_);
  nor _68420_ (_16928_, _13332_, _07908_);
  nor _68421_ (_16929_, _16928_, _16778_);
  nor _68422_ (_16931_, _16929_, _03589_);
  or _68423_ (_16932_, _16931_, _07405_);
  or _68424_ (_16933_, _16932_, _16927_);
  not _68425_ (_16934_, _07434_);
  and _68426_ (_16935_, _07437_, _16934_);
  or _68427_ (_16936_, _16935_, _07411_);
  and _68428_ (_16937_, _16936_, _16933_);
  or _68429_ (_16938_, _16937_, _03216_);
  and _68430_ (_16939_, _16938_, _16791_);
  or _68431_ (_16940_, _16939_, _03601_);
  nand _68432_ (_16942_, _16780_, _03601_);
  and _68433_ (_16943_, _16942_, _08364_);
  and _68434_ (_16944_, _16943_, _16940_);
  nor _68435_ (_16945_, _08364_, _03549_);
  or _68436_ (_16946_, _16945_, _08371_);
  or _68437_ (_16947_, _16946_, _16944_);
  and _68438_ (_16948_, _16947_, _16790_);
  or _68439_ (_16949_, _16948_, _08380_);
  or _68440_ (_16950_, _08664_, _04180_);
  and _68441_ (_16951_, _16950_, _16786_);
  and _68442_ (_16953_, _16951_, _16949_);
  or _68443_ (_16954_, _16953_, _16789_);
  and _68444_ (_16955_, _16954_, _08393_);
  and _68445_ (_16956_, _08392_, _08627_);
  or _68446_ (_16957_, _16956_, _03778_);
  or _68447_ (_16958_, _16957_, _16955_);
  or _68448_ (_16959_, _13353_, _03779_);
  and _68449_ (_16960_, _16959_, _07905_);
  and _68450_ (_16961_, _16960_, _16958_);
  nor _68451_ (_16962_, _08737_, _07905_);
  or _68452_ (_16964_, _16962_, _03600_);
  or _68453_ (_16965_, _16964_, _16961_);
  nand _68454_ (_16966_, _16965_, _16785_);
  and _68455_ (_16967_, _16966_, _07778_);
  nor _68456_ (_16968_, _16778_, _07778_);
  or _68457_ (_16969_, _16968_, _15103_);
  nor _68458_ (_16970_, _16969_, _16967_);
  or _68459_ (_16971_, _08662_, _04199_);
  and _68460_ (_16972_, _16971_, _08421_);
  or _68461_ (_16973_, _16972_, _16970_);
  or _68462_ (_16975_, _08662_, _15367_);
  and _68463_ (_16976_, _16975_, _16973_);
  or _68464_ (_16977_, _16976_, _08420_);
  or _68465_ (_16978_, _08425_, _08625_);
  and _68466_ (_16979_, _16978_, _03789_);
  and _68467_ (_16980_, _16979_, _16977_);
  or _68468_ (_16981_, _13351_, _08429_);
  and _68469_ (_16982_, _16981_, _08431_);
  or _68470_ (_16983_, _16982_, _16980_);
  or _68471_ (_16984_, _08435_, _08735_);
  and _68472_ (_16986_, _16984_, _07777_);
  and _68473_ (_16987_, _16986_, _16983_);
  or _68474_ (_16988_, _16987_, _16782_);
  and _68475_ (_16989_, _16988_, _08447_);
  nor _68476_ (_16990_, _08447_, _08663_);
  or _68477_ (_16991_, _16990_, _08450_);
  or _68478_ (_16992_, _16991_, _16989_);
  nand _68479_ (_16993_, _08450_, _08626_);
  and _68480_ (_16994_, _16993_, _03784_);
  and _68481_ (_16995_, _16994_, _16992_);
  nor _68482_ (_16997_, _13352_, _03784_);
  or _68483_ (_16998_, _16997_, _08458_);
  or _68484_ (_16999_, _16998_, _16995_);
  nand _68485_ (_17000_, _08458_, _08736_);
  and _68486_ (_17001_, _17000_, _16999_);
  or _68487_ (_17002_, _17001_, _03624_);
  nor _68488_ (_17003_, _13346_, _07908_);
  nor _68489_ (_17004_, _17003_, _16778_);
  nand _68490_ (_17005_, _17004_, _03624_);
  and _68491_ (_17006_, _17005_, _07898_);
  and _68492_ (_17008_, _17006_, _17002_);
  and _68493_ (_17009_, _07885_, _07832_);
  nor _68494_ (_17010_, _17009_, _07886_);
  or _68495_ (_17011_, _17010_, _08475_);
  and _68496_ (_17012_, _17011_, _11885_);
  or _68497_ (_17013_, _17012_, _17008_);
  and _68498_ (_17014_, _08497_, _08479_);
  nor _68499_ (_17015_, _17014_, _08498_);
  or _68500_ (_17016_, _17015_, _08477_);
  and _68501_ (_17017_, _17016_, _17013_);
  or _68502_ (_17019_, _17017_, _03776_);
  and _68503_ (_17020_, _08578_, _08531_);
  nor _68504_ (_17021_, _17020_, _08579_);
  or _68505_ (_17022_, _17021_, _03777_);
  and _68506_ (_17023_, _17022_, _08589_);
  and _68507_ (_17024_, _17023_, _17019_);
  and _68508_ (_17025_, _08608_, _08591_);
  nor _68509_ (_17026_, _17025_, _08609_);
  and _68510_ (_17027_, _17026_, _08506_);
  or _68511_ (_17028_, _17027_, _08587_);
  or _68512_ (_17030_, _17028_, _17024_);
  nand _68513_ (_17031_, _08587_, _07478_);
  and _68514_ (_17032_, _17031_, _08617_);
  and _68515_ (_17033_, _17032_, _17030_);
  nor _68516_ (_17034_, _08691_, _08664_);
  nor _68517_ (_17035_, _17034_, _08692_);
  and _68518_ (_17036_, _17035_, _08618_);
  or _68519_ (_17037_, _17036_, _17033_);
  and _68520_ (_17038_, _17037_, _08624_);
  nor _68521_ (_17039_, _08655_, _08627_);
  nor _68522_ (_17041_, _17039_, _08656_);
  and _68523_ (_17042_, _17041_, _08620_);
  or _68524_ (_17043_, _17042_, _03517_);
  or _68525_ (_17044_, _17043_, _17038_);
  and _68526_ (_17045_, _08723_, _08206_);
  nor _68527_ (_17046_, _17045_, _08724_);
  or _68528_ (_17047_, _17046_, _03518_);
  and _68529_ (_17048_, _17047_, _08734_);
  and _68530_ (_17049_, _17048_, _17044_);
  nor _68531_ (_17050_, _08763_, _08738_);
  nor _68532_ (_17052_, _17050_, _08764_);
  and _68533_ (_17053_, _17052_, _08701_);
  or _68534_ (_17054_, _17053_, _08732_);
  or _68535_ (_17055_, _17054_, _17049_);
  and _68536_ (_17056_, _17055_, _16777_);
  or _68537_ (_17057_, _17056_, _03815_);
  nand _68538_ (_17058_, _16816_, _03815_);
  and _68539_ (_17059_, _17058_, _08776_);
  and _68540_ (_17060_, _17059_, _17057_);
  nor _68541_ (_17061_, _08783_, _07433_);
  or _68542_ (_17063_, _17061_, _08784_);
  and _68543_ (_17064_, _17063_, _08775_);
  or _68544_ (_17065_, _17064_, _08780_);
  or _68545_ (_17066_, _17065_, _17060_);
  nand _68546_ (_17067_, _08780_, _06075_);
  and _68547_ (_17068_, _17067_, _03823_);
  and _68548_ (_17069_, _17068_, _17066_);
  nor _68549_ (_17070_, _16862_, _03823_);
  or _68550_ (_17071_, _17070_, _03447_);
  or _68551_ (_17072_, _17071_, _17069_);
  and _68552_ (_17074_, _13402_, _05254_);
  nor _68553_ (_17075_, _17074_, _16778_);
  nand _68554_ (_17076_, _17075_, _03447_);
  and _68555_ (_17077_, _17076_, _08799_);
  and _68556_ (_17078_, _17077_, _17072_);
  nor _68557_ (_17079_, _08809_, \oc8051_golden_model_1.ACC [6]);
  nor _68558_ (_17080_, _17079_, _08810_);
  nor _68559_ (_17081_, _17080_, _08805_);
  nor _68560_ (_17082_, _17081_, _11964_);
  or _68561_ (_17083_, _17082_, _17078_);
  nand _68562_ (_17085_, _08805_, _06075_);
  and _68563_ (_17086_, _17085_, _43000_);
  and _68564_ (_17087_, _17086_, _17083_);
  or _68565_ (_17088_, _17087_, _16775_);
  and _68566_ (_43497_, _17088_, _41806_);
  not _68567_ (_17089_, \oc8051_golden_model_1.DPL [0]);
  nor _68568_ (_17090_, _43000_, _17089_);
  nor _68569_ (_17091_, _05303_, _17089_);
  and _68570_ (_17092_, _05303_, _04620_);
  or _68571_ (_17093_, _17092_, _17091_);
  or _68572_ (_17095_, _17093_, _06838_);
  and _68573_ (_17096_, _05303_, \oc8051_golden_model_1.ACC [0]);
  or _68574_ (_17097_, _17096_, _17091_);
  or _68575_ (_17098_, _17097_, _03737_);
  nor _68576_ (_17099_, _05666_, _08824_);
  or _68577_ (_17100_, _17099_, _17091_);
  or _68578_ (_17101_, _17100_, _04081_);
  and _68579_ (_17102_, _17097_, _04409_);
  nor _68580_ (_17103_, _04409_, _17089_);
  or _68581_ (_17104_, _17103_, _03610_);
  or _68582_ (_17106_, _17104_, _17102_);
  and _68583_ (_17107_, _17106_, _03996_);
  and _68584_ (_17108_, _17107_, _17101_);
  and _68585_ (_17109_, _17093_, _03723_);
  or _68586_ (_17110_, _17109_, _03729_);
  or _68587_ (_17111_, _17110_, _17108_);
  and _68588_ (_17112_, _17111_, _17098_);
  or _68589_ (_17113_, _17112_, _08847_);
  nand _68590_ (_17114_, _08847_, \oc8051_golden_model_1.DPL [0]);
  and _68591_ (_17115_, _17114_, _08832_);
  and _68592_ (_17117_, _17115_, _17113_);
  nor _68593_ (_17118_, _04163_, _08832_);
  or _68594_ (_17119_, _17118_, _07390_);
  or _68595_ (_17120_, _17119_, _17117_);
  and _68596_ (_17121_, _17120_, _17095_);
  or _68597_ (_17122_, _17121_, _04481_);
  and _68598_ (_17123_, _06546_, _05303_);
  or _68599_ (_17124_, _17091_, _07400_);
  or _68600_ (_17125_, _17124_, _17123_);
  and _68601_ (_17126_, _17125_, _17122_);
  or _68602_ (_17128_, _17126_, _03222_);
  nor _68603_ (_17129_, _12109_, _08824_);
  or _68604_ (_17130_, _17129_, _17091_);
  or _68605_ (_17131_, _17130_, _03589_);
  and _68606_ (_17132_, _17131_, _05886_);
  and _68607_ (_17133_, _17132_, _17128_);
  and _68608_ (_17134_, _05303_, _06274_);
  or _68609_ (_17135_, _17134_, _17091_);
  and _68610_ (_17136_, _17135_, _03601_);
  or _68611_ (_17137_, _17136_, _03600_);
  or _68612_ (_17139_, _17137_, _17133_);
  and _68613_ (_17140_, _12124_, _05303_);
  or _68614_ (_17141_, _17140_, _17091_);
  or _68615_ (_17142_, _17141_, _07766_);
  and _68616_ (_17143_, _17142_, _17139_);
  or _68617_ (_17144_, _17143_, _03780_);
  and _68618_ (_17145_, _12128_, _05303_);
  or _68619_ (_17146_, _17145_, _17091_);
  or _68620_ (_17147_, _17146_, _07778_);
  and _68621_ (_17148_, _17147_, _07777_);
  and _68622_ (_17150_, _17148_, _17144_);
  nand _68623_ (_17151_, _17135_, _03622_);
  nor _68624_ (_17152_, _17151_, _17099_);
  or _68625_ (_17153_, _17152_, _17150_);
  and _68626_ (_17154_, _17153_, _06828_);
  or _68627_ (_17155_, _17091_, _05666_);
  and _68628_ (_17156_, _17097_, _03790_);
  and _68629_ (_17157_, _17156_, _17155_);
  or _68630_ (_17158_, _17157_, _03624_);
  or _68631_ (_17159_, _17158_, _17154_);
  nor _68632_ (_17161_, _12122_, _08824_);
  or _68633_ (_17162_, _17091_, _07795_);
  or _68634_ (_17163_, _17162_, _17161_);
  and _68635_ (_17164_, _17163_, _07793_);
  and _68636_ (_17165_, _17164_, _17159_);
  not _68637_ (_17166_, _03909_);
  nor _68638_ (_17167_, _12003_, _08824_);
  or _68639_ (_17168_, _17167_, _17091_);
  and _68640_ (_17169_, _17168_, _03785_);
  or _68641_ (_17170_, _17169_, _17166_);
  or _68642_ (_17172_, _17170_, _17165_);
  or _68643_ (_17173_, _17100_, _03909_);
  and _68644_ (_17174_, _17173_, _43000_);
  and _68645_ (_17175_, _17174_, _17172_);
  or _68646_ (_17176_, _17175_, _17090_);
  and _68647_ (_43498_, _17176_, _41806_);
  not _68648_ (_17177_, \oc8051_golden_model_1.DPL [1]);
  nor _68649_ (_17178_, _43000_, _17177_);
  nor _68650_ (_17179_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor _68651_ (_17180_, _17179_, _08852_);
  and _68652_ (_17182_, _17180_, _08847_);
  or _68653_ (_17183_, _05303_, \oc8051_golden_model_1.DPL [1]);
  and _68654_ (_17184_, _12213_, _05303_);
  not _68655_ (_17185_, _17184_);
  and _68656_ (_17186_, _17185_, _17183_);
  or _68657_ (_17187_, _17186_, _04081_);
  nand _68658_ (_17188_, _05303_, _03274_);
  and _68659_ (_17189_, _17188_, _17183_);
  and _68660_ (_17190_, _17189_, _04409_);
  nor _68661_ (_17191_, _04409_, _17177_);
  or _68662_ (_17193_, _17191_, _03610_);
  or _68663_ (_17194_, _17193_, _17190_);
  and _68664_ (_17195_, _17194_, _03996_);
  and _68665_ (_17196_, _17195_, _17187_);
  nor _68666_ (_17197_, _05303_, _17177_);
  and _68667_ (_17198_, _05303_, _06764_);
  or _68668_ (_17199_, _17198_, _17197_);
  and _68669_ (_17200_, _17199_, _03723_);
  or _68670_ (_17201_, _17200_, _03729_);
  or _68671_ (_17202_, _17201_, _17196_);
  or _68672_ (_17204_, _17189_, _03737_);
  and _68673_ (_17205_, _17204_, _08848_);
  and _68674_ (_17206_, _17205_, _17202_);
  or _68675_ (_17207_, _17206_, _17182_);
  and _68676_ (_17208_, _17207_, _08832_);
  nor _68677_ (_17209_, _04303_, _08832_);
  or _68678_ (_17210_, _17209_, _07390_);
  or _68679_ (_17211_, _17210_, _17208_);
  or _68680_ (_17212_, _17199_, _06838_);
  and _68681_ (_17213_, _17212_, _17211_);
  or _68682_ (_17215_, _17213_, _04481_);
  and _68683_ (_17216_, _06501_, _05303_);
  or _68684_ (_17217_, _17197_, _07400_);
  or _68685_ (_17218_, _17217_, _17216_);
  and _68686_ (_17219_, _17218_, _03589_);
  and _68687_ (_17220_, _17219_, _17215_);
  nor _68688_ (_17221_, _12313_, _08824_);
  or _68689_ (_17222_, _17221_, _17197_);
  and _68690_ (_17223_, _17222_, _03222_);
  or _68691_ (_17224_, _17223_, _17220_);
  and _68692_ (_17226_, _17224_, _03602_);
  nand _68693_ (_17227_, _05303_, _04303_);
  and _68694_ (_17228_, _17183_, _03601_);
  and _68695_ (_17229_, _17228_, _17227_);
  or _68696_ (_17230_, _12327_, _08824_);
  and _68697_ (_17231_, _17183_, _03600_);
  and _68698_ (_17232_, _17231_, _17230_);
  or _68699_ (_17233_, _17232_, _17229_);
  or _68700_ (_17234_, _17233_, _17226_);
  and _68701_ (_17235_, _17234_, _07778_);
  or _68702_ (_17237_, _12333_, _08824_);
  and _68703_ (_17238_, _17183_, _03780_);
  and _68704_ (_17239_, _17238_, _17237_);
  or _68705_ (_17240_, _17239_, _17235_);
  and _68706_ (_17241_, _17240_, _07777_);
  or _68707_ (_17242_, _12207_, _08824_);
  and _68708_ (_17243_, _17183_, _03622_);
  and _68709_ (_17244_, _17243_, _17242_);
  or _68710_ (_17245_, _17244_, _17241_);
  and _68711_ (_17246_, _17245_, _06828_);
  or _68712_ (_17248_, _17197_, _05618_);
  and _68713_ (_17249_, _17189_, _03790_);
  and _68714_ (_17250_, _17249_, _17248_);
  or _68715_ (_17251_, _17250_, _17246_);
  and _68716_ (_17252_, _17251_, _03786_);
  or _68717_ (_17253_, _17227_, _05618_);
  and _68718_ (_17254_, _17183_, _03624_);
  and _68719_ (_17255_, _17254_, _17253_);
  or _68720_ (_17256_, _17188_, _05618_);
  and _68721_ (_17257_, _17183_, _03785_);
  and _68722_ (_17259_, _17257_, _17256_);
  or _68723_ (_17260_, _17259_, _03815_);
  or _68724_ (_17261_, _17260_, _17255_);
  or _68725_ (_17262_, _17261_, _17252_);
  or _68726_ (_17263_, _17186_, _04246_);
  and _68727_ (_17264_, _17263_, _17262_);
  or _68728_ (_17265_, _17264_, _03447_);
  or _68729_ (_17266_, _17197_, _03514_);
  or _68730_ (_17267_, _17266_, _17184_);
  and _68731_ (_17268_, _17267_, _43000_);
  and _68732_ (_17269_, _17268_, _17265_);
  or _68733_ (_17270_, _17269_, _17178_);
  and _68734_ (_43499_, _17270_, _41806_);
  not _68735_ (_17271_, \oc8051_golden_model_1.DPL [2]);
  nor _68736_ (_17272_, _43000_, _17271_);
  nor _68737_ (_17273_, _05303_, _17271_);
  nor _68738_ (_17274_, _12538_, _08824_);
  or _68739_ (_17275_, _17274_, _17273_);
  and _68740_ (_17276_, _17275_, _03785_);
  and _68741_ (_17277_, _12539_, _05303_);
  or _68742_ (_17280_, _17277_, _17273_);
  and _68743_ (_17281_, _17280_, _03780_);
  nor _68744_ (_17282_, _08824_, _04875_);
  or _68745_ (_17283_, _17282_, _17273_);
  or _68746_ (_17284_, _17283_, _03996_);
  nor _68747_ (_17285_, _12416_, _08824_);
  or _68748_ (_17286_, _17285_, _17273_);
  and _68749_ (_17287_, _17286_, _03610_);
  nor _68750_ (_17288_, _04409_, _17271_);
  and _68751_ (_17289_, _05303_, \oc8051_golden_model_1.ACC [2]);
  or _68752_ (_17290_, _17289_, _17273_);
  and _68753_ (_17291_, _17290_, _04409_);
  or _68754_ (_17292_, _17291_, _17288_);
  and _68755_ (_17293_, _17292_, _04081_);
  or _68756_ (_17294_, _17293_, _03723_);
  or _68757_ (_17295_, _17294_, _17287_);
  and _68758_ (_17296_, _17295_, _17284_);
  or _68759_ (_17297_, _17296_, _03729_);
  or _68760_ (_17298_, _17290_, _03737_);
  and _68761_ (_17299_, _17298_, _08848_);
  and _68762_ (_17302_, _17299_, _17297_);
  nor _68763_ (_17303_, _08852_, \oc8051_golden_model_1.DPL [2]);
  nor _68764_ (_17304_, _17303_, _08853_);
  and _68765_ (_17305_, _17304_, _08847_);
  or _68766_ (_17306_, _17305_, _17302_);
  and _68767_ (_17307_, _17306_, _08832_);
  nor _68768_ (_17308_, _03946_, _08832_);
  or _68769_ (_17309_, _17308_, _07390_);
  or _68770_ (_17310_, _17309_, _17307_);
  or _68771_ (_17311_, _17283_, _06838_);
  and _68772_ (_17313_, _17311_, _17310_);
  or _68773_ (_17314_, _17313_, _04481_);
  and _68774_ (_17315_, _06637_, _05303_);
  or _68775_ (_17316_, _17273_, _07400_);
  or _68776_ (_17317_, _17316_, _17315_);
  and _68777_ (_17318_, _17317_, _03589_);
  and _68778_ (_17319_, _17318_, _17314_);
  nor _68779_ (_17320_, _12519_, _08824_);
  or _68780_ (_17321_, _17320_, _17273_);
  and _68781_ (_17322_, _17321_, _03222_);
  or _68782_ (_17324_, _17322_, _08828_);
  or _68783_ (_17325_, _17324_, _17319_);
  and _68784_ (_17326_, _12533_, _05303_);
  or _68785_ (_17327_, _17273_, _07766_);
  or _68786_ (_17328_, _17327_, _17326_);
  and _68787_ (_17329_, _05303_, _06332_);
  or _68788_ (_17330_, _17329_, _17273_);
  or _68789_ (_17331_, _17330_, _05886_);
  and _68790_ (_17332_, _17331_, _07778_);
  and _68791_ (_17333_, _17332_, _17328_);
  and _68792_ (_17335_, _17333_, _17325_);
  or _68793_ (_17336_, _17335_, _17281_);
  and _68794_ (_17337_, _17336_, _07777_);
  or _68795_ (_17338_, _17273_, _05718_);
  and _68796_ (_17339_, _17330_, _03622_);
  and _68797_ (_17340_, _17339_, _17338_);
  or _68798_ (_17341_, _17340_, _17337_);
  and _68799_ (_17342_, _17341_, _06828_);
  and _68800_ (_17343_, _17290_, _03790_);
  and _68801_ (_17344_, _17343_, _17338_);
  or _68802_ (_17346_, _17344_, _03624_);
  or _68803_ (_17347_, _17346_, _17342_);
  nor _68804_ (_17348_, _12532_, _08824_);
  or _68805_ (_17349_, _17273_, _07795_);
  or _68806_ (_17350_, _17349_, _17348_);
  and _68807_ (_17351_, _17350_, _07793_);
  and _68808_ (_17352_, _17351_, _17347_);
  or _68809_ (_17353_, _17352_, _17276_);
  and _68810_ (_17354_, _17353_, _04246_);
  and _68811_ (_17355_, _17286_, _03815_);
  or _68812_ (_17357_, _17355_, _03447_);
  or _68813_ (_17358_, _17357_, _17354_);
  and _68814_ (_17359_, _12592_, _05303_);
  or _68815_ (_17360_, _17273_, _03514_);
  or _68816_ (_17361_, _17360_, _17359_);
  and _68817_ (_17362_, _17361_, _43000_);
  and _68818_ (_17363_, _17362_, _17358_);
  or _68819_ (_17364_, _17363_, _17272_);
  and _68820_ (_43500_, _17364_, _41806_);
  not _68821_ (_17365_, \oc8051_golden_model_1.DPL [3]);
  nor _68822_ (_17367_, _43000_, _17365_);
  nor _68823_ (_17368_, _05303_, _17365_);
  nor _68824_ (_17369_, _12738_, _08824_);
  or _68825_ (_17370_, _17369_, _17368_);
  and _68826_ (_17371_, _17370_, _03785_);
  and _68827_ (_17372_, _12739_, _05303_);
  or _68828_ (_17373_, _17372_, _17368_);
  and _68829_ (_17374_, _17373_, _03780_);
  nor _68830_ (_17375_, _08853_, \oc8051_golden_model_1.DPL [3]);
  nor _68831_ (_17376_, _17375_, _08854_);
  and _68832_ (_17378_, _17376_, _08847_);
  nor _68833_ (_17379_, _12627_, _08824_);
  or _68834_ (_17380_, _17379_, _17368_);
  or _68835_ (_17381_, _17380_, _04081_);
  and _68836_ (_17382_, _05303_, \oc8051_golden_model_1.ACC [3]);
  or _68837_ (_17383_, _17382_, _17368_);
  and _68838_ (_17384_, _17383_, _04409_);
  nor _68839_ (_17385_, _04409_, _17365_);
  or _68840_ (_17386_, _17385_, _03610_);
  or _68841_ (_17387_, _17386_, _17384_);
  and _68842_ (_17389_, _17387_, _03996_);
  and _68843_ (_17390_, _17389_, _17381_);
  nor _68844_ (_17391_, _08824_, _05005_);
  or _68845_ (_17392_, _17391_, _17368_);
  and _68846_ (_17393_, _17392_, _03723_);
  or _68847_ (_17394_, _17393_, _03729_);
  or _68848_ (_17395_, _17394_, _17390_);
  or _68849_ (_17396_, _17383_, _03737_);
  and _68850_ (_17397_, _17396_, _08848_);
  and _68851_ (_17398_, _17397_, _17395_);
  or _68852_ (_17400_, _17398_, _17378_);
  and _68853_ (_17401_, _17400_, _08832_);
  nor _68854_ (_17402_, _03708_, _08832_);
  or _68855_ (_17403_, _17402_, _07390_);
  or _68856_ (_17404_, _17403_, _17401_);
  or _68857_ (_17405_, _17392_, _06838_);
  and _68858_ (_17406_, _17405_, _17404_);
  or _68859_ (_17407_, _17406_, _04481_);
  and _68860_ (_17408_, _06592_, _05303_);
  or _68861_ (_17409_, _17368_, _07400_);
  or _68862_ (_17411_, _17409_, _17408_);
  and _68863_ (_17412_, _17411_, _03589_);
  and _68864_ (_17413_, _17412_, _17407_);
  nor _68865_ (_17414_, _12718_, _08824_);
  or _68866_ (_17415_, _17414_, _17368_);
  and _68867_ (_17416_, _17415_, _03222_);
  or _68868_ (_17417_, _17416_, _08828_);
  or _68869_ (_17418_, _17417_, _17413_);
  and _68870_ (_17419_, _12733_, _05303_);
  or _68871_ (_17420_, _17368_, _07766_);
  or _68872_ (_17422_, _17420_, _17419_);
  and _68873_ (_17423_, _05303_, _06276_);
  or _68874_ (_17424_, _17423_, _17368_);
  or _68875_ (_17425_, _17424_, _05886_);
  and _68876_ (_17426_, _17425_, _07778_);
  and _68877_ (_17427_, _17426_, _17422_);
  and _68878_ (_17428_, _17427_, _17418_);
  or _68879_ (_17429_, _17428_, _17374_);
  and _68880_ (_17430_, _17429_, _07777_);
  or _68881_ (_17431_, _17368_, _05567_);
  and _68882_ (_17433_, _17424_, _03622_);
  and _68883_ (_17434_, _17433_, _17431_);
  or _68884_ (_17435_, _17434_, _17430_);
  and _68885_ (_17436_, _17435_, _06828_);
  and _68886_ (_17437_, _17383_, _03790_);
  and _68887_ (_17438_, _17437_, _17431_);
  or _68888_ (_17439_, _17438_, _03624_);
  or _68889_ (_17440_, _17439_, _17436_);
  nor _68890_ (_17441_, _12732_, _08824_);
  or _68891_ (_17442_, _17368_, _07795_);
  or _68892_ (_17444_, _17442_, _17441_);
  and _68893_ (_17445_, _17444_, _07793_);
  and _68894_ (_17446_, _17445_, _17440_);
  or _68895_ (_17447_, _17446_, _17371_);
  and _68896_ (_17448_, _17447_, _04246_);
  and _68897_ (_17449_, _17380_, _03815_);
  or _68898_ (_17450_, _17449_, _03447_);
  or _68899_ (_17451_, _17450_, _17448_);
  and _68900_ (_17452_, _12794_, _05303_);
  or _68901_ (_17453_, _17368_, _03514_);
  or _68902_ (_17455_, _17453_, _17452_);
  and _68903_ (_17456_, _17455_, _43000_);
  and _68904_ (_17457_, _17456_, _17451_);
  or _68905_ (_17458_, _17457_, _17367_);
  and _68906_ (_43501_, _17458_, _41806_);
  not _68907_ (_17459_, \oc8051_golden_model_1.DPL [4]);
  nor _68908_ (_17460_, _43000_, _17459_);
  nor _68909_ (_17461_, _05303_, _17459_);
  nor _68910_ (_17462_, _12816_, _08824_);
  or _68911_ (_17463_, _17462_, _17461_);
  and _68912_ (_17465_, _17463_, _03785_);
  nor _68913_ (_17466_, _05777_, _08824_);
  or _68914_ (_17467_, _17466_, _17461_);
  or _68915_ (_17468_, _17467_, _06838_);
  nor _68916_ (_17469_, _12841_, _08824_);
  or _68917_ (_17470_, _17469_, _17461_);
  or _68918_ (_17471_, _17470_, _04081_);
  and _68919_ (_17472_, _05303_, \oc8051_golden_model_1.ACC [4]);
  or _68920_ (_17473_, _17472_, _17461_);
  and _68921_ (_17474_, _17473_, _04409_);
  nor _68922_ (_17476_, _04409_, _17459_);
  or _68923_ (_17477_, _17476_, _03610_);
  or _68924_ (_17478_, _17477_, _17474_);
  and _68925_ (_17479_, _17478_, _03996_);
  and _68926_ (_17480_, _17479_, _17471_);
  and _68927_ (_17481_, _17467_, _03723_);
  or _68928_ (_17482_, _17481_, _03729_);
  or _68929_ (_17483_, _17482_, _17480_);
  or _68930_ (_17484_, _17473_, _03737_);
  and _68931_ (_17485_, _17484_, _08848_);
  and _68932_ (_17487_, _17485_, _17483_);
  nor _68933_ (_17488_, _08854_, \oc8051_golden_model_1.DPL [4]);
  nor _68934_ (_17489_, _17488_, _08855_);
  and _68935_ (_17490_, _17489_, _08847_);
  or _68936_ (_17491_, _17490_, _17487_);
  and _68937_ (_17492_, _17491_, _08832_);
  nor _68938_ (_17493_, _06236_, _08832_);
  or _68939_ (_17494_, _17493_, _07390_);
  or _68940_ (_17495_, _17494_, _17492_);
  and _68941_ (_17496_, _17495_, _17468_);
  or _68942_ (_17498_, _17496_, _04481_);
  and _68943_ (_17499_, _06730_, _05303_);
  or _68944_ (_17500_, _17461_, _07400_);
  or _68945_ (_17501_, _17500_, _17499_);
  and _68946_ (_17502_, _17501_, _03589_);
  and _68947_ (_17503_, _17502_, _17498_);
  nor _68948_ (_17504_, _12933_, _08824_);
  or _68949_ (_17505_, _17504_, _17461_);
  and _68950_ (_17506_, _17505_, _03222_);
  or _68951_ (_17507_, _17506_, _17503_);
  or _68952_ (_17509_, _17507_, _08828_);
  and _68953_ (_17510_, _12821_, _05303_);
  or _68954_ (_17511_, _17461_, _07766_);
  or _68955_ (_17512_, _17511_, _17510_);
  and _68956_ (_17513_, _06298_, _05303_);
  or _68957_ (_17514_, _17513_, _17461_);
  or _68958_ (_17515_, _17514_, _05886_);
  and _68959_ (_17516_, _17515_, _07778_);
  and _68960_ (_17517_, _17516_, _17512_);
  and _68961_ (_17518_, _17517_, _17509_);
  and _68962_ (_17520_, _12817_, _05303_);
  or _68963_ (_17521_, _17520_, _17461_);
  and _68964_ (_17522_, _17521_, _03780_);
  or _68965_ (_17523_, _17522_, _17518_);
  and _68966_ (_17524_, _17523_, _07777_);
  or _68967_ (_17525_, _17461_, _05825_);
  and _68968_ (_17526_, _17514_, _03622_);
  and _68969_ (_17527_, _17526_, _17525_);
  or _68970_ (_17528_, _17527_, _17524_);
  and _68971_ (_17529_, _17528_, _06828_);
  and _68972_ (_17531_, _17473_, _03790_);
  and _68973_ (_17532_, _17531_, _17525_);
  or _68974_ (_17533_, _17532_, _03624_);
  or _68975_ (_17534_, _17533_, _17529_);
  nor _68976_ (_17535_, _12819_, _08824_);
  or _68977_ (_17536_, _17461_, _07795_);
  or _68978_ (_17537_, _17536_, _17535_);
  and _68979_ (_17538_, _17537_, _07793_);
  and _68980_ (_17539_, _17538_, _17534_);
  or _68981_ (_17540_, _17539_, _17465_);
  and _68982_ (_17542_, _17540_, _04246_);
  and _68983_ (_17543_, _17470_, _03815_);
  or _68984_ (_17544_, _17543_, _03447_);
  or _68985_ (_17545_, _17544_, _17542_);
  and _68986_ (_17546_, _13003_, _05303_);
  or _68987_ (_17547_, _17461_, _03514_);
  or _68988_ (_17548_, _17547_, _17546_);
  and _68989_ (_17549_, _17548_, _43000_);
  and _68990_ (_17550_, _17549_, _17545_);
  or _68991_ (_17551_, _17550_, _17460_);
  and _68992_ (_43502_, _17551_, _41806_);
  not _68993_ (_17553_, \oc8051_golden_model_1.DPL [5]);
  nor _68994_ (_17554_, _43000_, _17553_);
  nor _68995_ (_17555_, _05303_, _17553_);
  nor _68996_ (_17556_, _13146_, _08824_);
  or _68997_ (_17557_, _17556_, _17555_);
  and _68998_ (_17558_, _17557_, _03785_);
  nor _68999_ (_17559_, _05469_, _08824_);
  or _69000_ (_17560_, _17559_, _17555_);
  or _69001_ (_17561_, _17560_, _06838_);
  nor _69002_ (_17563_, _13014_, _08824_);
  or _69003_ (_17564_, _17563_, _17555_);
  or _69004_ (_17565_, _17564_, _04081_);
  and _69005_ (_17566_, _05303_, \oc8051_golden_model_1.ACC [5]);
  or _69006_ (_17567_, _17566_, _17555_);
  and _69007_ (_17568_, _17567_, _04409_);
  nor _69008_ (_17569_, _04409_, _17553_);
  or _69009_ (_17570_, _17569_, _03610_);
  or _69010_ (_17571_, _17570_, _17568_);
  and _69011_ (_17572_, _17571_, _03996_);
  and _69012_ (_17574_, _17572_, _17565_);
  and _69013_ (_17575_, _17560_, _03723_);
  or _69014_ (_17576_, _17575_, _03729_);
  or _69015_ (_17577_, _17576_, _17574_);
  or _69016_ (_17578_, _17567_, _03737_);
  and _69017_ (_17579_, _17578_, _08848_);
  and _69018_ (_17580_, _17579_, _17577_);
  nor _69019_ (_17581_, _08855_, \oc8051_golden_model_1.DPL [5]);
  nor _69020_ (_17582_, _17581_, _08856_);
  and _69021_ (_17583_, _17582_, _08847_);
  or _69022_ (_17585_, _17583_, _17580_);
  and _69023_ (_17586_, _17585_, _08832_);
  nor _69024_ (_17587_, _06267_, _08832_);
  or _69025_ (_17588_, _17587_, _07390_);
  or _69026_ (_17589_, _17588_, _17586_);
  and _69027_ (_17590_, _17589_, _17561_);
  or _69028_ (_17591_, _17590_, _04481_);
  and _69029_ (_17592_, _06684_, _05303_);
  or _69030_ (_17593_, _17555_, _07400_);
  or _69031_ (_17594_, _17593_, _17592_);
  and _69032_ (_17596_, _17594_, _03589_);
  and _69033_ (_17597_, _17596_, _17591_);
  nor _69034_ (_17598_, _13127_, _08824_);
  or _69035_ (_17599_, _17598_, _17555_);
  and _69036_ (_17600_, _17599_, _03222_);
  or _69037_ (_17601_, _17600_, _17597_);
  or _69038_ (_17602_, _17601_, _08828_);
  and _69039_ (_17603_, _13141_, _05303_);
  or _69040_ (_17604_, _17555_, _07766_);
  or _69041_ (_17605_, _17604_, _17603_);
  and _69042_ (_17607_, _06306_, _05303_);
  or _69043_ (_17608_, _17607_, _17555_);
  or _69044_ (_17609_, _17608_, _05886_);
  and _69045_ (_17610_, _17609_, _07778_);
  and _69046_ (_17611_, _17610_, _17605_);
  and _69047_ (_17612_, _17611_, _17602_);
  and _69048_ (_17613_, _13147_, _05303_);
  or _69049_ (_17614_, _17613_, _17555_);
  and _69050_ (_17615_, _17614_, _03780_);
  or _69051_ (_17616_, _17615_, _17612_);
  and _69052_ (_17618_, _17616_, _07777_);
  or _69053_ (_17619_, _17555_, _05518_);
  and _69054_ (_17620_, _17608_, _03622_);
  and _69055_ (_17621_, _17620_, _17619_);
  or _69056_ (_17622_, _17621_, _17618_);
  and _69057_ (_17623_, _17622_, _06828_);
  and _69058_ (_17624_, _17567_, _03790_);
  and _69059_ (_17625_, _17624_, _17619_);
  or _69060_ (_17626_, _17625_, _03624_);
  or _69061_ (_17627_, _17626_, _17623_);
  nor _69062_ (_17629_, _13140_, _08824_);
  or _69063_ (_17630_, _17555_, _07795_);
  or _69064_ (_17631_, _17630_, _17629_);
  and _69065_ (_17632_, _17631_, _07793_);
  and _69066_ (_17633_, _17632_, _17627_);
  or _69067_ (_17634_, _17633_, _17558_);
  and _69068_ (_17635_, _17634_, _04246_);
  and _69069_ (_17636_, _17564_, _03815_);
  or _69070_ (_17637_, _17636_, _03447_);
  or _69071_ (_17638_, _17637_, _17635_);
  and _69072_ (_17640_, _13199_, _05303_);
  or _69073_ (_17641_, _17555_, _03514_);
  or _69074_ (_17642_, _17641_, _17640_);
  and _69075_ (_17643_, _17642_, _43000_);
  and _69076_ (_17644_, _17643_, _17638_);
  or _69077_ (_17645_, _17644_, _17554_);
  and _69078_ (_43505_, _17645_, _41806_);
  not _69079_ (_17646_, \oc8051_golden_model_1.DPL [6]);
  nor _69080_ (_17647_, _43000_, _17646_);
  nor _69081_ (_17648_, _05303_, _17646_);
  nor _69082_ (_17650_, _13352_, _08824_);
  or _69083_ (_17651_, _17650_, _17648_);
  and _69084_ (_17652_, _17651_, _03785_);
  nor _69085_ (_17653_, _05363_, _08824_);
  or _69086_ (_17654_, _17653_, _17648_);
  or _69087_ (_17655_, _17654_, _06838_);
  nor _69088_ (_17656_, _13242_, _08824_);
  or _69089_ (_17657_, _17656_, _17648_);
  or _69090_ (_17658_, _17657_, _04081_);
  and _69091_ (_17659_, _05303_, \oc8051_golden_model_1.ACC [6]);
  or _69092_ (_17661_, _17659_, _17648_);
  and _69093_ (_17662_, _17661_, _04409_);
  nor _69094_ (_17663_, _04409_, _17646_);
  or _69095_ (_17664_, _17663_, _03610_);
  or _69096_ (_17665_, _17664_, _17662_);
  and _69097_ (_17666_, _17665_, _03996_);
  and _69098_ (_17667_, _17666_, _17658_);
  and _69099_ (_17668_, _17654_, _03723_);
  or _69100_ (_17669_, _17668_, _03729_);
  or _69101_ (_17670_, _17669_, _17667_);
  or _69102_ (_17672_, _17661_, _03737_);
  and _69103_ (_17673_, _17672_, _08848_);
  and _69104_ (_17674_, _17673_, _17670_);
  nor _69105_ (_17675_, _08856_, \oc8051_golden_model_1.DPL [6]);
  nor _69106_ (_17676_, _17675_, _08857_);
  and _69107_ (_17677_, _17676_, _08847_);
  or _69108_ (_17678_, _17677_, _17674_);
  and _69109_ (_17679_, _17678_, _08832_);
  nor _69110_ (_17680_, _06204_, _08832_);
  or _69111_ (_17681_, _17680_, _07390_);
  or _69112_ (_17683_, _17681_, _17679_);
  and _69113_ (_17684_, _17683_, _17655_);
  or _69114_ (_17685_, _17684_, _04481_);
  and _69115_ (_17686_, _06455_, _05303_);
  or _69116_ (_17687_, _17648_, _07400_);
  or _69117_ (_17688_, _17687_, _17686_);
  and _69118_ (_17689_, _17688_, _03589_);
  and _69119_ (_17690_, _17689_, _17685_);
  nor _69120_ (_17691_, _13332_, _08824_);
  or _69121_ (_17692_, _17691_, _17648_);
  and _69122_ (_17694_, _17692_, _03222_);
  or _69123_ (_17695_, _17694_, _17690_);
  or _69124_ (_17696_, _17695_, _08828_);
  and _69125_ (_17697_, _13347_, _05303_);
  or _69126_ (_17698_, _17648_, _07766_);
  or _69127_ (_17699_, _17698_, _17697_);
  and _69128_ (_17700_, _13339_, _05303_);
  or _69129_ (_17701_, _17700_, _17648_);
  or _69130_ (_17702_, _17701_, _05886_);
  and _69131_ (_17703_, _17702_, _07778_);
  and _69132_ (_17705_, _17703_, _17699_);
  and _69133_ (_17706_, _17705_, _17696_);
  and _69134_ (_17707_, _13353_, _05303_);
  or _69135_ (_17708_, _17707_, _17648_);
  and _69136_ (_17709_, _17708_, _03780_);
  or _69137_ (_17710_, _17709_, _17706_);
  and _69138_ (_17711_, _17710_, _07777_);
  or _69139_ (_17712_, _17648_, _05412_);
  and _69140_ (_17713_, _17701_, _03622_);
  and _69141_ (_17714_, _17713_, _17712_);
  or _69142_ (_17716_, _17714_, _17711_);
  and _69143_ (_17717_, _17716_, _06828_);
  and _69144_ (_17718_, _17661_, _03790_);
  and _69145_ (_17719_, _17718_, _17712_);
  or _69146_ (_17720_, _17719_, _03624_);
  or _69147_ (_17721_, _17720_, _17717_);
  nor _69148_ (_17722_, _13346_, _08824_);
  or _69149_ (_17723_, _17648_, _07795_);
  or _69150_ (_17724_, _17723_, _17722_);
  and _69151_ (_17725_, _17724_, _07793_);
  and _69152_ (_17727_, _17725_, _17721_);
  or _69153_ (_17728_, _17727_, _17652_);
  and _69154_ (_17729_, _17728_, _04246_);
  and _69155_ (_17730_, _17657_, _03815_);
  or _69156_ (_17731_, _17730_, _03447_);
  or _69157_ (_17732_, _17731_, _17729_);
  and _69158_ (_17733_, _13402_, _05303_);
  or _69159_ (_17734_, _17648_, _03514_);
  or _69160_ (_17735_, _17734_, _17733_);
  and _69161_ (_17736_, _17735_, _43000_);
  and _69162_ (_17738_, _17736_, _17732_);
  or _69163_ (_17739_, _17738_, _17647_);
  and _69164_ (_43506_, _17739_, _41806_);
  not _69165_ (_17740_, \oc8051_golden_model_1.DPH [0]);
  nor _69166_ (_17741_, _43000_, _17740_);
  nor _69167_ (_17742_, _08859_, \oc8051_golden_model_1.DPH [0]);
  nor _69168_ (_17743_, _17742_, _08947_);
  and _69169_ (_17744_, _17743_, _08847_);
  nor _69170_ (_17745_, _05297_, _17740_);
  nor _69171_ (_17746_, _05666_, _08921_);
  or _69172_ (_17748_, _17746_, _17745_);
  or _69173_ (_17749_, _17748_, _04081_);
  and _69174_ (_17750_, _05297_, \oc8051_golden_model_1.ACC [0]);
  or _69175_ (_17751_, _17750_, _17745_);
  and _69176_ (_17752_, _17751_, _04409_);
  nor _69177_ (_17753_, _04409_, _17740_);
  or _69178_ (_17754_, _17753_, _03610_);
  or _69179_ (_17755_, _17754_, _17752_);
  and _69180_ (_17756_, _17755_, _03996_);
  and _69181_ (_17757_, _17756_, _17749_);
  and _69182_ (_17759_, _05297_, _04620_);
  or _69183_ (_17760_, _17759_, _17745_);
  and _69184_ (_17761_, _17760_, _03723_);
  or _69185_ (_17762_, _17761_, _03729_);
  or _69186_ (_17763_, _17762_, _17757_);
  or _69187_ (_17764_, _17751_, _03737_);
  and _69188_ (_17765_, _17764_, _08848_);
  and _69189_ (_17766_, _17765_, _17763_);
  or _69190_ (_17767_, _17766_, _17744_);
  and _69191_ (_17768_, _17767_, _08832_);
  nor _69192_ (_17770_, _04048_, _08832_);
  or _69193_ (_17771_, _17770_, _07390_);
  or _69194_ (_17772_, _17771_, _17768_);
  or _69195_ (_17773_, _17760_, _06838_);
  and _69196_ (_17774_, _17773_, _17772_);
  or _69197_ (_17775_, _17774_, _04481_);
  and _69198_ (_17776_, _06546_, _05297_);
  or _69199_ (_17777_, _17745_, _07400_);
  or _69200_ (_17778_, _17777_, _17776_);
  and _69201_ (_17779_, _17778_, _17775_);
  or _69202_ (_17781_, _17779_, _03222_);
  nor _69203_ (_17782_, _12109_, _08921_);
  or _69204_ (_17783_, _17782_, _17745_);
  or _69205_ (_17784_, _17783_, _03589_);
  and _69206_ (_17785_, _17784_, _05886_);
  and _69207_ (_17786_, _17785_, _17781_);
  and _69208_ (_17787_, _05297_, _06274_);
  or _69209_ (_17788_, _17787_, _17745_);
  and _69210_ (_17789_, _17788_, _03601_);
  or _69211_ (_17790_, _17789_, _03600_);
  or _69212_ (_17792_, _17790_, _17786_);
  and _69213_ (_17793_, _12124_, _05297_);
  or _69214_ (_17794_, _17793_, _17745_);
  or _69215_ (_17795_, _17794_, _07766_);
  and _69216_ (_17796_, _17795_, _17792_);
  or _69217_ (_17797_, _17796_, _03780_);
  and _69218_ (_17798_, _12128_, _05297_);
  or _69219_ (_17799_, _17798_, _17745_);
  or _69220_ (_17800_, _17799_, _07778_);
  and _69221_ (_17801_, _17800_, _07777_);
  and _69222_ (_17803_, _17801_, _17797_);
  nand _69223_ (_17804_, _17788_, _03622_);
  nor _69224_ (_17805_, _17804_, _17746_);
  or _69225_ (_17806_, _17805_, _17803_);
  and _69226_ (_17807_, _17806_, _06828_);
  or _69227_ (_17808_, _17745_, _05666_);
  and _69228_ (_17809_, _17751_, _03790_);
  and _69229_ (_17810_, _17809_, _17808_);
  or _69230_ (_17811_, _17810_, _03624_);
  or _69231_ (_17812_, _17811_, _17807_);
  nor _69232_ (_17814_, _12122_, _08921_);
  or _69233_ (_17815_, _17745_, _07795_);
  or _69234_ (_17816_, _17815_, _17814_);
  and _69235_ (_17817_, _17816_, _07793_);
  and _69236_ (_17818_, _17817_, _17812_);
  nor _69237_ (_17819_, _12003_, _08921_);
  or _69238_ (_17820_, _17819_, _17745_);
  and _69239_ (_17821_, _17820_, _03785_);
  or _69240_ (_17822_, _17821_, _17166_);
  or _69241_ (_17823_, _17822_, _17818_);
  or _69242_ (_17825_, _17748_, _03909_);
  and _69243_ (_17826_, _17825_, _43000_);
  and _69244_ (_17827_, _17826_, _17823_);
  or _69245_ (_17828_, _17827_, _17741_);
  and _69246_ (_43507_, _17828_, _41806_);
  not _69247_ (_17829_, \oc8051_golden_model_1.DPH [1]);
  nor _69248_ (_17830_, _43000_, _17829_);
  nor _69249_ (_17831_, _05297_, _17829_);
  and _69250_ (_17832_, _05297_, _06764_);
  or _69251_ (_17833_, _17832_, _17831_);
  or _69252_ (_17835_, _17833_, _03996_);
  or _69253_ (_17836_, _05297_, \oc8051_golden_model_1.DPH [1]);
  and _69254_ (_17837_, _12213_, _05297_);
  not _69255_ (_17838_, _17837_);
  and _69256_ (_17839_, _17838_, _17836_);
  and _69257_ (_17840_, _17839_, _03610_);
  nand _69258_ (_17841_, _05297_, _03274_);
  and _69259_ (_17842_, _17841_, _17836_);
  and _69260_ (_17843_, _17842_, _04409_);
  nor _69261_ (_17844_, _04409_, _17829_);
  or _69262_ (_17846_, _17844_, _17843_);
  and _69263_ (_17847_, _17846_, _04081_);
  or _69264_ (_17848_, _17847_, _03723_);
  or _69265_ (_17849_, _17848_, _17840_);
  and _69266_ (_17850_, _17849_, _17835_);
  or _69267_ (_17851_, _17850_, _03729_);
  or _69268_ (_17852_, _17842_, _03737_);
  and _69269_ (_17853_, _17852_, _08848_);
  and _69270_ (_17854_, _17853_, _17851_);
  nor _69271_ (_17855_, _08947_, \oc8051_golden_model_1.DPH [1]);
  nor _69272_ (_17857_, _17855_, _08948_);
  and _69273_ (_17858_, _17857_, _08847_);
  or _69274_ (_17859_, _17858_, _17854_);
  and _69275_ (_17860_, _17859_, _08832_);
  nor _69276_ (_17861_, _03414_, _08832_);
  or _69277_ (_17862_, _17861_, _07390_);
  or _69278_ (_17863_, _17862_, _17860_);
  or _69279_ (_17864_, _17833_, _06838_);
  and _69280_ (_17865_, _17864_, _17863_);
  or _69281_ (_17866_, _17865_, _04481_);
  and _69282_ (_17868_, _06501_, _05297_);
  or _69283_ (_17869_, _17831_, _07400_);
  or _69284_ (_17870_, _17869_, _17868_);
  and _69285_ (_17871_, _17870_, _03589_);
  and _69286_ (_17872_, _17871_, _17866_);
  nand _69287_ (_17873_, _12313_, _05297_);
  and _69288_ (_17874_, _17836_, _03222_);
  and _69289_ (_17875_, _17874_, _17873_);
  or _69290_ (_17876_, _17875_, _17872_);
  and _69291_ (_17877_, _17876_, _03602_);
  or _69292_ (_17879_, _12327_, _08921_);
  and _69293_ (_17880_, _17879_, _03600_);
  nand _69294_ (_17881_, _05297_, _04303_);
  and _69295_ (_17882_, _17881_, _03601_);
  or _69296_ (_17883_, _17882_, _17880_);
  and _69297_ (_17884_, _17883_, _17836_);
  or _69298_ (_17885_, _17884_, _17877_);
  and _69299_ (_17886_, _17885_, _07778_);
  or _69300_ (_17887_, _12333_, _08921_);
  and _69301_ (_17888_, _17836_, _03780_);
  and _69302_ (_17890_, _17888_, _17887_);
  or _69303_ (_17891_, _17890_, _17886_);
  and _69304_ (_17892_, _17891_, _07777_);
  or _69305_ (_17893_, _12207_, _08921_);
  and _69306_ (_17894_, _17836_, _03622_);
  and _69307_ (_17895_, _17894_, _17893_);
  or _69308_ (_17896_, _17895_, _17892_);
  and _69309_ (_17897_, _17896_, _06828_);
  or _69310_ (_17898_, _17831_, _05618_);
  and _69311_ (_17899_, _17842_, _03790_);
  and _69312_ (_17901_, _17899_, _17898_);
  or _69313_ (_17902_, _17901_, _17897_);
  and _69314_ (_17903_, _17902_, _03786_);
  or _69315_ (_17904_, _17881_, _05618_);
  and _69316_ (_17905_, _17836_, _03624_);
  and _69317_ (_17906_, _17905_, _17904_);
  or _69318_ (_17907_, _17841_, _05618_);
  and _69319_ (_17908_, _17836_, _03785_);
  and _69320_ (_17909_, _17908_, _17907_);
  or _69321_ (_17910_, _17909_, _03815_);
  or _69322_ (_17912_, _17910_, _17906_);
  or _69323_ (_17913_, _17912_, _17903_);
  or _69324_ (_17914_, _17839_, _04246_);
  and _69325_ (_17915_, _17914_, _17913_);
  or _69326_ (_17916_, _17915_, _03447_);
  or _69327_ (_17917_, _17831_, _03514_);
  or _69328_ (_17918_, _17917_, _17837_);
  and _69329_ (_17919_, _17918_, _43000_);
  and _69330_ (_17920_, _17919_, _17916_);
  or _69331_ (_17921_, _17920_, _17830_);
  and _69332_ (_43510_, _17921_, _41806_);
  not _69333_ (_17923_, \oc8051_golden_model_1.DPH [2]);
  nor _69334_ (_17924_, _43000_, _17923_);
  nor _69335_ (_17925_, _05297_, _17923_);
  nor _69336_ (_17926_, _12538_, _08921_);
  or _69337_ (_17927_, _17926_, _17925_);
  and _69338_ (_17928_, _17927_, _03785_);
  and _69339_ (_17929_, _12539_, _05297_);
  or _69340_ (_17930_, _17929_, _17925_);
  and _69341_ (_17931_, _17930_, _03780_);
  nor _69342_ (_17933_, _08921_, _04875_);
  or _69343_ (_17934_, _17933_, _17925_);
  or _69344_ (_17935_, _17934_, _06838_);
  nor _69345_ (_17936_, _12416_, _08921_);
  or _69346_ (_17937_, _17936_, _17925_);
  or _69347_ (_17938_, _17937_, _04081_);
  and _69348_ (_17939_, _05297_, \oc8051_golden_model_1.ACC [2]);
  or _69349_ (_17940_, _17939_, _17925_);
  and _69350_ (_17941_, _17940_, _04409_);
  nor _69351_ (_17942_, _04409_, _17923_);
  or _69352_ (_17944_, _17942_, _03610_);
  or _69353_ (_17945_, _17944_, _17941_);
  and _69354_ (_17946_, _17945_, _03996_);
  and _69355_ (_17947_, _17946_, _17938_);
  and _69356_ (_17948_, _17934_, _03723_);
  or _69357_ (_17949_, _17948_, _03729_);
  or _69358_ (_17950_, _17949_, _17947_);
  or _69359_ (_17951_, _17940_, _03737_);
  and _69360_ (_17952_, _17951_, _08848_);
  and _69361_ (_17953_, _17952_, _17950_);
  or _69362_ (_17955_, _08948_, \oc8051_golden_model_1.DPH [2]);
  nor _69363_ (_17956_, _08949_, _08848_);
  and _69364_ (_17957_, _17956_, _17955_);
  or _69365_ (_17958_, _17957_, _17953_);
  and _69366_ (_17959_, _17958_, _08832_);
  nor _69367_ (_17960_, _03904_, _08832_);
  or _69368_ (_17961_, _17960_, _07390_);
  or _69369_ (_17962_, _17961_, _17959_);
  and _69370_ (_17963_, _17962_, _17935_);
  or _69371_ (_17964_, _17963_, _04481_);
  and _69372_ (_17966_, _06637_, _05297_);
  or _69373_ (_17967_, _17925_, _07400_);
  or _69374_ (_17968_, _17967_, _17966_);
  and _69375_ (_17969_, _17968_, _03589_);
  and _69376_ (_17970_, _17969_, _17964_);
  nor _69377_ (_17971_, _12519_, _08921_);
  or _69378_ (_17972_, _17971_, _17925_);
  and _69379_ (_17973_, _17972_, _03222_);
  or _69380_ (_17974_, _17973_, _17970_);
  or _69381_ (_17975_, _17974_, _08828_);
  and _69382_ (_17977_, _12533_, _05297_);
  or _69383_ (_17978_, _17925_, _07766_);
  or _69384_ (_17979_, _17978_, _17977_);
  and _69385_ (_17980_, _05297_, _06332_);
  or _69386_ (_17981_, _17980_, _17925_);
  or _69387_ (_17982_, _17981_, _05886_);
  and _69388_ (_17983_, _17982_, _07778_);
  and _69389_ (_17984_, _17983_, _17979_);
  and _69390_ (_17985_, _17984_, _17975_);
  or _69391_ (_17986_, _17985_, _17931_);
  and _69392_ (_17988_, _17986_, _07777_);
  or _69393_ (_17989_, _17925_, _05718_);
  and _69394_ (_17990_, _17981_, _03622_);
  and _69395_ (_17991_, _17990_, _17989_);
  or _69396_ (_17992_, _17991_, _17988_);
  and _69397_ (_17993_, _17992_, _06828_);
  and _69398_ (_17994_, _17940_, _03790_);
  and _69399_ (_17995_, _17994_, _17989_);
  or _69400_ (_17996_, _17995_, _03624_);
  or _69401_ (_17997_, _17996_, _17993_);
  nor _69402_ (_17999_, _12532_, _08921_);
  or _69403_ (_18000_, _17925_, _07795_);
  or _69404_ (_18001_, _18000_, _17999_);
  and _69405_ (_18002_, _18001_, _07793_);
  and _69406_ (_18003_, _18002_, _17997_);
  or _69407_ (_18004_, _18003_, _17928_);
  and _69408_ (_18005_, _18004_, _04246_);
  and _69409_ (_18006_, _17937_, _03815_);
  or _69410_ (_18007_, _18006_, _03447_);
  or _69411_ (_18008_, _18007_, _18005_);
  and _69412_ (_18010_, _12592_, _05297_);
  or _69413_ (_18011_, _17925_, _03514_);
  or _69414_ (_18012_, _18011_, _18010_);
  and _69415_ (_18013_, _18012_, _43000_);
  and _69416_ (_18014_, _18013_, _18008_);
  or _69417_ (_18015_, _18014_, _17924_);
  and _69418_ (_43511_, _18015_, _41806_);
  not _69419_ (_18016_, \oc8051_golden_model_1.DPH [3]);
  nor _69420_ (_18017_, _43000_, _18016_);
  nor _69421_ (_18018_, _05297_, _18016_);
  nor _69422_ (_18020_, _12738_, _08921_);
  or _69423_ (_18021_, _18020_, _18018_);
  and _69424_ (_18022_, _18021_, _03785_);
  and _69425_ (_18023_, _12739_, _05297_);
  or _69426_ (_18024_, _18023_, _18018_);
  and _69427_ (_18025_, _18024_, _03780_);
  nor _69428_ (_18026_, _12627_, _08921_);
  or _69429_ (_18027_, _18026_, _18018_);
  or _69430_ (_18028_, _18027_, _04081_);
  and _69431_ (_18029_, _05297_, \oc8051_golden_model_1.ACC [3]);
  or _69432_ (_18031_, _18029_, _18018_);
  and _69433_ (_18032_, _18031_, _04409_);
  nor _69434_ (_18033_, _04409_, _18016_);
  or _69435_ (_18034_, _18033_, _03610_);
  or _69436_ (_18035_, _18034_, _18032_);
  and _69437_ (_18036_, _18035_, _03996_);
  and _69438_ (_18037_, _18036_, _18028_);
  nor _69439_ (_18038_, _08921_, _05005_);
  or _69440_ (_18039_, _18038_, _18018_);
  and _69441_ (_18040_, _18039_, _03723_);
  or _69442_ (_18042_, _18040_, _03729_);
  or _69443_ (_18043_, _18042_, _18037_);
  or _69444_ (_18044_, _18031_, _03737_);
  and _69445_ (_18045_, _18044_, _08848_);
  and _69446_ (_18046_, _18045_, _18043_);
  or _69447_ (_18047_, _08949_, \oc8051_golden_model_1.DPH [3]);
  nor _69448_ (_18048_, _08950_, _08848_);
  and _69449_ (_18049_, _18048_, _18047_);
  or _69450_ (_18050_, _18049_, _18046_);
  and _69451_ (_18051_, _18050_, _08832_);
  nor _69452_ (_18053_, _08832_, _03581_);
  or _69453_ (_18054_, _18053_, _07390_);
  or _69454_ (_18055_, _18054_, _18051_);
  or _69455_ (_18056_, _18039_, _06838_);
  and _69456_ (_18057_, _18056_, _18055_);
  or _69457_ (_18058_, _18057_, _04481_);
  and _69458_ (_18059_, _06592_, _05297_);
  or _69459_ (_18060_, _18018_, _07400_);
  or _69460_ (_18061_, _18060_, _18059_);
  and _69461_ (_18062_, _18061_, _03589_);
  and _69462_ (_18064_, _18062_, _18058_);
  nor _69463_ (_18065_, _12718_, _08921_);
  or _69464_ (_18066_, _18065_, _18018_);
  and _69465_ (_18067_, _18066_, _03222_);
  or _69466_ (_18068_, _18067_, _08828_);
  or _69467_ (_18069_, _18068_, _18064_);
  and _69468_ (_18070_, _12733_, _05297_);
  or _69469_ (_18071_, _18018_, _07766_);
  or _69470_ (_18072_, _18071_, _18070_);
  and _69471_ (_18073_, _05297_, _06276_);
  or _69472_ (_18075_, _18073_, _18018_);
  or _69473_ (_18076_, _18075_, _05886_);
  and _69474_ (_18077_, _18076_, _07778_);
  and _69475_ (_18078_, _18077_, _18072_);
  and _69476_ (_18079_, _18078_, _18069_);
  or _69477_ (_18080_, _18079_, _18025_);
  and _69478_ (_18081_, _18080_, _07777_);
  or _69479_ (_18082_, _18018_, _05567_);
  and _69480_ (_18083_, _18075_, _03622_);
  and _69481_ (_18084_, _18083_, _18082_);
  or _69482_ (_18086_, _18084_, _18081_);
  and _69483_ (_18087_, _18086_, _06828_);
  and _69484_ (_18088_, _18031_, _03790_);
  and _69485_ (_18089_, _18088_, _18082_);
  or _69486_ (_18090_, _18089_, _03624_);
  or _69487_ (_18091_, _18090_, _18087_);
  nor _69488_ (_18092_, _12732_, _08921_);
  or _69489_ (_18093_, _18018_, _07795_);
  or _69490_ (_18094_, _18093_, _18092_);
  and _69491_ (_18095_, _18094_, _07793_);
  and _69492_ (_18097_, _18095_, _18091_);
  or _69493_ (_18098_, _18097_, _18022_);
  and _69494_ (_18099_, _18098_, _04246_);
  and _69495_ (_18100_, _18027_, _03815_);
  or _69496_ (_18101_, _18100_, _03447_);
  or _69497_ (_18102_, _18101_, _18099_);
  and _69498_ (_18103_, _12794_, _05297_);
  or _69499_ (_18104_, _18018_, _03514_);
  or _69500_ (_18105_, _18104_, _18103_);
  and _69501_ (_18106_, _18105_, _43000_);
  and _69502_ (_18108_, _18106_, _18102_);
  or _69503_ (_18109_, _18108_, _18017_);
  and _69504_ (_43512_, _18109_, _41806_);
  not _69505_ (_18110_, \oc8051_golden_model_1.DPH [4]);
  nor _69506_ (_18111_, _43000_, _18110_);
  nor _69507_ (_18112_, _05297_, _18110_);
  nor _69508_ (_18113_, _12816_, _08921_);
  or _69509_ (_18114_, _18113_, _18112_);
  and _69510_ (_18115_, _18114_, _03785_);
  nor _69511_ (_18116_, _05777_, _08921_);
  or _69512_ (_18118_, _18116_, _18112_);
  or _69513_ (_18119_, _18118_, _06838_);
  nor _69514_ (_18120_, _12841_, _08921_);
  or _69515_ (_18121_, _18120_, _18112_);
  or _69516_ (_18122_, _18121_, _04081_);
  and _69517_ (_18123_, _05297_, \oc8051_golden_model_1.ACC [4]);
  or _69518_ (_18124_, _18123_, _18112_);
  and _69519_ (_18125_, _18124_, _04409_);
  nor _69520_ (_18126_, _04409_, _18110_);
  or _69521_ (_18127_, _18126_, _03610_);
  or _69522_ (_18129_, _18127_, _18125_);
  and _69523_ (_18130_, _18129_, _03996_);
  and _69524_ (_18131_, _18130_, _18122_);
  and _69525_ (_18132_, _18118_, _03723_);
  or _69526_ (_18133_, _18132_, _03729_);
  or _69527_ (_18134_, _18133_, _18131_);
  or _69528_ (_18135_, _18124_, _03737_);
  and _69529_ (_18136_, _18135_, _08848_);
  and _69530_ (_18137_, _18136_, _18134_);
  or _69531_ (_18138_, _08950_, \oc8051_golden_model_1.DPH [4]);
  nor _69532_ (_18140_, _08951_, _08848_);
  and _69533_ (_18141_, _18140_, _18138_);
  or _69534_ (_18142_, _18141_, _18137_);
  and _69535_ (_18143_, _18142_, _08832_);
  nor _69536_ (_18144_, _03486_, _08832_);
  or _69537_ (_18145_, _18144_, _07390_);
  or _69538_ (_18146_, _18145_, _18143_);
  and _69539_ (_18147_, _18146_, _18119_);
  or _69540_ (_18148_, _18147_, _04481_);
  and _69541_ (_18149_, _06730_, _05297_);
  or _69542_ (_18151_, _18112_, _07400_);
  or _69543_ (_18152_, _18151_, _18149_);
  and _69544_ (_18153_, _18152_, _03589_);
  and _69545_ (_18154_, _18153_, _18148_);
  nor _69546_ (_18155_, _12933_, _08921_);
  or _69547_ (_18156_, _18155_, _18112_);
  and _69548_ (_18157_, _18156_, _03222_);
  or _69549_ (_18158_, _18157_, _18154_);
  or _69550_ (_18159_, _18158_, _08828_);
  and _69551_ (_18160_, _12821_, _05297_);
  or _69552_ (_18162_, _18112_, _07766_);
  or _69553_ (_18163_, _18162_, _18160_);
  and _69554_ (_18164_, _06298_, _05297_);
  or _69555_ (_18165_, _18164_, _18112_);
  or _69556_ (_18166_, _18165_, _05886_);
  and _69557_ (_18167_, _18166_, _07778_);
  and _69558_ (_18168_, _18167_, _18163_);
  and _69559_ (_18169_, _18168_, _18159_);
  and _69560_ (_18170_, _12817_, _05297_);
  or _69561_ (_18171_, _18170_, _18112_);
  and _69562_ (_18173_, _18171_, _03780_);
  or _69563_ (_18174_, _18173_, _18169_);
  and _69564_ (_18175_, _18174_, _07777_);
  or _69565_ (_18176_, _18112_, _05825_);
  and _69566_ (_18177_, _18165_, _03622_);
  and _69567_ (_18178_, _18177_, _18176_);
  or _69568_ (_18179_, _18178_, _18175_);
  and _69569_ (_18180_, _18179_, _06828_);
  and _69570_ (_18181_, _18124_, _03790_);
  and _69571_ (_18182_, _18181_, _18176_);
  or _69572_ (_18184_, _18182_, _03624_);
  or _69573_ (_18185_, _18184_, _18180_);
  nor _69574_ (_18186_, _12819_, _08921_);
  or _69575_ (_18187_, _18112_, _07795_);
  or _69576_ (_18188_, _18187_, _18186_);
  and _69577_ (_18189_, _18188_, _07793_);
  and _69578_ (_18190_, _18189_, _18185_);
  or _69579_ (_18191_, _18190_, _18115_);
  and _69580_ (_18192_, _18191_, _04246_);
  and _69581_ (_18193_, _18121_, _03815_);
  or _69582_ (_18195_, _18193_, _03447_);
  or _69583_ (_18196_, _18195_, _18192_);
  and _69584_ (_18197_, _13003_, _05297_);
  or _69585_ (_18198_, _18112_, _03514_);
  or _69586_ (_18199_, _18198_, _18197_);
  and _69587_ (_18200_, _18199_, _43000_);
  and _69588_ (_18201_, _18200_, _18196_);
  or _69589_ (_18202_, _18201_, _18111_);
  and _69590_ (_43513_, _18202_, _41806_);
  not _69591_ (_18203_, \oc8051_golden_model_1.DPH [5]);
  nor _69592_ (_18205_, _43000_, _18203_);
  nor _69593_ (_18206_, _05297_, _18203_);
  nor _69594_ (_18207_, _13146_, _08921_);
  or _69595_ (_18208_, _18207_, _18206_);
  and _69596_ (_18209_, _18208_, _03785_);
  nor _69597_ (_18210_, _05469_, _08921_);
  or _69598_ (_18211_, _18210_, _18206_);
  or _69599_ (_18212_, _18211_, _06838_);
  nor _69600_ (_18213_, _13014_, _08921_);
  or _69601_ (_18214_, _18213_, _18206_);
  or _69602_ (_18216_, _18214_, _04081_);
  and _69603_ (_18217_, _05297_, \oc8051_golden_model_1.ACC [5]);
  or _69604_ (_18218_, _18217_, _18206_);
  and _69605_ (_18219_, _18218_, _04409_);
  nor _69606_ (_18220_, _04409_, _18203_);
  or _69607_ (_18221_, _18220_, _03610_);
  or _69608_ (_18222_, _18221_, _18219_);
  and _69609_ (_18223_, _18222_, _03996_);
  and _69610_ (_18224_, _18223_, _18216_);
  and _69611_ (_18225_, _18211_, _03723_);
  or _69612_ (_18227_, _18225_, _03729_);
  or _69613_ (_18228_, _18227_, _18224_);
  or _69614_ (_18229_, _18218_, _03737_);
  and _69615_ (_18230_, _18229_, _08848_);
  and _69616_ (_18231_, _18230_, _18228_);
  or _69617_ (_18232_, _08951_, \oc8051_golden_model_1.DPH [5]);
  nor _69618_ (_18233_, _08952_, _08848_);
  and _69619_ (_18234_, _18233_, _18232_);
  or _69620_ (_18235_, _18234_, _18231_);
  and _69621_ (_18236_, _18235_, _08832_);
  nor _69622_ (_18238_, _03860_, _08832_);
  or _69623_ (_18239_, _18238_, _07390_);
  or _69624_ (_18240_, _18239_, _18236_);
  and _69625_ (_18241_, _18240_, _18212_);
  or _69626_ (_18242_, _18241_, _04481_);
  and _69627_ (_18243_, _06684_, _05297_);
  or _69628_ (_18244_, _18206_, _07400_);
  or _69629_ (_18245_, _18244_, _18243_);
  and _69630_ (_18246_, _18245_, _03589_);
  and _69631_ (_18247_, _18246_, _18242_);
  nor _69632_ (_18249_, _13127_, _08921_);
  or _69633_ (_18250_, _18249_, _18206_);
  and _69634_ (_18251_, _18250_, _03222_);
  or _69635_ (_18252_, _18251_, _18247_);
  or _69636_ (_18253_, _18252_, _08828_);
  and _69637_ (_18254_, _13141_, _05297_);
  or _69638_ (_18255_, _18206_, _07766_);
  or _69639_ (_18256_, _18255_, _18254_);
  and _69640_ (_18257_, _06306_, _05297_);
  or _69641_ (_18258_, _18257_, _18206_);
  or _69642_ (_18260_, _18258_, _05886_);
  and _69643_ (_18261_, _18260_, _07778_);
  and _69644_ (_18262_, _18261_, _18256_);
  and _69645_ (_18263_, _18262_, _18253_);
  and _69646_ (_18264_, _13147_, _05297_);
  or _69647_ (_18265_, _18264_, _18206_);
  and _69648_ (_18266_, _18265_, _03780_);
  or _69649_ (_18267_, _18266_, _18263_);
  and _69650_ (_18268_, _18267_, _07777_);
  or _69651_ (_18269_, _18206_, _05518_);
  and _69652_ (_18271_, _18258_, _03622_);
  and _69653_ (_18272_, _18271_, _18269_);
  or _69654_ (_18273_, _18272_, _18268_);
  and _69655_ (_18274_, _18273_, _06828_);
  and _69656_ (_18275_, _18218_, _03790_);
  and _69657_ (_18276_, _18275_, _18269_);
  or _69658_ (_18277_, _18276_, _03624_);
  or _69659_ (_18278_, _18277_, _18274_);
  nor _69660_ (_18279_, _13140_, _08921_);
  or _69661_ (_18280_, _18206_, _07795_);
  or _69662_ (_18282_, _18280_, _18279_);
  and _69663_ (_18283_, _18282_, _07793_);
  and _69664_ (_18284_, _18283_, _18278_);
  or _69665_ (_18285_, _18284_, _18209_);
  and _69666_ (_18286_, _18285_, _04246_);
  and _69667_ (_18287_, _18214_, _03815_);
  or _69668_ (_18288_, _18287_, _03447_);
  or _69669_ (_18289_, _18288_, _18286_);
  and _69670_ (_18290_, _13199_, _05297_);
  or _69671_ (_18291_, _18206_, _03514_);
  or _69672_ (_18293_, _18291_, _18290_);
  and _69673_ (_18294_, _18293_, _43000_);
  and _69674_ (_18295_, _18294_, _18289_);
  or _69675_ (_18296_, _18295_, _18205_);
  and _69676_ (_43514_, _18296_, _41806_);
  not _69677_ (_18297_, \oc8051_golden_model_1.DPH [6]);
  nor _69678_ (_18298_, _43000_, _18297_);
  nor _69679_ (_18299_, _05297_, _18297_);
  nor _69680_ (_18300_, _13352_, _08921_);
  or _69681_ (_18301_, _18300_, _18299_);
  and _69682_ (_18303_, _18301_, _03785_);
  nor _69683_ (_18304_, _05363_, _08921_);
  or _69684_ (_18305_, _18304_, _18299_);
  or _69685_ (_18306_, _18305_, _06838_);
  nor _69686_ (_18307_, _13242_, _08921_);
  or _69687_ (_18308_, _18307_, _18299_);
  or _69688_ (_18309_, _18308_, _04081_);
  and _69689_ (_18310_, _05297_, \oc8051_golden_model_1.ACC [6]);
  or _69690_ (_18311_, _18310_, _18299_);
  and _69691_ (_18312_, _18311_, _04409_);
  nor _69692_ (_18314_, _04409_, _18297_);
  or _69693_ (_18315_, _18314_, _03610_);
  or _69694_ (_18316_, _18315_, _18312_);
  and _69695_ (_18317_, _18316_, _03996_);
  and _69696_ (_18318_, _18317_, _18309_);
  and _69697_ (_18319_, _18305_, _03723_);
  or _69698_ (_18320_, _18319_, _03729_);
  or _69699_ (_18321_, _18320_, _18318_);
  or _69700_ (_18322_, _18311_, _03737_);
  and _69701_ (_18323_, _18322_, _08848_);
  and _69702_ (_18325_, _18323_, _18321_);
  or _69703_ (_18326_, _08952_, \oc8051_golden_model_1.DPH [6]);
  nor _69704_ (_18327_, _08953_, _08848_);
  and _69705_ (_18328_, _18327_, _18326_);
  or _69706_ (_18329_, _18328_, _18325_);
  and _69707_ (_18330_, _18329_, _08832_);
  nor _69708_ (_18331_, _08832_, _03549_);
  or _69709_ (_18332_, _18331_, _07390_);
  or _69710_ (_18333_, _18332_, _18330_);
  and _69711_ (_18334_, _18333_, _18306_);
  or _69712_ (_18336_, _18334_, _04481_);
  and _69713_ (_18337_, _06455_, _05297_);
  or _69714_ (_18338_, _18299_, _07400_);
  or _69715_ (_18339_, _18338_, _18337_);
  and _69716_ (_18340_, _18339_, _03589_);
  and _69717_ (_18341_, _18340_, _18336_);
  nor _69718_ (_18342_, _13332_, _08921_);
  or _69719_ (_18343_, _18342_, _18299_);
  and _69720_ (_18344_, _18343_, _03222_);
  or _69721_ (_18345_, _18344_, _18341_);
  or _69722_ (_18347_, _18345_, _08828_);
  and _69723_ (_18348_, _13347_, _05297_);
  or _69724_ (_18349_, _18299_, _07766_);
  or _69725_ (_18350_, _18349_, _18348_);
  and _69726_ (_18351_, _13339_, _05297_);
  or _69727_ (_18352_, _18351_, _18299_);
  or _69728_ (_18353_, _18352_, _05886_);
  and _69729_ (_18354_, _18353_, _07778_);
  and _69730_ (_18355_, _18354_, _18350_);
  and _69731_ (_18356_, _18355_, _18347_);
  and _69732_ (_18358_, _13353_, _05297_);
  or _69733_ (_18359_, _18358_, _18299_);
  and _69734_ (_18360_, _18359_, _03780_);
  or _69735_ (_18361_, _18360_, _18356_);
  and _69736_ (_18362_, _18361_, _07777_);
  or _69737_ (_18363_, _18299_, _05412_);
  and _69738_ (_18364_, _18352_, _03622_);
  and _69739_ (_18365_, _18364_, _18363_);
  or _69740_ (_18366_, _18365_, _18362_);
  and _69741_ (_18367_, _18366_, _06828_);
  and _69742_ (_18369_, _18311_, _03790_);
  and _69743_ (_18370_, _18369_, _18363_);
  or _69744_ (_18371_, _18370_, _03624_);
  or _69745_ (_18372_, _18371_, _18367_);
  nor _69746_ (_18373_, _13346_, _08921_);
  or _69747_ (_18374_, _18299_, _07795_);
  or _69748_ (_18375_, _18374_, _18373_);
  and _69749_ (_18376_, _18375_, _07793_);
  and _69750_ (_18377_, _18376_, _18372_);
  or _69751_ (_18378_, _18377_, _18303_);
  and _69752_ (_18380_, _18378_, _04246_);
  and _69753_ (_18381_, _18308_, _03815_);
  or _69754_ (_18382_, _18381_, _03447_);
  or _69755_ (_18383_, _18382_, _18380_);
  and _69756_ (_18384_, _13402_, _05297_);
  or _69757_ (_18385_, _18299_, _03514_);
  or _69758_ (_18386_, _18385_, _18384_);
  and _69759_ (_18387_, _18386_, _43000_);
  and _69760_ (_18388_, _18387_, _18383_);
  or _69761_ (_18389_, _18388_, _18298_);
  and _69762_ (_43515_, _18389_, _41806_);
  not _69763_ (_18391_, \oc8051_golden_model_1.IE [0]);
  nor _69764_ (_18392_, _05229_, _18391_);
  nor _69765_ (_18393_, _05666_, _09021_);
  nor _69766_ (_18394_, _18393_, _18392_);
  and _69767_ (_18395_, _18394_, _03447_);
  and _69768_ (_18396_, _12128_, _05229_);
  nor _69769_ (_18397_, _18396_, _18392_);
  nor _69770_ (_18398_, _18397_, _07778_);
  and _69771_ (_18399_, _05229_, _06274_);
  nor _69772_ (_18401_, _18399_, _18392_);
  and _69773_ (_18402_, _18401_, _03601_);
  and _69774_ (_18403_, _05229_, _04620_);
  nor _69775_ (_18404_, _18403_, _18392_);
  and _69776_ (_18405_, _18404_, _07390_);
  and _69777_ (_18406_, _05229_, \oc8051_golden_model_1.ACC [0]);
  nor _69778_ (_18407_, _18406_, _18392_);
  nor _69779_ (_18408_, _18407_, _09029_);
  nor _69780_ (_18409_, _04409_, _18391_);
  or _69781_ (_18410_, _18409_, _18408_);
  and _69782_ (_18412_, _18410_, _04081_);
  nor _69783_ (_18413_, _18394_, _04081_);
  or _69784_ (_18414_, _18413_, _18412_);
  and _69785_ (_18415_, _18414_, _04055_);
  nor _69786_ (_18416_, _05924_, _18391_);
  and _69787_ (_18417_, _12021_, _05924_);
  nor _69788_ (_18418_, _18417_, _18416_);
  nor _69789_ (_18419_, _18418_, _04055_);
  nor _69790_ (_18420_, _18419_, _18415_);
  nor _69791_ (_18421_, _18420_, _03723_);
  nor _69792_ (_18423_, _18404_, _03996_);
  or _69793_ (_18424_, _18423_, _18421_);
  and _69794_ (_18425_, _18424_, _03737_);
  nor _69795_ (_18426_, _18407_, _03737_);
  or _69796_ (_18427_, _18426_, _18425_);
  and _69797_ (_18428_, _18427_, _03736_);
  and _69798_ (_18429_, _18392_, _03714_);
  or _69799_ (_18430_, _18429_, _18428_);
  and _69800_ (_18431_, _18430_, _06840_);
  nor _69801_ (_18432_, _18394_, _06840_);
  or _69802_ (_18434_, _18432_, _18431_);
  and _69803_ (_18435_, _18434_, _03710_);
  nor _69804_ (_18436_, _12052_, _09059_);
  nor _69805_ (_18437_, _18436_, _18416_);
  nor _69806_ (_18438_, _18437_, _03710_);
  or _69807_ (_18439_, _18438_, _07390_);
  nor _69808_ (_18440_, _18439_, _18435_);
  nor _69809_ (_18441_, _18440_, _18405_);
  nor _69810_ (_18442_, _18441_, _04481_);
  and _69811_ (_18443_, _06546_, _05229_);
  nor _69812_ (_18445_, _18392_, _07400_);
  not _69813_ (_18446_, _18445_);
  nor _69814_ (_18447_, _18446_, _18443_);
  or _69815_ (_18448_, _18447_, _03222_);
  nor _69816_ (_18449_, _18448_, _18442_);
  nor _69817_ (_18450_, _12109_, _09021_);
  nor _69818_ (_18451_, _18450_, _18392_);
  nor _69819_ (_18452_, _18451_, _03589_);
  or _69820_ (_18453_, _18452_, _03601_);
  nor _69821_ (_18454_, _18453_, _18449_);
  nor _69822_ (_18456_, _18454_, _18402_);
  or _69823_ (_18457_, _18456_, _03600_);
  and _69824_ (_18458_, _12124_, _05229_);
  or _69825_ (_18459_, _18458_, _18392_);
  or _69826_ (_18460_, _18459_, _07766_);
  and _69827_ (_18461_, _18460_, _07778_);
  and _69828_ (_18462_, _18461_, _18457_);
  nor _69829_ (_18463_, _18462_, _18398_);
  nor _69830_ (_18464_, _18463_, _03622_);
  or _69831_ (_18465_, _18401_, _07777_);
  nor _69832_ (_18467_, _18465_, _18393_);
  nor _69833_ (_18468_, _18467_, _18464_);
  nor _69834_ (_18469_, _18468_, _03790_);
  and _69835_ (_18470_, _12005_, _05229_);
  or _69836_ (_18471_, _18470_, _18392_);
  and _69837_ (_18472_, _18471_, _03790_);
  or _69838_ (_18473_, _18472_, _18469_);
  and _69839_ (_18474_, _18473_, _07795_);
  nor _69840_ (_18475_, _12122_, _09021_);
  nor _69841_ (_18476_, _18475_, _18392_);
  nor _69842_ (_18478_, _18476_, _07795_);
  or _69843_ (_18479_, _18478_, _18474_);
  and _69844_ (_18480_, _18479_, _07793_);
  nor _69845_ (_18481_, _12003_, _09021_);
  nor _69846_ (_18482_, _18481_, _18392_);
  nor _69847_ (_18483_, _18482_, _07793_);
  or _69848_ (_18484_, _18483_, _18480_);
  and _69849_ (_18485_, _18484_, _04246_);
  nor _69850_ (_18486_, _18394_, _04246_);
  or _69851_ (_18487_, _18486_, _18485_);
  and _69852_ (_18489_, _18487_, _03823_);
  and _69853_ (_18490_, _18392_, _03453_);
  nor _69854_ (_18491_, _18490_, _03447_);
  not _69855_ (_18492_, _18491_);
  nor _69856_ (_18493_, _18492_, _18489_);
  nor _69857_ (_18494_, _18493_, _18395_);
  or _69858_ (_18495_, _18494_, _43004_);
  or _69859_ (_18496_, _43000_, \oc8051_golden_model_1.IE [0]);
  and _69860_ (_18497_, _18496_, _41806_);
  and _69861_ (_43516_, _18497_, _18495_);
  not _69862_ (_18499_, _03786_);
  not _69863_ (_18500_, \oc8051_golden_model_1.IE [1]);
  nor _69864_ (_18501_, _05229_, _18500_);
  and _69865_ (_18502_, _06501_, _05229_);
  or _69866_ (_18503_, _18502_, _18501_);
  and _69867_ (_18504_, _18503_, _04481_);
  nor _69868_ (_18505_, _05229_, \oc8051_golden_model_1.IE [1]);
  and _69869_ (_18506_, _05229_, _03274_);
  nor _69870_ (_18507_, _18506_, _18505_);
  and _69871_ (_18508_, _18507_, _04409_);
  nor _69872_ (_18510_, _04409_, _18500_);
  or _69873_ (_18511_, _18510_, _18508_);
  and _69874_ (_18512_, _18511_, _04081_);
  and _69875_ (_18513_, _12213_, _05229_);
  nor _69876_ (_18514_, _18513_, _18505_);
  and _69877_ (_18515_, _18514_, _03610_);
  or _69878_ (_18516_, _18515_, _18512_);
  and _69879_ (_18517_, _18516_, _04055_);
  and _69880_ (_18518_, _12224_, _05924_);
  nor _69881_ (_18519_, _05924_, _18500_);
  or _69882_ (_18521_, _18519_, _03723_);
  or _69883_ (_18522_, _18521_, _18518_);
  and _69884_ (_18523_, _18522_, _14265_);
  nor _69885_ (_18524_, _18523_, _18517_);
  and _69886_ (_18525_, _05229_, _06764_);
  nor _69887_ (_18526_, _18525_, _18501_);
  and _69888_ (_18527_, _18526_, _03723_);
  nor _69889_ (_18528_, _18527_, _18524_);
  and _69890_ (_18529_, _18528_, _03737_);
  and _69891_ (_18530_, _18507_, _03729_);
  or _69892_ (_18532_, _18530_, _18529_);
  and _69893_ (_18533_, _18532_, _03736_);
  and _69894_ (_18534_, _12211_, _05924_);
  nor _69895_ (_18535_, _18534_, _18519_);
  nor _69896_ (_18536_, _18535_, _03736_);
  or _69897_ (_18537_, _18536_, _03719_);
  or _69898_ (_18538_, _18537_, _18533_);
  and _69899_ (_18539_, _18518_, _12239_);
  or _69900_ (_18540_, _18519_, _06840_);
  or _69901_ (_18541_, _18540_, _18539_);
  and _69902_ (_18543_, _18541_, _18538_);
  and _69903_ (_18544_, _18543_, _03710_);
  nor _69904_ (_18545_, _12256_, _09059_);
  nor _69905_ (_18546_, _18519_, _18545_);
  nor _69906_ (_18547_, _18546_, _03710_);
  or _69907_ (_18548_, _18547_, _07390_);
  nor _69908_ (_18549_, _18548_, _18544_);
  and _69909_ (_18550_, _18526_, _07390_);
  or _69910_ (_18551_, _18550_, _04481_);
  nor _69911_ (_18552_, _18551_, _18549_);
  or _69912_ (_18554_, _18552_, _18504_);
  and _69913_ (_18555_, _18554_, _03589_);
  nor _69914_ (_18556_, _12313_, _09021_);
  nor _69915_ (_18557_, _18556_, _18501_);
  nor _69916_ (_18558_, _18557_, _03589_);
  nor _69917_ (_18559_, _18558_, _18555_);
  nor _69918_ (_18560_, _18559_, _08828_);
  not _69919_ (_18561_, _18505_);
  nor _69920_ (_18562_, _12327_, _09021_);
  nor _69921_ (_18563_, _18562_, _07766_);
  and _69922_ (_18565_, _05229_, _04303_);
  nor _69923_ (_18566_, _18565_, _05886_);
  or _69924_ (_18567_, _18566_, _18563_);
  and _69925_ (_18568_, _18567_, _18561_);
  nor _69926_ (_18569_, _18568_, _18560_);
  nor _69927_ (_18570_, _18569_, _03780_);
  nor _69928_ (_18571_, _12333_, _09021_);
  nor _69929_ (_18572_, _18571_, _07778_);
  and _69930_ (_18573_, _18572_, _18561_);
  nor _69931_ (_18574_, _18573_, _18570_);
  nor _69932_ (_18576_, _18574_, _03622_);
  nor _69933_ (_18577_, _12207_, _09021_);
  nor _69934_ (_18578_, _18577_, _07777_);
  and _69935_ (_18579_, _18578_, _18561_);
  nor _69936_ (_18580_, _18579_, _18576_);
  nor _69937_ (_18581_, _18580_, _03790_);
  nor _69938_ (_18582_, _18501_, _05618_);
  nor _69939_ (_18583_, _18582_, _06828_);
  and _69940_ (_18584_, _18583_, _18507_);
  nor _69941_ (_18585_, _18584_, _18581_);
  or _69942_ (_18587_, _18585_, _18499_);
  and _69943_ (_18588_, _18565_, _05617_);
  nor _69944_ (_18589_, _18588_, _07795_);
  and _69945_ (_18590_, _18589_, _18561_);
  and _69946_ (_18591_, _18506_, _05617_);
  or _69947_ (_18592_, _18505_, _07793_);
  nor _69948_ (_18593_, _18592_, _18591_);
  or _69949_ (_18594_, _18593_, _03815_);
  nor _69950_ (_18595_, _18594_, _18590_);
  and _69951_ (_18596_, _18595_, _18587_);
  nor _69952_ (_18598_, _18514_, _04246_);
  or _69953_ (_18599_, _18598_, _03453_);
  nor _69954_ (_18600_, _18599_, _18596_);
  nor _69955_ (_18601_, _18535_, _03823_);
  or _69956_ (_18602_, _18601_, _03447_);
  nor _69957_ (_18603_, _18602_, _18600_);
  or _69958_ (_18604_, _18501_, _03514_);
  nor _69959_ (_18605_, _18604_, _18513_);
  nor _69960_ (_18606_, _18605_, _18603_);
  or _69961_ (_18607_, _18606_, _43004_);
  or _69962_ (_18609_, _43000_, \oc8051_golden_model_1.IE [1]);
  and _69963_ (_18610_, _18609_, _41806_);
  and _69964_ (_43517_, _18610_, _18607_);
  not _69965_ (_18611_, \oc8051_golden_model_1.IE [2]);
  nor _69966_ (_18612_, _05229_, _18611_);
  and _69967_ (_18613_, _05229_, _06332_);
  nor _69968_ (_18614_, _18613_, _18612_);
  and _69969_ (_18615_, _18614_, _03601_);
  nor _69970_ (_18616_, _09021_, _04875_);
  nor _69971_ (_18617_, _18616_, _18612_);
  and _69972_ (_18619_, _18617_, _07390_);
  and _69973_ (_18620_, _05229_, \oc8051_golden_model_1.ACC [2]);
  nor _69974_ (_18621_, _18620_, _18612_);
  nor _69975_ (_18622_, _18621_, _09029_);
  nor _69976_ (_18623_, _04409_, _18611_);
  or _69977_ (_18624_, _18623_, _18622_);
  and _69978_ (_18625_, _18624_, _04081_);
  nor _69979_ (_18626_, _12416_, _09021_);
  nor _69980_ (_18627_, _18626_, _18612_);
  nor _69981_ (_18628_, _18627_, _04081_);
  or _69982_ (_18630_, _18628_, _18625_);
  and _69983_ (_18631_, _18630_, _04055_);
  nor _69984_ (_18632_, _05924_, _18611_);
  and _69985_ (_18633_, _12411_, _05924_);
  nor _69986_ (_18634_, _18633_, _18632_);
  nor _69987_ (_18635_, _18634_, _04055_);
  or _69988_ (_18636_, _18635_, _18631_);
  and _69989_ (_18637_, _18636_, _03996_);
  nor _69990_ (_18638_, _18617_, _03996_);
  or _69991_ (_18639_, _18638_, _18637_);
  and _69992_ (_18641_, _18639_, _03737_);
  nor _69993_ (_18642_, _18621_, _03737_);
  or _69994_ (_18643_, _18642_, _18641_);
  and _69995_ (_18644_, _18643_, _03736_);
  and _69996_ (_18645_, _12409_, _05924_);
  nor _69997_ (_18646_, _18645_, _18632_);
  nor _69998_ (_18647_, _18646_, _03736_);
  or _69999_ (_18648_, _18647_, _03719_);
  or _70000_ (_18649_, _18648_, _18644_);
  and _70001_ (_18650_, _18633_, _12443_);
  or _70002_ (_18652_, _18632_, _06840_);
  or _70003_ (_18653_, _18652_, _18650_);
  and _70004_ (_18654_, _18653_, _03710_);
  and _70005_ (_18655_, _18654_, _18649_);
  nor _70006_ (_18656_, _12461_, _09059_);
  nor _70007_ (_18657_, _18656_, _18632_);
  nor _70008_ (_18658_, _18657_, _03710_);
  nor _70009_ (_18659_, _18658_, _07390_);
  not _70010_ (_18660_, _18659_);
  nor _70011_ (_18661_, _18660_, _18655_);
  nor _70012_ (_18663_, _18661_, _18619_);
  nor _70013_ (_18664_, _18663_, _04481_);
  and _70014_ (_18665_, _06637_, _05229_);
  nor _70015_ (_18666_, _18612_, _07400_);
  not _70016_ (_18667_, _18666_);
  nor _70017_ (_18668_, _18667_, _18665_);
  or _70018_ (_18669_, _18668_, _03222_);
  nor _70019_ (_18670_, _18669_, _18664_);
  nor _70020_ (_18671_, _12519_, _09021_);
  nor _70021_ (_18672_, _18612_, _18671_);
  nor _70022_ (_18674_, _18672_, _03589_);
  or _70023_ (_18675_, _18674_, _03601_);
  nor _70024_ (_18676_, _18675_, _18670_);
  nor _70025_ (_18677_, _18676_, _18615_);
  or _70026_ (_18678_, _18677_, _03600_);
  and _70027_ (_18679_, _12533_, _05229_);
  or _70028_ (_18680_, _18679_, _18612_);
  or _70029_ (_18681_, _18680_, _07766_);
  and _70030_ (_18682_, _18681_, _07778_);
  and _70031_ (_18683_, _18682_, _18678_);
  and _70032_ (_18685_, _12539_, _05229_);
  nor _70033_ (_18686_, _18685_, _18612_);
  nor _70034_ (_18687_, _18686_, _07778_);
  nor _70035_ (_18688_, _18687_, _18683_);
  nor _70036_ (_18689_, _18688_, _03622_);
  nor _70037_ (_18690_, _18612_, _05718_);
  not _70038_ (_18691_, _18690_);
  nor _70039_ (_18692_, _18614_, _07777_);
  and _70040_ (_18693_, _18692_, _18691_);
  nor _70041_ (_18694_, _18693_, _18689_);
  nor _70042_ (_18696_, _18694_, _03790_);
  nor _70043_ (_18697_, _18621_, _06828_);
  and _70044_ (_18698_, _18697_, _18691_);
  or _70045_ (_18699_, _18698_, _18696_);
  and _70046_ (_18700_, _18699_, _07795_);
  nor _70047_ (_18701_, _12532_, _09021_);
  nor _70048_ (_18702_, _18701_, _18612_);
  nor _70049_ (_18703_, _18702_, _07795_);
  or _70050_ (_18704_, _18703_, _18700_);
  and _70051_ (_18705_, _18704_, _07793_);
  nor _70052_ (_18707_, _12538_, _09021_);
  nor _70053_ (_18708_, _18707_, _18612_);
  nor _70054_ (_18709_, _18708_, _07793_);
  or _70055_ (_18710_, _18709_, _18705_);
  and _70056_ (_18711_, _18710_, _04246_);
  nor _70057_ (_18712_, _18627_, _04246_);
  or _70058_ (_18713_, _18712_, _18711_);
  and _70059_ (_18714_, _18713_, _03823_);
  nor _70060_ (_18715_, _18646_, _03823_);
  or _70061_ (_18716_, _18715_, _18714_);
  and _70062_ (_18718_, _18716_, _03514_);
  and _70063_ (_18719_, _12592_, _05229_);
  nor _70064_ (_18720_, _18719_, _18612_);
  nor _70065_ (_18721_, _18720_, _03514_);
  or _70066_ (_18722_, _18721_, _18718_);
  or _70067_ (_18723_, _18722_, _43004_);
  or _70068_ (_18724_, _43000_, \oc8051_golden_model_1.IE [2]);
  and _70069_ (_18725_, _18724_, _41806_);
  and _70070_ (_43518_, _18725_, _18723_);
  not _70071_ (_18726_, \oc8051_golden_model_1.IE [3]);
  nor _70072_ (_18728_, _05229_, _18726_);
  and _70073_ (_18729_, _05229_, _06276_);
  nor _70074_ (_18730_, _18729_, _18728_);
  and _70075_ (_18731_, _18730_, _03601_);
  nor _70076_ (_18732_, _09021_, _05005_);
  nor _70077_ (_18733_, _18732_, _18728_);
  and _70078_ (_18734_, _18733_, _07390_);
  and _70079_ (_18735_, _05229_, \oc8051_golden_model_1.ACC [3]);
  nor _70080_ (_18736_, _18735_, _18728_);
  nor _70081_ (_18737_, _18736_, _09029_);
  nor _70082_ (_18739_, _04409_, _18726_);
  or _70083_ (_18740_, _18739_, _18737_);
  and _70084_ (_18741_, _18740_, _04081_);
  nor _70085_ (_18742_, _12627_, _09021_);
  nor _70086_ (_18743_, _18742_, _18728_);
  nor _70087_ (_18744_, _18743_, _04081_);
  or _70088_ (_18745_, _18744_, _18741_);
  and _70089_ (_18746_, _18745_, _04055_);
  nor _70090_ (_18747_, _05924_, _18726_);
  and _70091_ (_18748_, _12631_, _05924_);
  nor _70092_ (_18750_, _18748_, _18747_);
  nor _70093_ (_18751_, _18750_, _04055_);
  or _70094_ (_18752_, _18751_, _03723_);
  or _70095_ (_18753_, _18752_, _18746_);
  nand _70096_ (_18754_, _18733_, _03723_);
  and _70097_ (_18755_, _18754_, _18753_);
  and _70098_ (_18756_, _18755_, _03737_);
  nor _70099_ (_18757_, _18736_, _03737_);
  or _70100_ (_18758_, _18757_, _18756_);
  and _70101_ (_18759_, _18758_, _03736_);
  and _70102_ (_18761_, _12641_, _05924_);
  nor _70103_ (_18762_, _18761_, _18747_);
  nor _70104_ (_18763_, _18762_, _03736_);
  or _70105_ (_18764_, _18763_, _03719_);
  or _70106_ (_18765_, _18764_, _18759_);
  nor _70107_ (_18766_, _18747_, _12648_);
  nor _70108_ (_18767_, _18766_, _18750_);
  or _70109_ (_18768_, _18767_, _06840_);
  and _70110_ (_18769_, _18768_, _03710_);
  and _70111_ (_18770_, _18769_, _18765_);
  nor _70112_ (_18772_, _12612_, _09059_);
  nor _70113_ (_18773_, _18772_, _18747_);
  nor _70114_ (_18774_, _18773_, _03710_);
  nor _70115_ (_18775_, _18774_, _07390_);
  not _70116_ (_18776_, _18775_);
  nor _70117_ (_18777_, _18776_, _18770_);
  nor _70118_ (_18778_, _18777_, _18734_);
  nor _70119_ (_18779_, _18778_, _04481_);
  and _70120_ (_18780_, _06592_, _05229_);
  nor _70121_ (_18781_, _18728_, _07400_);
  not _70122_ (_18783_, _18781_);
  nor _70123_ (_18784_, _18783_, _18780_);
  or _70124_ (_18785_, _18784_, _03222_);
  nor _70125_ (_18786_, _18785_, _18779_);
  nor _70126_ (_18787_, _12718_, _09021_);
  nor _70127_ (_18788_, _18728_, _18787_);
  nor _70128_ (_18789_, _18788_, _03589_);
  or _70129_ (_18790_, _18789_, _03601_);
  nor _70130_ (_18791_, _18790_, _18786_);
  nor _70131_ (_18792_, _18791_, _18731_);
  or _70132_ (_18794_, _18792_, _03600_);
  and _70133_ (_18795_, _12733_, _05229_);
  or _70134_ (_18796_, _18795_, _18728_);
  or _70135_ (_18797_, _18796_, _07766_);
  and _70136_ (_18798_, _18797_, _07778_);
  and _70137_ (_18799_, _18798_, _18794_);
  and _70138_ (_18800_, _12739_, _05229_);
  nor _70139_ (_18801_, _18800_, _18728_);
  nor _70140_ (_18802_, _18801_, _07778_);
  nor _70141_ (_18803_, _18802_, _18799_);
  nor _70142_ (_18805_, _18803_, _03622_);
  nor _70143_ (_18806_, _18728_, _05567_);
  not _70144_ (_18807_, _18806_);
  nor _70145_ (_18808_, _18730_, _07777_);
  and _70146_ (_18809_, _18808_, _18807_);
  nor _70147_ (_18810_, _18809_, _18805_);
  nor _70148_ (_18811_, _18810_, _03790_);
  nor _70149_ (_18812_, _18736_, _06828_);
  and _70150_ (_18813_, _18812_, _18807_);
  nor _70151_ (_18814_, _18813_, _03624_);
  not _70152_ (_18816_, _18814_);
  nor _70153_ (_18817_, _18816_, _18811_);
  nor _70154_ (_18818_, _12732_, _09021_);
  or _70155_ (_18819_, _18728_, _07795_);
  nor _70156_ (_18820_, _18819_, _18818_);
  or _70157_ (_18821_, _18820_, _03785_);
  nor _70158_ (_18822_, _18821_, _18817_);
  nor _70159_ (_18823_, _12738_, _09021_);
  nor _70160_ (_18824_, _18823_, _18728_);
  nor _70161_ (_18825_, _18824_, _07793_);
  or _70162_ (_18827_, _18825_, _18822_);
  and _70163_ (_18828_, _18827_, _04246_);
  nor _70164_ (_18829_, _18743_, _04246_);
  or _70165_ (_18830_, _18829_, _18828_);
  and _70166_ (_18831_, _18830_, _03823_);
  nor _70167_ (_18832_, _18762_, _03823_);
  or _70168_ (_18833_, _18832_, _18831_);
  and _70169_ (_18834_, _18833_, _03514_);
  and _70170_ (_18835_, _12794_, _05229_);
  nor _70171_ (_18836_, _18835_, _18728_);
  nor _70172_ (_18838_, _18836_, _03514_);
  or _70173_ (_18839_, _18838_, _18834_);
  or _70174_ (_18840_, _18839_, _43004_);
  or _70175_ (_18841_, _43000_, \oc8051_golden_model_1.IE [3]);
  and _70176_ (_18842_, _18841_, _41806_);
  and _70177_ (_43519_, _18842_, _18840_);
  not _70178_ (_18843_, \oc8051_golden_model_1.IE [4]);
  nor _70179_ (_18844_, _05229_, _18843_);
  nor _70180_ (_18845_, _05777_, _09021_);
  nor _70181_ (_18846_, _18845_, _18844_);
  and _70182_ (_18848_, _18846_, _07390_);
  nor _70183_ (_18849_, _05924_, _18843_);
  and _70184_ (_18850_, _12827_, _05924_);
  nor _70185_ (_18851_, _18850_, _18849_);
  nor _70186_ (_18852_, _18851_, _03736_);
  and _70187_ (_18853_, _05229_, \oc8051_golden_model_1.ACC [4]);
  nor _70188_ (_18854_, _18853_, _18844_);
  nor _70189_ (_18855_, _18854_, _09029_);
  nor _70190_ (_18856_, _04409_, _18843_);
  or _70191_ (_18857_, _18856_, _18855_);
  and _70192_ (_18859_, _18857_, _04081_);
  nor _70193_ (_18860_, _12841_, _09021_);
  nor _70194_ (_18861_, _18860_, _18844_);
  nor _70195_ (_18862_, _18861_, _04081_);
  or _70196_ (_18863_, _18862_, _18859_);
  and _70197_ (_18864_, _18863_, _04055_);
  and _70198_ (_18865_, _12845_, _05924_);
  nor _70199_ (_18866_, _18865_, _18849_);
  nor _70200_ (_18867_, _18866_, _04055_);
  or _70201_ (_18868_, _18867_, _03723_);
  or _70202_ (_18870_, _18868_, _18864_);
  nand _70203_ (_18871_, _18846_, _03723_);
  and _70204_ (_18872_, _18871_, _18870_);
  and _70205_ (_18873_, _18872_, _03737_);
  nor _70206_ (_18874_, _18854_, _03737_);
  or _70207_ (_18875_, _18874_, _18873_);
  and _70208_ (_18876_, _18875_, _03736_);
  nor _70209_ (_18877_, _18876_, _18852_);
  nor _70210_ (_18878_, _18877_, _03719_);
  and _70211_ (_18879_, _12861_, _05924_);
  nor _70212_ (_18881_, _18879_, _18849_);
  nor _70213_ (_18882_, _18881_, _06840_);
  nor _70214_ (_18883_, _18882_, _18878_);
  nor _70215_ (_18884_, _18883_, _03505_);
  nor _70216_ (_18885_, _12825_, _09059_);
  nor _70217_ (_18886_, _18885_, _18849_);
  nor _70218_ (_18887_, _18886_, _03710_);
  nor _70219_ (_18888_, _18887_, _07390_);
  not _70220_ (_18889_, _18888_);
  nor _70221_ (_18890_, _18889_, _18884_);
  nor _70222_ (_18892_, _18890_, _18848_);
  nor _70223_ (_18893_, _18892_, _04481_);
  and _70224_ (_18894_, _06730_, _05229_);
  nor _70225_ (_18895_, _18844_, _07400_);
  not _70226_ (_18896_, _18895_);
  nor _70227_ (_18897_, _18896_, _18894_);
  nor _70228_ (_18898_, _18897_, _03222_);
  not _70229_ (_18899_, _18898_);
  nor _70230_ (_18900_, _18899_, _18893_);
  nor _70231_ (_18901_, _12933_, _09021_);
  nor _70232_ (_18903_, _18901_, _18844_);
  nor _70233_ (_18904_, _18903_, _03589_);
  or _70234_ (_18905_, _18904_, _08828_);
  or _70235_ (_18906_, _18905_, _18900_);
  and _70236_ (_18907_, _12821_, _05229_);
  or _70237_ (_18908_, _18844_, _07766_);
  or _70238_ (_18909_, _18908_, _18907_);
  and _70239_ (_18910_, _06298_, _05229_);
  nor _70240_ (_18911_, _18910_, _18844_);
  and _70241_ (_18912_, _18911_, _03601_);
  nor _70242_ (_18914_, _18912_, _03780_);
  and _70243_ (_18915_, _18914_, _18909_);
  and _70244_ (_18916_, _18915_, _18906_);
  and _70245_ (_18917_, _12817_, _05229_);
  nor _70246_ (_18918_, _18917_, _18844_);
  nor _70247_ (_18919_, _18918_, _07778_);
  nor _70248_ (_18920_, _18919_, _18916_);
  nor _70249_ (_18921_, _18920_, _03622_);
  nor _70250_ (_18922_, _18844_, _05825_);
  not _70251_ (_18923_, _18922_);
  nor _70252_ (_18925_, _18911_, _07777_);
  and _70253_ (_18926_, _18925_, _18923_);
  nor _70254_ (_18927_, _18926_, _18921_);
  nor _70255_ (_18928_, _18927_, _03790_);
  nor _70256_ (_18929_, _18854_, _06828_);
  and _70257_ (_18930_, _18929_, _18923_);
  or _70258_ (_18931_, _18930_, _18928_);
  and _70259_ (_18932_, _18931_, _07795_);
  nor _70260_ (_18933_, _12819_, _09021_);
  nor _70261_ (_18934_, _18933_, _18844_);
  nor _70262_ (_18936_, _18934_, _07795_);
  or _70263_ (_18937_, _18936_, _18932_);
  and _70264_ (_18938_, _18937_, _07793_);
  nor _70265_ (_18939_, _12816_, _09021_);
  nor _70266_ (_18940_, _18939_, _18844_);
  nor _70267_ (_18941_, _18940_, _07793_);
  or _70268_ (_18942_, _18941_, _18938_);
  and _70269_ (_18943_, _18942_, _04246_);
  nor _70270_ (_18944_, _18861_, _04246_);
  or _70271_ (_18945_, _18944_, _18943_);
  and _70272_ (_18947_, _18945_, _03823_);
  nor _70273_ (_18948_, _18851_, _03823_);
  or _70274_ (_18949_, _18948_, _18947_);
  and _70275_ (_18950_, _18949_, _03514_);
  and _70276_ (_18951_, _13003_, _05229_);
  nor _70277_ (_18952_, _18951_, _18844_);
  nor _70278_ (_18953_, _18952_, _03514_);
  or _70279_ (_18954_, _18953_, _18950_);
  or _70280_ (_18955_, _18954_, _43004_);
  or _70281_ (_18956_, _43000_, \oc8051_golden_model_1.IE [4]);
  and _70282_ (_18958_, _18956_, _41806_);
  and _70283_ (_43520_, _18958_, _18955_);
  not _70284_ (_18959_, \oc8051_golden_model_1.IE [5]);
  nor _70285_ (_18960_, _05229_, _18959_);
  and _70286_ (_18961_, _06684_, _05229_);
  or _70287_ (_18962_, _18961_, _18960_);
  and _70288_ (_18963_, _18962_, _04481_);
  and _70289_ (_18964_, _05229_, \oc8051_golden_model_1.ACC [5]);
  nor _70290_ (_18965_, _18964_, _18960_);
  nor _70291_ (_18966_, _18965_, _09029_);
  nor _70292_ (_18968_, _04409_, _18959_);
  or _70293_ (_18969_, _18968_, _18966_);
  and _70294_ (_18970_, _18969_, _04081_);
  nor _70295_ (_18971_, _13014_, _09021_);
  nor _70296_ (_18972_, _18971_, _18960_);
  nor _70297_ (_18973_, _18972_, _04081_);
  or _70298_ (_18974_, _18973_, _18970_);
  and _70299_ (_18975_, _18974_, _04055_);
  nor _70300_ (_18976_, _05924_, _18959_);
  and _70301_ (_18977_, _13037_, _05924_);
  nor _70302_ (_18979_, _18977_, _18976_);
  nor _70303_ (_18980_, _18979_, _04055_);
  or _70304_ (_18981_, _18980_, _03723_);
  or _70305_ (_18982_, _18981_, _18975_);
  nor _70306_ (_18983_, _05469_, _09021_);
  nor _70307_ (_18984_, _18983_, _18960_);
  nand _70308_ (_18985_, _18984_, _03723_);
  and _70309_ (_18986_, _18985_, _18982_);
  and _70310_ (_18987_, _18986_, _03737_);
  nor _70311_ (_18988_, _18965_, _03737_);
  or _70312_ (_18990_, _18988_, _18987_);
  and _70313_ (_18991_, _18990_, _03736_);
  and _70314_ (_18992_, _13047_, _05924_);
  nor _70315_ (_18993_, _18992_, _18976_);
  nor _70316_ (_18994_, _18993_, _03736_);
  or _70317_ (_18995_, _18994_, _03719_);
  or _70318_ (_18996_, _18995_, _18991_);
  nor _70319_ (_18997_, _18976_, _13054_);
  nor _70320_ (_18998_, _18997_, _18979_);
  or _70321_ (_18999_, _18998_, _06840_);
  and _70322_ (_19001_, _18999_, _03710_);
  and _70323_ (_19002_, _19001_, _18996_);
  nor _70324_ (_19003_, _13020_, _09059_);
  nor _70325_ (_19004_, _19003_, _18976_);
  nor _70326_ (_19005_, _19004_, _03710_);
  nor _70327_ (_19006_, _19005_, _07390_);
  not _70328_ (_19007_, _19006_);
  nor _70329_ (_19008_, _19007_, _19002_);
  and _70330_ (_19009_, _18984_, _07390_);
  or _70331_ (_19010_, _19009_, _04481_);
  nor _70332_ (_19012_, _19010_, _19008_);
  or _70333_ (_19013_, _19012_, _18963_);
  and _70334_ (_19014_, _19013_, _03589_);
  nor _70335_ (_19015_, _13127_, _09021_);
  nor _70336_ (_19016_, _19015_, _18960_);
  nor _70337_ (_19017_, _19016_, _03589_);
  or _70338_ (_19018_, _19017_, _08828_);
  or _70339_ (_19019_, _19018_, _19014_);
  and _70340_ (_19020_, _13141_, _05229_);
  or _70341_ (_19021_, _18960_, _07766_);
  or _70342_ (_19023_, _19021_, _19020_);
  and _70343_ (_19024_, _06306_, _05229_);
  nor _70344_ (_19025_, _19024_, _18960_);
  and _70345_ (_19026_, _19025_, _03601_);
  nor _70346_ (_19027_, _19026_, _03780_);
  and _70347_ (_19028_, _19027_, _19023_);
  and _70348_ (_19029_, _19028_, _19019_);
  and _70349_ (_19030_, _13147_, _05229_);
  nor _70350_ (_19031_, _19030_, _18960_);
  nor _70351_ (_19032_, _19031_, _07778_);
  nor _70352_ (_19034_, _19032_, _19029_);
  nor _70353_ (_19035_, _19034_, _03622_);
  nor _70354_ (_19036_, _18960_, _05518_);
  not _70355_ (_19037_, _19036_);
  nor _70356_ (_19038_, _19025_, _07777_);
  and _70357_ (_19039_, _19038_, _19037_);
  nor _70358_ (_19040_, _19039_, _19035_);
  nor _70359_ (_19041_, _19040_, _03790_);
  nor _70360_ (_19042_, _18965_, _06828_);
  and _70361_ (_19043_, _19042_, _19037_);
  or _70362_ (_19045_, _19043_, _19041_);
  and _70363_ (_19046_, _19045_, _07795_);
  nor _70364_ (_19047_, _13140_, _09021_);
  nor _70365_ (_19048_, _19047_, _18960_);
  nor _70366_ (_19049_, _19048_, _07795_);
  or _70367_ (_19050_, _19049_, _19046_);
  and _70368_ (_19051_, _19050_, _07793_);
  nor _70369_ (_19052_, _13146_, _09021_);
  nor _70370_ (_19053_, _19052_, _18960_);
  nor _70371_ (_19054_, _19053_, _07793_);
  or _70372_ (_19056_, _19054_, _19051_);
  and _70373_ (_19057_, _19056_, _04246_);
  nor _70374_ (_19058_, _18972_, _04246_);
  or _70375_ (_19059_, _19058_, _19057_);
  and _70376_ (_19060_, _19059_, _03823_);
  nor _70377_ (_19061_, _18993_, _03823_);
  or _70378_ (_19062_, _19061_, _19060_);
  and _70379_ (_19063_, _19062_, _03514_);
  and _70380_ (_19064_, _13199_, _05229_);
  nor _70381_ (_19065_, _19064_, _18960_);
  nor _70382_ (_19067_, _19065_, _03514_);
  or _70383_ (_19068_, _19067_, _19063_);
  or _70384_ (_19069_, _19068_, _43004_);
  or _70385_ (_19070_, _43000_, \oc8051_golden_model_1.IE [5]);
  and _70386_ (_19071_, _19070_, _41806_);
  and _70387_ (_43521_, _19071_, _19069_);
  not _70388_ (_19072_, \oc8051_golden_model_1.IE [6]);
  nor _70389_ (_19073_, _05229_, _19072_);
  and _70390_ (_19074_, _06455_, _05229_);
  or _70391_ (_19075_, _19074_, _19073_);
  and _70392_ (_19077_, _19075_, _04481_);
  and _70393_ (_19078_, _05229_, \oc8051_golden_model_1.ACC [6]);
  nor _70394_ (_19079_, _19078_, _19073_);
  nor _70395_ (_19080_, _19079_, _09029_);
  nor _70396_ (_19081_, _04409_, _19072_);
  or _70397_ (_19082_, _19081_, _19080_);
  and _70398_ (_19083_, _19082_, _04081_);
  nor _70399_ (_19084_, _13242_, _09021_);
  nor _70400_ (_19085_, _19084_, _19073_);
  nor _70401_ (_19086_, _19085_, _04081_);
  or _70402_ (_19088_, _19086_, _19083_);
  and _70403_ (_19089_, _19088_, _04055_);
  nor _70404_ (_19090_, _05924_, _19072_);
  and _70405_ (_19091_, _13229_, _05924_);
  nor _70406_ (_19092_, _19091_, _19090_);
  nor _70407_ (_19093_, _19092_, _04055_);
  or _70408_ (_19094_, _19093_, _03723_);
  or _70409_ (_19095_, _19094_, _19089_);
  nor _70410_ (_19096_, _05363_, _09021_);
  nor _70411_ (_19097_, _19096_, _19073_);
  nand _70412_ (_19099_, _19097_, _03723_);
  and _70413_ (_19100_, _19099_, _19095_);
  and _70414_ (_19101_, _19100_, _03737_);
  nor _70415_ (_19102_, _19079_, _03737_);
  or _70416_ (_19103_, _19102_, _19101_);
  and _70417_ (_19104_, _19103_, _03736_);
  and _70418_ (_19105_, _13253_, _05924_);
  nor _70419_ (_19106_, _19105_, _19090_);
  nor _70420_ (_19107_, _19106_, _03736_);
  or _70421_ (_19108_, _19107_, _19104_);
  and _70422_ (_19110_, _19108_, _06840_);
  nor _70423_ (_19111_, _19090_, _13260_);
  nor _70424_ (_19112_, _19111_, _19092_);
  and _70425_ (_19113_, _19112_, _03719_);
  or _70426_ (_19114_, _19113_, _19110_);
  and _70427_ (_19115_, _19114_, _03710_);
  nor _70428_ (_19116_, _13226_, _09059_);
  nor _70429_ (_19117_, _19116_, _19090_);
  nor _70430_ (_19118_, _19117_, _03710_);
  nor _70431_ (_19119_, _19118_, _07390_);
  not _70432_ (_19121_, _19119_);
  nor _70433_ (_19122_, _19121_, _19115_);
  and _70434_ (_19123_, _19097_, _07390_);
  or _70435_ (_19124_, _19123_, _04481_);
  nor _70436_ (_19125_, _19124_, _19122_);
  or _70437_ (_19126_, _19125_, _19077_);
  and _70438_ (_19127_, _19126_, _03589_);
  nor _70439_ (_19128_, _13332_, _09021_);
  nor _70440_ (_19129_, _19128_, _19073_);
  nor _70441_ (_19130_, _19129_, _03589_);
  or _70442_ (_19132_, _19130_, _08828_);
  or _70443_ (_19133_, _19132_, _19127_);
  and _70444_ (_19134_, _13347_, _05229_);
  or _70445_ (_19135_, _19073_, _07766_);
  or _70446_ (_19136_, _19135_, _19134_);
  and _70447_ (_19137_, _13339_, _05229_);
  nor _70448_ (_19138_, _19137_, _19073_);
  and _70449_ (_19139_, _19138_, _03601_);
  nor _70450_ (_19140_, _19139_, _03780_);
  and _70451_ (_19141_, _19140_, _19136_);
  and _70452_ (_19143_, _19141_, _19133_);
  and _70453_ (_19144_, _13353_, _05229_);
  nor _70454_ (_19145_, _19144_, _19073_);
  nor _70455_ (_19146_, _19145_, _07778_);
  nor _70456_ (_19147_, _19146_, _19143_);
  nor _70457_ (_19148_, _19147_, _03622_);
  nor _70458_ (_19149_, _19073_, _05412_);
  not _70459_ (_19150_, _19149_);
  nor _70460_ (_19151_, _19138_, _07777_);
  and _70461_ (_19152_, _19151_, _19150_);
  nor _70462_ (_19154_, _19152_, _19148_);
  nor _70463_ (_19155_, _19154_, _03790_);
  nor _70464_ (_19156_, _19079_, _06828_);
  and _70465_ (_19157_, _19156_, _19150_);
  nor _70466_ (_19158_, _19157_, _03624_);
  not _70467_ (_19159_, _19158_);
  nor _70468_ (_19160_, _19159_, _19155_);
  nor _70469_ (_19161_, _13346_, _09021_);
  or _70470_ (_19162_, _19073_, _07795_);
  nor _70471_ (_19163_, _19162_, _19161_);
  or _70472_ (_19165_, _19163_, _03785_);
  nor _70473_ (_19166_, _19165_, _19160_);
  nor _70474_ (_19167_, _13352_, _09021_);
  nor _70475_ (_19168_, _19167_, _19073_);
  nor _70476_ (_19169_, _19168_, _07793_);
  or _70477_ (_19170_, _19169_, _19166_);
  and _70478_ (_19171_, _19170_, _04246_);
  nor _70479_ (_19172_, _19085_, _04246_);
  or _70480_ (_19173_, _19172_, _19171_);
  and _70481_ (_19174_, _19173_, _03823_);
  nor _70482_ (_19176_, _19106_, _03823_);
  or _70483_ (_19177_, _19176_, _19174_);
  and _70484_ (_19178_, _19177_, _03514_);
  and _70485_ (_19179_, _13402_, _05229_);
  nor _70486_ (_19180_, _19179_, _19073_);
  nor _70487_ (_19181_, _19180_, _03514_);
  or _70488_ (_19182_, _19181_, _19178_);
  or _70489_ (_19183_, _19182_, _43004_);
  or _70490_ (_19184_, _43000_, \oc8051_golden_model_1.IE [6]);
  and _70491_ (_19185_, _19184_, _41806_);
  and _70492_ (_43522_, _19185_, _19183_);
  not _70493_ (_19187_, \oc8051_golden_model_1.IP [0]);
  nor _70494_ (_19188_, _05251_, _19187_);
  and _70495_ (_19189_, _12128_, _05251_);
  nor _70496_ (_19190_, _19189_, _19188_);
  nor _70497_ (_19191_, _19190_, _07778_);
  and _70498_ (_19192_, _05251_, _06274_);
  nor _70499_ (_19193_, _19192_, _19188_);
  and _70500_ (_19194_, _19193_, _03601_);
  and _70501_ (_19195_, _05251_, _04620_);
  nor _70502_ (_19197_, _19195_, _19188_);
  and _70503_ (_19198_, _19197_, _07390_);
  nor _70504_ (_19199_, _05666_, _09129_);
  nor _70505_ (_19200_, _19199_, _19188_);
  nor _70506_ (_19201_, _19200_, _04081_);
  nor _70507_ (_19202_, _04409_, _19187_);
  and _70508_ (_19203_, _05251_, \oc8051_golden_model_1.ACC [0]);
  nor _70509_ (_19204_, _19203_, _19188_);
  nor _70510_ (_19205_, _19204_, _09029_);
  nor _70511_ (_19206_, _19205_, _19202_);
  nor _70512_ (_19208_, _19206_, _03610_);
  or _70513_ (_19209_, _19208_, _03715_);
  nor _70514_ (_19210_, _19209_, _19201_);
  and _70515_ (_19211_, _12021_, _05908_);
  nor _70516_ (_19212_, _05908_, _19187_);
  or _70517_ (_19213_, _19212_, _04055_);
  nor _70518_ (_19214_, _19213_, _19211_);
  or _70519_ (_19215_, _19214_, _03723_);
  nor _70520_ (_19216_, _19215_, _19210_);
  nor _70521_ (_19217_, _19197_, _03996_);
  or _70522_ (_19219_, _19217_, _19216_);
  and _70523_ (_19220_, _19219_, _03737_);
  nor _70524_ (_19221_, _19204_, _03737_);
  or _70525_ (_19222_, _19221_, _19220_);
  and _70526_ (_19223_, _19222_, _03736_);
  and _70527_ (_19224_, _19188_, _03714_);
  or _70528_ (_19225_, _19224_, _19223_);
  and _70529_ (_19226_, _19225_, _06840_);
  nor _70530_ (_19227_, _19200_, _06840_);
  or _70531_ (_19228_, _19227_, _19226_);
  and _70532_ (_19230_, _19228_, _03710_);
  nor _70533_ (_19231_, _12052_, _09166_);
  nor _70534_ (_19232_, _19231_, _19212_);
  nor _70535_ (_19233_, _19232_, _03710_);
  or _70536_ (_19234_, _19233_, _07390_);
  nor _70537_ (_19235_, _19234_, _19230_);
  nor _70538_ (_19236_, _19235_, _19198_);
  nor _70539_ (_19237_, _19236_, _04481_);
  and _70540_ (_19238_, _06546_, _05251_);
  nor _70541_ (_19239_, _19188_, _07400_);
  not _70542_ (_19241_, _19239_);
  nor _70543_ (_19242_, _19241_, _19238_);
  or _70544_ (_19243_, _19242_, _03222_);
  nor _70545_ (_19244_, _19243_, _19237_);
  nor _70546_ (_19245_, _12109_, _09129_);
  nor _70547_ (_19246_, _19245_, _19188_);
  nor _70548_ (_19247_, _19246_, _03589_);
  or _70549_ (_19248_, _19247_, _03601_);
  nor _70550_ (_19249_, _19248_, _19244_);
  nor _70551_ (_19250_, _19249_, _19194_);
  or _70552_ (_19252_, _19250_, _03600_);
  and _70553_ (_19253_, _12124_, _05251_);
  or _70554_ (_19254_, _19253_, _19188_);
  or _70555_ (_19255_, _19254_, _07766_);
  and _70556_ (_19256_, _19255_, _07778_);
  and _70557_ (_19257_, _19256_, _19252_);
  nor _70558_ (_19258_, _19257_, _19191_);
  nor _70559_ (_19259_, _19258_, _03622_);
  or _70560_ (_19260_, _19193_, _07777_);
  nor _70561_ (_19261_, _19260_, _19199_);
  nor _70562_ (_19263_, _19261_, _19259_);
  nor _70563_ (_19264_, _19263_, _03790_);
  and _70564_ (_19265_, _12005_, _05251_);
  or _70565_ (_19266_, _19265_, _19188_);
  and _70566_ (_19267_, _19266_, _03790_);
  or _70567_ (_19268_, _19267_, _19264_);
  and _70568_ (_19269_, _19268_, _07795_);
  nor _70569_ (_19270_, _12122_, _09129_);
  nor _70570_ (_19271_, _19270_, _19188_);
  nor _70571_ (_19272_, _19271_, _07795_);
  or _70572_ (_19274_, _19272_, _19269_);
  and _70573_ (_19275_, _19274_, _07793_);
  nor _70574_ (_19276_, _12003_, _09129_);
  nor _70575_ (_19277_, _19276_, _19188_);
  nor _70576_ (_19278_, _19277_, _07793_);
  or _70577_ (_19279_, _19278_, _19275_);
  and _70578_ (_19280_, _19279_, _04246_);
  nor _70579_ (_19281_, _19200_, _04246_);
  or _70580_ (_19282_, _19281_, _19280_);
  and _70581_ (_19283_, _19282_, _03823_);
  and _70582_ (_19285_, _19188_, _03453_);
  or _70583_ (_19286_, _19285_, _19283_);
  and _70584_ (_19287_, _19286_, _03514_);
  nor _70585_ (_19288_, _19200_, _03514_);
  or _70586_ (_19289_, _19288_, _19287_);
  or _70587_ (_19290_, _19289_, _43004_);
  or _70588_ (_19291_, _43000_, \oc8051_golden_model_1.IP [0]);
  and _70589_ (_19292_, _19291_, _41806_);
  and _70590_ (_43525_, _19292_, _19290_);
  not _70591_ (_19293_, \oc8051_golden_model_1.IP [1]);
  nor _70592_ (_19295_, _05251_, _19293_);
  and _70593_ (_19296_, _06501_, _05251_);
  or _70594_ (_19297_, _19296_, _19295_);
  and _70595_ (_19298_, _19297_, _04481_);
  nor _70596_ (_19299_, _05251_, \oc8051_golden_model_1.IP [1]);
  and _70597_ (_19300_, _05251_, _03274_);
  nor _70598_ (_19301_, _19300_, _19299_);
  and _70599_ (_19302_, _19301_, _04409_);
  nor _70600_ (_19303_, _04409_, _19293_);
  or _70601_ (_19304_, _19303_, _19302_);
  and _70602_ (_19306_, _19304_, _04081_);
  and _70603_ (_19307_, _12213_, _05251_);
  nor _70604_ (_19308_, _19307_, _19299_);
  and _70605_ (_19309_, _19308_, _03610_);
  or _70606_ (_19310_, _19309_, _19306_);
  and _70607_ (_19311_, _19310_, _04055_);
  and _70608_ (_19312_, _12224_, _05908_);
  nor _70609_ (_19313_, _05908_, _19293_);
  or _70610_ (_19314_, _19313_, _03723_);
  or _70611_ (_19315_, _19314_, _19312_);
  and _70612_ (_19317_, _19315_, _14265_);
  nor _70613_ (_19318_, _19317_, _19311_);
  and _70614_ (_19319_, _05251_, _06764_);
  nor _70615_ (_19320_, _19319_, _19295_);
  and _70616_ (_19321_, _19320_, _03723_);
  nor _70617_ (_19322_, _19321_, _19318_);
  and _70618_ (_19323_, _19322_, _03737_);
  and _70619_ (_19324_, _19301_, _03729_);
  or _70620_ (_19325_, _19324_, _19323_);
  and _70621_ (_19326_, _19325_, _03736_);
  and _70622_ (_19328_, _12211_, _05908_);
  nor _70623_ (_19329_, _19328_, _19313_);
  nor _70624_ (_19330_, _19329_, _03736_);
  or _70625_ (_19331_, _19330_, _19326_);
  and _70626_ (_19332_, _19331_, _06840_);
  and _70627_ (_19333_, _19312_, _12239_);
  or _70628_ (_19334_, _19333_, _19313_);
  and _70629_ (_19335_, _19334_, _03719_);
  or _70630_ (_19336_, _19335_, _19332_);
  and _70631_ (_19337_, _19336_, _03710_);
  nor _70632_ (_19339_, _12256_, _09166_);
  nor _70633_ (_19340_, _19313_, _19339_);
  nor _70634_ (_19341_, _19340_, _03710_);
  or _70635_ (_19342_, _19341_, _07390_);
  nor _70636_ (_19343_, _19342_, _19337_);
  and _70637_ (_19344_, _19320_, _07390_);
  or _70638_ (_19345_, _19344_, _04481_);
  nor _70639_ (_19346_, _19345_, _19343_);
  or _70640_ (_19347_, _19346_, _19298_);
  and _70641_ (_19348_, _19347_, _03589_);
  nor _70642_ (_19350_, _12313_, _09129_);
  nor _70643_ (_19351_, _19350_, _19295_);
  nor _70644_ (_19352_, _19351_, _03589_);
  nor _70645_ (_19353_, _19352_, _19348_);
  nor _70646_ (_19354_, _19353_, _08828_);
  nor _70647_ (_19355_, _12327_, _09129_);
  nor _70648_ (_19356_, _19355_, _07766_);
  and _70649_ (_19357_, _05251_, _04303_);
  nor _70650_ (_19358_, _19357_, _05886_);
  nor _70651_ (_19359_, _19358_, _19356_);
  nor _70652_ (_19361_, _19359_, _19299_);
  nor _70653_ (_19362_, _19361_, _19354_);
  nor _70654_ (_19363_, _19362_, _03780_);
  not _70655_ (_19364_, _19299_);
  nor _70656_ (_19365_, _12333_, _09129_);
  nor _70657_ (_19366_, _19365_, _07778_);
  and _70658_ (_19367_, _19366_, _19364_);
  nor _70659_ (_19368_, _19367_, _19363_);
  nor _70660_ (_19369_, _19368_, _03622_);
  nor _70661_ (_19370_, _12207_, _09129_);
  nor _70662_ (_19372_, _19370_, _07777_);
  and _70663_ (_19373_, _19372_, _19364_);
  nor _70664_ (_19374_, _19373_, _19369_);
  nor _70665_ (_19375_, _19374_, _03790_);
  nor _70666_ (_19376_, _19295_, _05618_);
  nor _70667_ (_19377_, _19376_, _06828_);
  and _70668_ (_19378_, _19377_, _19301_);
  nor _70669_ (_19379_, _19378_, _19375_);
  or _70670_ (_19380_, _19379_, _18499_);
  and _70671_ (_19381_, _19357_, _05617_);
  or _70672_ (_19383_, _19299_, _07795_);
  or _70673_ (_19384_, _19383_, _19381_);
  and _70674_ (_19385_, _19300_, _05617_);
  or _70675_ (_19386_, _19299_, _07793_);
  or _70676_ (_19387_, _19386_, _19385_);
  and _70677_ (_19388_, _19387_, _04246_);
  and _70678_ (_19389_, _19388_, _19384_);
  and _70679_ (_19390_, _19389_, _19380_);
  nor _70680_ (_19391_, _19308_, _04246_);
  or _70681_ (_19392_, _19391_, _03453_);
  nor _70682_ (_19394_, _19392_, _19390_);
  nor _70683_ (_19395_, _19329_, _03823_);
  or _70684_ (_19396_, _19395_, _03447_);
  nor _70685_ (_19397_, _19396_, _19394_);
  or _70686_ (_19398_, _19295_, _03514_);
  nor _70687_ (_19399_, _19398_, _19307_);
  nor _70688_ (_19400_, _19399_, _19397_);
  or _70689_ (_19401_, _19400_, _43004_);
  or _70690_ (_19402_, _43000_, \oc8051_golden_model_1.IP [1]);
  and _70691_ (_19403_, _19402_, _41806_);
  and _70692_ (_43526_, _19403_, _19401_);
  not _70693_ (_19405_, \oc8051_golden_model_1.IP [2]);
  nor _70694_ (_19406_, _05251_, _19405_);
  and _70695_ (_19407_, _05251_, _06332_);
  nor _70696_ (_19408_, _19407_, _19406_);
  and _70697_ (_19409_, _19408_, _03601_);
  nor _70698_ (_19410_, _09129_, _04875_);
  nor _70699_ (_19411_, _19410_, _19406_);
  and _70700_ (_19412_, _19411_, _07390_);
  and _70701_ (_19413_, _05251_, \oc8051_golden_model_1.ACC [2]);
  nor _70702_ (_19415_, _19413_, _19406_);
  nor _70703_ (_19416_, _19415_, _09029_);
  nor _70704_ (_19417_, _04409_, _19405_);
  or _70705_ (_19418_, _19417_, _19416_);
  and _70706_ (_19419_, _19418_, _04081_);
  nor _70707_ (_19420_, _12416_, _09129_);
  nor _70708_ (_19421_, _19420_, _19406_);
  nor _70709_ (_19422_, _19421_, _04081_);
  or _70710_ (_19423_, _19422_, _19419_);
  and _70711_ (_19424_, _19423_, _04055_);
  nor _70712_ (_19426_, _05908_, _19405_);
  and _70713_ (_19427_, _12411_, _05908_);
  nor _70714_ (_19428_, _19427_, _19426_);
  nor _70715_ (_19429_, _19428_, _04055_);
  or _70716_ (_19430_, _19429_, _19424_);
  and _70717_ (_19431_, _19430_, _03996_);
  nor _70718_ (_19432_, _19411_, _03996_);
  or _70719_ (_19433_, _19432_, _19431_);
  and _70720_ (_19434_, _19433_, _03737_);
  nor _70721_ (_19435_, _19415_, _03737_);
  or _70722_ (_19437_, _19435_, _19434_);
  and _70723_ (_19438_, _19437_, _03736_);
  and _70724_ (_19439_, _12409_, _05908_);
  nor _70725_ (_19440_, _19439_, _19426_);
  nor _70726_ (_19441_, _19440_, _03736_);
  or _70727_ (_19442_, _19441_, _03719_);
  or _70728_ (_19443_, _19442_, _19438_);
  and _70729_ (_19444_, _19427_, _12443_);
  or _70730_ (_19445_, _19426_, _06840_);
  or _70731_ (_19446_, _19445_, _19444_);
  and _70732_ (_19448_, _19446_, _03710_);
  and _70733_ (_19449_, _19448_, _19443_);
  nor _70734_ (_19450_, _12461_, _09166_);
  nor _70735_ (_19451_, _19450_, _19426_);
  nor _70736_ (_19452_, _19451_, _03710_);
  nor _70737_ (_19453_, _19452_, _07390_);
  not _70738_ (_19454_, _19453_);
  nor _70739_ (_19455_, _19454_, _19449_);
  nor _70740_ (_19456_, _19455_, _19412_);
  nor _70741_ (_19457_, _19456_, _04481_);
  and _70742_ (_19459_, _06637_, _05251_);
  nor _70743_ (_19460_, _19406_, _07400_);
  not _70744_ (_19461_, _19460_);
  nor _70745_ (_19462_, _19461_, _19459_);
  or _70746_ (_19463_, _19462_, _03222_);
  nor _70747_ (_19464_, _19463_, _19457_);
  nor _70748_ (_19465_, _12519_, _09129_);
  nor _70749_ (_19466_, _19406_, _19465_);
  nor _70750_ (_19467_, _19466_, _03589_);
  or _70751_ (_19468_, _19467_, _03601_);
  nor _70752_ (_19470_, _19468_, _19464_);
  nor _70753_ (_19471_, _19470_, _19409_);
  or _70754_ (_19472_, _19471_, _03600_);
  and _70755_ (_19473_, _12533_, _05251_);
  or _70756_ (_19474_, _19473_, _19406_);
  or _70757_ (_19475_, _19474_, _07766_);
  and _70758_ (_19476_, _19475_, _07778_);
  and _70759_ (_19477_, _19476_, _19472_);
  and _70760_ (_19478_, _12539_, _05251_);
  nor _70761_ (_19479_, _19478_, _19406_);
  nor _70762_ (_19481_, _19479_, _07778_);
  nor _70763_ (_19482_, _19481_, _19477_);
  nor _70764_ (_19483_, _19482_, _03622_);
  nor _70765_ (_19484_, _19406_, _05718_);
  not _70766_ (_19485_, _19484_);
  nor _70767_ (_19486_, _19408_, _07777_);
  and _70768_ (_19487_, _19486_, _19485_);
  nor _70769_ (_19488_, _19487_, _19483_);
  nor _70770_ (_19489_, _19488_, _03790_);
  nor _70771_ (_19490_, _19415_, _06828_);
  and _70772_ (_19492_, _19490_, _19485_);
  nor _70773_ (_19493_, _19492_, _03624_);
  not _70774_ (_19494_, _19493_);
  nor _70775_ (_19495_, _19494_, _19489_);
  nor _70776_ (_19496_, _12532_, _09129_);
  or _70777_ (_19497_, _19406_, _07795_);
  nor _70778_ (_19498_, _19497_, _19496_);
  or _70779_ (_19499_, _19498_, _03785_);
  nor _70780_ (_19500_, _19499_, _19495_);
  nor _70781_ (_19501_, _12538_, _09129_);
  nor _70782_ (_19503_, _19501_, _19406_);
  nor _70783_ (_19504_, _19503_, _07793_);
  or _70784_ (_19505_, _19504_, _19500_);
  and _70785_ (_19506_, _19505_, _04246_);
  nor _70786_ (_19507_, _19421_, _04246_);
  or _70787_ (_19508_, _19507_, _19506_);
  and _70788_ (_19509_, _19508_, _03823_);
  nor _70789_ (_19510_, _19440_, _03823_);
  or _70790_ (_19511_, _19510_, _19509_);
  and _70791_ (_19512_, _19511_, _03514_);
  and _70792_ (_19514_, _12592_, _05251_);
  nor _70793_ (_19515_, _19514_, _19406_);
  nor _70794_ (_19516_, _19515_, _03514_);
  or _70795_ (_19517_, _19516_, _19512_);
  or _70796_ (_19518_, _19517_, _43004_);
  or _70797_ (_19519_, _43000_, \oc8051_golden_model_1.IP [2]);
  and _70798_ (_19520_, _19519_, _41806_);
  and _70799_ (_43527_, _19520_, _19518_);
  not _70800_ (_19521_, \oc8051_golden_model_1.IP [3]);
  nor _70801_ (_19522_, _05251_, _19521_);
  and _70802_ (_19524_, _05251_, _06276_);
  nor _70803_ (_19525_, _19524_, _19522_);
  and _70804_ (_19526_, _19525_, _03601_);
  nor _70805_ (_19527_, _09129_, _05005_);
  nor _70806_ (_19528_, _19527_, _19522_);
  and _70807_ (_19529_, _19528_, _07390_);
  and _70808_ (_19530_, _05251_, \oc8051_golden_model_1.ACC [3]);
  nor _70809_ (_19531_, _19530_, _19522_);
  nor _70810_ (_19532_, _19531_, _09029_);
  nor _70811_ (_19533_, _04409_, _19521_);
  or _70812_ (_19535_, _19533_, _19532_);
  and _70813_ (_19536_, _19535_, _04081_);
  nor _70814_ (_19537_, _12627_, _09129_);
  nor _70815_ (_19538_, _19537_, _19522_);
  nor _70816_ (_19539_, _19538_, _04081_);
  or _70817_ (_19540_, _19539_, _19536_);
  and _70818_ (_19541_, _19540_, _04055_);
  nor _70819_ (_19542_, _05908_, _19521_);
  and _70820_ (_19543_, _12631_, _05908_);
  nor _70821_ (_19544_, _19543_, _19542_);
  nor _70822_ (_19546_, _19544_, _04055_);
  or _70823_ (_19547_, _19546_, _03723_);
  or _70824_ (_19548_, _19547_, _19541_);
  nand _70825_ (_19549_, _19528_, _03723_);
  and _70826_ (_19550_, _19549_, _19548_);
  and _70827_ (_19551_, _19550_, _03737_);
  nor _70828_ (_19552_, _19531_, _03737_);
  or _70829_ (_19553_, _19552_, _19551_);
  and _70830_ (_19554_, _19553_, _03736_);
  and _70831_ (_19555_, _12641_, _05908_);
  nor _70832_ (_19557_, _19555_, _19542_);
  nor _70833_ (_19558_, _19557_, _03736_);
  or _70834_ (_19559_, _19558_, _19554_);
  and _70835_ (_19560_, _19559_, _06840_);
  nor _70836_ (_19561_, _19542_, _12648_);
  nor _70837_ (_19562_, _19561_, _19544_);
  and _70838_ (_19563_, _19562_, _03719_);
  or _70839_ (_19564_, _19563_, _19560_);
  and _70840_ (_19565_, _19564_, _03710_);
  nor _70841_ (_19566_, _12612_, _09166_);
  nor _70842_ (_19568_, _19566_, _19542_);
  nor _70843_ (_19569_, _19568_, _03710_);
  nor _70844_ (_19570_, _19569_, _07390_);
  not _70845_ (_19571_, _19570_);
  nor _70846_ (_19572_, _19571_, _19565_);
  nor _70847_ (_19573_, _19572_, _19529_);
  nor _70848_ (_19574_, _19573_, _04481_);
  and _70849_ (_19575_, _06592_, _05251_);
  nor _70850_ (_19576_, _19522_, _07400_);
  not _70851_ (_19577_, _19576_);
  nor _70852_ (_19579_, _19577_, _19575_);
  or _70853_ (_19580_, _19579_, _03222_);
  nor _70854_ (_19581_, _19580_, _19574_);
  nor _70855_ (_19582_, _12718_, _09129_);
  nor _70856_ (_19583_, _19522_, _19582_);
  nor _70857_ (_19584_, _19583_, _03589_);
  or _70858_ (_19585_, _19584_, _03601_);
  nor _70859_ (_19586_, _19585_, _19581_);
  nor _70860_ (_19587_, _19586_, _19526_);
  or _70861_ (_19588_, _19587_, _03600_);
  and _70862_ (_19590_, _12733_, _05251_);
  or _70863_ (_19591_, _19590_, _19522_);
  or _70864_ (_19592_, _19591_, _07766_);
  and _70865_ (_19593_, _19592_, _07778_);
  and _70866_ (_19594_, _19593_, _19588_);
  and _70867_ (_19595_, _12739_, _05251_);
  nor _70868_ (_19596_, _19595_, _19522_);
  nor _70869_ (_19597_, _19596_, _07778_);
  nor _70870_ (_19598_, _19597_, _19594_);
  nor _70871_ (_19599_, _19598_, _03622_);
  nor _70872_ (_19601_, _19522_, _05567_);
  not _70873_ (_19602_, _19601_);
  nor _70874_ (_19603_, _19525_, _07777_);
  and _70875_ (_19604_, _19603_, _19602_);
  nor _70876_ (_19605_, _19604_, _19599_);
  nor _70877_ (_19606_, _19605_, _03790_);
  nor _70878_ (_19607_, _19531_, _06828_);
  and _70879_ (_19608_, _19607_, _19602_);
  nor _70880_ (_19609_, _19608_, _03624_);
  not _70881_ (_19610_, _19609_);
  nor _70882_ (_19612_, _19610_, _19606_);
  nor _70883_ (_19613_, _12732_, _09129_);
  or _70884_ (_19614_, _19522_, _07795_);
  nor _70885_ (_19615_, _19614_, _19613_);
  or _70886_ (_19616_, _19615_, _03785_);
  nor _70887_ (_19617_, _19616_, _19612_);
  nor _70888_ (_19618_, _12738_, _09129_);
  nor _70889_ (_19619_, _19618_, _19522_);
  nor _70890_ (_19620_, _19619_, _07793_);
  or _70891_ (_19621_, _19620_, _19617_);
  and _70892_ (_19623_, _19621_, _04246_);
  nor _70893_ (_19624_, _19538_, _04246_);
  or _70894_ (_19625_, _19624_, _19623_);
  and _70895_ (_19626_, _19625_, _03823_);
  nor _70896_ (_19627_, _19557_, _03823_);
  or _70897_ (_19628_, _19627_, _19626_);
  and _70898_ (_19629_, _19628_, _03514_);
  and _70899_ (_19630_, _12794_, _05251_);
  nor _70900_ (_19631_, _19630_, _19522_);
  nor _70901_ (_19632_, _19631_, _03514_);
  or _70902_ (_19634_, _19632_, _19629_);
  or _70903_ (_19635_, _19634_, _43004_);
  or _70904_ (_19636_, _43000_, \oc8051_golden_model_1.IP [3]);
  and _70905_ (_19637_, _19636_, _41806_);
  and _70906_ (_43530_, _19637_, _19635_);
  not _70907_ (_19638_, \oc8051_golden_model_1.IP [4]);
  nor _70908_ (_19639_, _05251_, _19638_);
  nor _70909_ (_19640_, _05777_, _09129_);
  nor _70910_ (_19641_, _19640_, _19639_);
  and _70911_ (_19642_, _19641_, _07390_);
  nor _70912_ (_19644_, _05908_, _19638_);
  and _70913_ (_19645_, _12827_, _05908_);
  nor _70914_ (_19646_, _19645_, _19644_);
  nor _70915_ (_19647_, _19646_, _03736_);
  and _70916_ (_19648_, _05251_, \oc8051_golden_model_1.ACC [4]);
  nor _70917_ (_19649_, _19648_, _19639_);
  nor _70918_ (_19650_, _19649_, _09029_);
  nor _70919_ (_19651_, _04409_, _19638_);
  or _70920_ (_19652_, _19651_, _19650_);
  and _70921_ (_19653_, _19652_, _04081_);
  nor _70922_ (_19655_, _12841_, _09129_);
  nor _70923_ (_19656_, _19655_, _19639_);
  nor _70924_ (_19657_, _19656_, _04081_);
  or _70925_ (_19658_, _19657_, _19653_);
  and _70926_ (_19659_, _19658_, _04055_);
  and _70927_ (_19660_, _12845_, _05908_);
  nor _70928_ (_19661_, _19660_, _19644_);
  nor _70929_ (_19662_, _19661_, _04055_);
  or _70930_ (_19663_, _19662_, _03723_);
  or _70931_ (_19664_, _19663_, _19659_);
  nand _70932_ (_19666_, _19641_, _03723_);
  and _70933_ (_19667_, _19666_, _19664_);
  and _70934_ (_19668_, _19667_, _03737_);
  nor _70935_ (_19669_, _19649_, _03737_);
  or _70936_ (_19670_, _19669_, _19668_);
  and _70937_ (_19671_, _19670_, _03736_);
  nor _70938_ (_19672_, _19671_, _19647_);
  nor _70939_ (_19673_, _19672_, _03719_);
  nor _70940_ (_19674_, _19644_, _12860_);
  or _70941_ (_19675_, _19661_, _06840_);
  nor _70942_ (_19677_, _19675_, _19674_);
  nor _70943_ (_19678_, _19677_, _19673_);
  nor _70944_ (_19679_, _19678_, _03505_);
  nor _70945_ (_19680_, _12825_, _09166_);
  nor _70946_ (_19681_, _19680_, _19644_);
  nor _70947_ (_19682_, _19681_, _03710_);
  nor _70948_ (_19683_, _19682_, _07390_);
  not _70949_ (_19684_, _19683_);
  nor _70950_ (_19685_, _19684_, _19679_);
  nor _70951_ (_19686_, _19685_, _19642_);
  nor _70952_ (_19688_, _19686_, _04481_);
  and _70953_ (_19689_, _06730_, _05251_);
  nor _70954_ (_19690_, _19639_, _07400_);
  not _70955_ (_19691_, _19690_);
  nor _70956_ (_19692_, _19691_, _19689_);
  nor _70957_ (_19693_, _19692_, _03222_);
  not _70958_ (_19694_, _19693_);
  nor _70959_ (_19695_, _19694_, _19688_);
  nor _70960_ (_19696_, _12933_, _09129_);
  nor _70961_ (_19697_, _19696_, _19639_);
  nor _70962_ (_19699_, _19697_, _03589_);
  or _70963_ (_19700_, _19699_, _08828_);
  or _70964_ (_19701_, _19700_, _19695_);
  and _70965_ (_19702_, _12821_, _05251_);
  or _70966_ (_19703_, _19639_, _07766_);
  or _70967_ (_19704_, _19703_, _19702_);
  and _70968_ (_19705_, _06298_, _05251_);
  nor _70969_ (_19706_, _19705_, _19639_);
  and _70970_ (_19707_, _19706_, _03601_);
  nor _70971_ (_19708_, _19707_, _03780_);
  and _70972_ (_19710_, _19708_, _19704_);
  and _70973_ (_19711_, _19710_, _19701_);
  and _70974_ (_19712_, _12817_, _05251_);
  nor _70975_ (_19713_, _19712_, _19639_);
  nor _70976_ (_19714_, _19713_, _07778_);
  nor _70977_ (_19715_, _19714_, _19711_);
  nor _70978_ (_19716_, _19715_, _03622_);
  nor _70979_ (_19717_, _19639_, _05825_);
  not _70980_ (_19718_, _19717_);
  nor _70981_ (_19719_, _19706_, _07777_);
  and _70982_ (_19721_, _19719_, _19718_);
  nor _70983_ (_19722_, _19721_, _19716_);
  nor _70984_ (_19723_, _19722_, _03790_);
  nor _70985_ (_19724_, _19649_, _06828_);
  and _70986_ (_19725_, _19724_, _19718_);
  or _70987_ (_19726_, _19725_, _19723_);
  and _70988_ (_19727_, _19726_, _07795_);
  nor _70989_ (_19728_, _12819_, _09129_);
  nor _70990_ (_19729_, _19728_, _19639_);
  nor _70991_ (_19730_, _19729_, _07795_);
  or _70992_ (_19732_, _19730_, _19727_);
  and _70993_ (_19733_, _19732_, _07793_);
  nor _70994_ (_19734_, _12816_, _09129_);
  nor _70995_ (_19735_, _19734_, _19639_);
  nor _70996_ (_19736_, _19735_, _07793_);
  or _70997_ (_19737_, _19736_, _19733_);
  and _70998_ (_19738_, _19737_, _04246_);
  nor _70999_ (_19739_, _19656_, _04246_);
  or _71000_ (_19740_, _19739_, _19738_);
  and _71001_ (_19741_, _19740_, _03823_);
  nor _71002_ (_19743_, _19646_, _03823_);
  or _71003_ (_19744_, _19743_, _19741_);
  and _71004_ (_19745_, _19744_, _03514_);
  and _71005_ (_19746_, _13003_, _05251_);
  nor _71006_ (_19747_, _19746_, _19639_);
  nor _71007_ (_19748_, _19747_, _03514_);
  or _71008_ (_19749_, _19748_, _19745_);
  or _71009_ (_19750_, _19749_, _43004_);
  or _71010_ (_19751_, _43000_, \oc8051_golden_model_1.IP [4]);
  and _71011_ (_19752_, _19751_, _41806_);
  and _71012_ (_43531_, _19752_, _19750_);
  not _71013_ (_19754_, \oc8051_golden_model_1.IP [5]);
  nor _71014_ (_19755_, _05251_, _19754_);
  and _71015_ (_19756_, _06684_, _05251_);
  or _71016_ (_19757_, _19756_, _19755_);
  and _71017_ (_19758_, _19757_, _04481_);
  and _71018_ (_19759_, _05251_, \oc8051_golden_model_1.ACC [5]);
  nor _71019_ (_19760_, _19759_, _19755_);
  nor _71020_ (_19761_, _19760_, _09029_);
  nor _71021_ (_19762_, _04409_, _19754_);
  or _71022_ (_19764_, _19762_, _19761_);
  and _71023_ (_19765_, _19764_, _04081_);
  nor _71024_ (_19766_, _13014_, _09129_);
  nor _71025_ (_19767_, _19766_, _19755_);
  nor _71026_ (_19768_, _19767_, _04081_);
  or _71027_ (_19769_, _19768_, _19765_);
  and _71028_ (_19770_, _19769_, _04055_);
  nor _71029_ (_19771_, _05908_, _19754_);
  and _71030_ (_19772_, _13037_, _05908_);
  nor _71031_ (_19773_, _19772_, _19771_);
  nor _71032_ (_19775_, _19773_, _04055_);
  or _71033_ (_19776_, _19775_, _03723_);
  or _71034_ (_19777_, _19776_, _19770_);
  nor _71035_ (_19778_, _05469_, _09129_);
  nor _71036_ (_19779_, _19778_, _19755_);
  nand _71037_ (_19780_, _19779_, _03723_);
  and _71038_ (_19781_, _19780_, _19777_);
  and _71039_ (_19782_, _19781_, _03737_);
  nor _71040_ (_19783_, _19760_, _03737_);
  or _71041_ (_19784_, _19783_, _19782_);
  and _71042_ (_19786_, _19784_, _03736_);
  and _71043_ (_19787_, _13047_, _05908_);
  nor _71044_ (_19788_, _19787_, _19771_);
  nor _71045_ (_19789_, _19788_, _03736_);
  or _71046_ (_19790_, _19789_, _19786_);
  and _71047_ (_19791_, _19790_, _06840_);
  nor _71048_ (_19792_, _19771_, _13054_);
  nor _71049_ (_19793_, _19792_, _19773_);
  and _71050_ (_19794_, _19793_, _03719_);
  or _71051_ (_19795_, _19794_, _19791_);
  and _71052_ (_19797_, _19795_, _03710_);
  nor _71053_ (_19798_, _13020_, _09166_);
  nor _71054_ (_19799_, _19798_, _19771_);
  nor _71055_ (_19800_, _19799_, _03710_);
  nor _71056_ (_19801_, _19800_, _07390_);
  not _71057_ (_19802_, _19801_);
  nor _71058_ (_19803_, _19802_, _19797_);
  and _71059_ (_19804_, _19779_, _07390_);
  or _71060_ (_19805_, _19804_, _04481_);
  nor _71061_ (_19806_, _19805_, _19803_);
  or _71062_ (_19808_, _19806_, _19758_);
  and _71063_ (_19809_, _19808_, _03589_);
  nor _71064_ (_19810_, _13127_, _09129_);
  nor _71065_ (_19811_, _19810_, _19755_);
  nor _71066_ (_19812_, _19811_, _03589_);
  or _71067_ (_19813_, _19812_, _08828_);
  or _71068_ (_19814_, _19813_, _19809_);
  and _71069_ (_19815_, _13141_, _05251_);
  or _71070_ (_19816_, _19755_, _07766_);
  or _71071_ (_19817_, _19816_, _19815_);
  and _71072_ (_19819_, _06306_, _05251_);
  nor _71073_ (_19820_, _19819_, _19755_);
  and _71074_ (_19821_, _19820_, _03601_);
  nor _71075_ (_19822_, _19821_, _03780_);
  and _71076_ (_19823_, _19822_, _19817_);
  and _71077_ (_19824_, _19823_, _19814_);
  and _71078_ (_19825_, _13147_, _05251_);
  nor _71079_ (_19826_, _19825_, _19755_);
  nor _71080_ (_19827_, _19826_, _07778_);
  nor _71081_ (_19828_, _19827_, _19824_);
  nor _71082_ (_19830_, _19828_, _03622_);
  nor _71083_ (_19831_, _19755_, _05518_);
  not _71084_ (_19832_, _19831_);
  nor _71085_ (_19833_, _19820_, _07777_);
  and _71086_ (_19834_, _19833_, _19832_);
  nor _71087_ (_19835_, _19834_, _19830_);
  nor _71088_ (_19836_, _19835_, _03790_);
  nor _71089_ (_19837_, _19760_, _06828_);
  and _71090_ (_19838_, _19837_, _19832_);
  or _71091_ (_19839_, _19838_, _19836_);
  and _71092_ (_19841_, _19839_, _07795_);
  nor _71093_ (_19842_, _13140_, _09129_);
  nor _71094_ (_19843_, _19842_, _19755_);
  nor _71095_ (_19844_, _19843_, _07795_);
  or _71096_ (_19845_, _19844_, _19841_);
  and _71097_ (_19846_, _19845_, _07793_);
  nor _71098_ (_19847_, _13146_, _09129_);
  nor _71099_ (_19848_, _19847_, _19755_);
  nor _71100_ (_19849_, _19848_, _07793_);
  or _71101_ (_19850_, _19849_, _19846_);
  and _71102_ (_19852_, _19850_, _04246_);
  nor _71103_ (_19853_, _19767_, _04246_);
  or _71104_ (_19854_, _19853_, _19852_);
  and _71105_ (_19855_, _19854_, _03823_);
  nor _71106_ (_19856_, _19788_, _03823_);
  or _71107_ (_19857_, _19856_, _19855_);
  and _71108_ (_19858_, _19857_, _03514_);
  and _71109_ (_19859_, _13199_, _05251_);
  nor _71110_ (_19860_, _19859_, _19755_);
  nor _71111_ (_19861_, _19860_, _03514_);
  or _71112_ (_19863_, _19861_, _19858_);
  or _71113_ (_19864_, _19863_, _43004_);
  or _71114_ (_19865_, _43000_, \oc8051_golden_model_1.IP [5]);
  and _71115_ (_19866_, _19865_, _41806_);
  and _71116_ (_43532_, _19866_, _19864_);
  not _71117_ (_19867_, \oc8051_golden_model_1.IP [6]);
  nor _71118_ (_19868_, _05251_, _19867_);
  and _71119_ (_19869_, _06455_, _05251_);
  or _71120_ (_19870_, _19869_, _19868_);
  and _71121_ (_19871_, _19870_, _04481_);
  and _71122_ (_19873_, _05251_, \oc8051_golden_model_1.ACC [6]);
  nor _71123_ (_19874_, _19873_, _19868_);
  nor _71124_ (_19875_, _19874_, _09029_);
  nor _71125_ (_19876_, _04409_, _19867_);
  or _71126_ (_19877_, _19876_, _19875_);
  and _71127_ (_19878_, _19877_, _04081_);
  nor _71128_ (_19879_, _13242_, _09129_);
  nor _71129_ (_19880_, _19879_, _19868_);
  nor _71130_ (_19881_, _19880_, _04081_);
  or _71131_ (_19882_, _19881_, _19878_);
  and _71132_ (_19884_, _19882_, _04055_);
  nor _71133_ (_19885_, _05908_, _19867_);
  and _71134_ (_19886_, _13229_, _05908_);
  nor _71135_ (_19887_, _19886_, _19885_);
  nor _71136_ (_19888_, _19887_, _04055_);
  or _71137_ (_19889_, _19888_, _03723_);
  or _71138_ (_19890_, _19889_, _19884_);
  nor _71139_ (_19891_, _05363_, _09129_);
  nor _71140_ (_19892_, _19891_, _19868_);
  nand _71141_ (_19893_, _19892_, _03723_);
  and _71142_ (_19895_, _19893_, _19890_);
  and _71143_ (_19896_, _19895_, _03737_);
  nor _71144_ (_19897_, _19874_, _03737_);
  or _71145_ (_19898_, _19897_, _19896_);
  and _71146_ (_19899_, _19898_, _03736_);
  and _71147_ (_19900_, _13253_, _05908_);
  nor _71148_ (_19901_, _19900_, _19885_);
  nor _71149_ (_19902_, _19901_, _03736_);
  or _71150_ (_19903_, _19902_, _03719_);
  or _71151_ (_19904_, _19903_, _19899_);
  nor _71152_ (_19906_, _19885_, _13260_);
  nor _71153_ (_19907_, _19906_, _19887_);
  or _71154_ (_19908_, _19907_, _06840_);
  and _71155_ (_19909_, _19908_, _03710_);
  and _71156_ (_19910_, _19909_, _19904_);
  nor _71157_ (_19911_, _13226_, _09166_);
  nor _71158_ (_19912_, _19911_, _19885_);
  nor _71159_ (_19913_, _19912_, _03710_);
  nor _71160_ (_19914_, _19913_, _07390_);
  not _71161_ (_19915_, _19914_);
  nor _71162_ (_19917_, _19915_, _19910_);
  and _71163_ (_19918_, _19892_, _07390_);
  or _71164_ (_19919_, _19918_, _04481_);
  nor _71165_ (_19920_, _19919_, _19917_);
  or _71166_ (_19921_, _19920_, _19871_);
  and _71167_ (_19922_, _19921_, _03589_);
  nor _71168_ (_19923_, _13332_, _09129_);
  nor _71169_ (_19924_, _19923_, _19868_);
  nor _71170_ (_19925_, _19924_, _03589_);
  or _71171_ (_19926_, _19925_, _08828_);
  or _71172_ (_19928_, _19926_, _19922_);
  and _71173_ (_19929_, _13347_, _05251_);
  or _71174_ (_19930_, _19868_, _07766_);
  or _71175_ (_19931_, _19930_, _19929_);
  and _71176_ (_19932_, _13339_, _05251_);
  nor _71177_ (_19933_, _19932_, _19868_);
  and _71178_ (_19934_, _19933_, _03601_);
  nor _71179_ (_19935_, _19934_, _03780_);
  and _71180_ (_19936_, _19935_, _19931_);
  and _71181_ (_19937_, _19936_, _19928_);
  and _71182_ (_19939_, _13353_, _05251_);
  nor _71183_ (_19940_, _19939_, _19868_);
  nor _71184_ (_19941_, _19940_, _07778_);
  nor _71185_ (_19942_, _19941_, _19937_);
  nor _71186_ (_19943_, _19942_, _03622_);
  nor _71187_ (_19944_, _19868_, _05412_);
  not _71188_ (_19945_, _19944_);
  nor _71189_ (_19946_, _19933_, _07777_);
  and _71190_ (_19947_, _19946_, _19945_);
  nor _71191_ (_19948_, _19947_, _19943_);
  nor _71192_ (_19950_, _19948_, _03790_);
  nor _71193_ (_19951_, _19874_, _06828_);
  and _71194_ (_19952_, _19951_, _19945_);
  or _71195_ (_19953_, _19952_, _19950_);
  and _71196_ (_19954_, _19953_, _07795_);
  nor _71197_ (_19955_, _13346_, _09129_);
  nor _71198_ (_19956_, _19955_, _19868_);
  nor _71199_ (_19957_, _19956_, _07795_);
  or _71200_ (_19958_, _19957_, _19954_);
  and _71201_ (_19959_, _19958_, _07793_);
  nor _71202_ (_19961_, _13352_, _09129_);
  nor _71203_ (_19962_, _19961_, _19868_);
  nor _71204_ (_19963_, _19962_, _07793_);
  or _71205_ (_19964_, _19963_, _19959_);
  and _71206_ (_19965_, _19964_, _04246_);
  nor _71207_ (_19966_, _19880_, _04246_);
  or _71208_ (_19967_, _19966_, _19965_);
  and _71209_ (_19968_, _19967_, _03823_);
  nor _71210_ (_19969_, _19901_, _03823_);
  or _71211_ (_19970_, _19969_, _19968_);
  and _71212_ (_19972_, _19970_, _03514_);
  and _71213_ (_19973_, _13402_, _05251_);
  nor _71214_ (_19974_, _19973_, _19868_);
  nor _71215_ (_19975_, _19974_, _03514_);
  or _71216_ (_19976_, _19975_, _19972_);
  or _71217_ (_19977_, _19976_, _43004_);
  or _71218_ (_19978_, _43000_, \oc8051_golden_model_1.IP [6]);
  and _71219_ (_19979_, _19978_, _41806_);
  and _71220_ (_43533_, _19979_, _19977_);
  not _71221_ (_19980_, \oc8051_golden_model_1.P0 [0]);
  nor _71222_ (_19982_, _43000_, _19980_);
  or _71223_ (_19983_, _19982_, rst);
  nor _71224_ (_19984_, _05293_, _19980_);
  and _71225_ (_19985_, _12128_, _05293_);
  or _71226_ (_19986_, _19985_, _19984_);
  and _71227_ (_19987_, _19986_, _03780_);
  and _71228_ (_19988_, _05293_, _04620_);
  or _71229_ (_19989_, _19988_, _19984_);
  or _71230_ (_19990_, _19989_, _06838_);
  nor _71231_ (_19991_, _05666_, _09236_);
  or _71232_ (_19993_, _19991_, _19984_);
  and _71233_ (_19994_, _19993_, _03610_);
  nor _71234_ (_19995_, _04409_, _19980_);
  and _71235_ (_19996_, _05293_, \oc8051_golden_model_1.ACC [0]);
  or _71236_ (_19997_, _19996_, _19984_);
  and _71237_ (_19998_, _19997_, _04409_);
  or _71238_ (_19999_, _19998_, _19995_);
  and _71239_ (_20000_, _19999_, _04081_);
  or _71240_ (_20001_, _20000_, _03715_);
  or _71241_ (_20002_, _20001_, _19994_);
  and _71242_ (_20004_, _12021_, _05209_);
  nor _71243_ (_20005_, _05209_, _19980_);
  or _71244_ (_20006_, _20005_, _04055_);
  or _71245_ (_20007_, _20006_, _20004_);
  and _71246_ (_20008_, _20007_, _03996_);
  and _71247_ (_20009_, _20008_, _20002_);
  and _71248_ (_20010_, _19989_, _03723_);
  or _71249_ (_20011_, _20010_, _03729_);
  or _71250_ (_20012_, _20011_, _20009_);
  or _71251_ (_20013_, _19997_, _03737_);
  and _71252_ (_20015_, _20013_, _03736_);
  and _71253_ (_20016_, _20015_, _20012_);
  and _71254_ (_20017_, _19984_, _03714_);
  or _71255_ (_20018_, _20017_, _03719_);
  or _71256_ (_20019_, _20018_, _20016_);
  or _71257_ (_20020_, _19993_, _06840_);
  and _71258_ (_20021_, _20020_, _03710_);
  and _71259_ (_20022_, _20021_, _20019_);
  or _71260_ (_20023_, _12051_, _12009_);
  and _71261_ (_20024_, _20023_, _05209_);
  or _71262_ (_20026_, _20024_, _20005_);
  and _71263_ (_20027_, _20026_, _03505_);
  or _71264_ (_20028_, _20027_, _07390_);
  or _71265_ (_20029_, _20028_, _20022_);
  and _71266_ (_20030_, _20029_, _19990_);
  or _71267_ (_20031_, _20030_, _04481_);
  and _71268_ (_20032_, _06546_, _05293_);
  or _71269_ (_20033_, _19984_, _07400_);
  or _71270_ (_20034_, _20033_, _20032_);
  and _71271_ (_20035_, _20034_, _03589_);
  and _71272_ (_20037_, _20035_, _20031_);
  and _71273_ (_20038_, _06340_, \oc8051_golden_model_1.P1 [0]);
  and _71274_ (_20039_, _06343_, \oc8051_golden_model_1.P0 [0]);
  and _71275_ (_20040_, _06346_, \oc8051_golden_model_1.P2 [0]);
  and _71276_ (_20041_, _06348_, \oc8051_golden_model_1.P3 [0]);
  or _71277_ (_20042_, _20041_, _20040_);
  or _71278_ (_20043_, _20042_, _20039_);
  nor _71279_ (_20044_, _20043_, _20038_);
  and _71280_ (_20045_, _20044_, _12076_);
  and _71281_ (_20046_, _20045_, _12090_);
  nand _71282_ (_20048_, _20046_, _12106_);
  or _71283_ (_20049_, _20048_, _12064_);
  and _71284_ (_20050_, _20049_, _05293_);
  or _71285_ (_20051_, _20050_, _19984_);
  and _71286_ (_20052_, _20051_, _03222_);
  or _71287_ (_20053_, _20052_, _20037_);
  or _71288_ (_20054_, _20053_, _08828_);
  and _71289_ (_20055_, _12124_, _05293_);
  or _71290_ (_20056_, _19984_, _07766_);
  or _71291_ (_20057_, _20056_, _20055_);
  and _71292_ (_20059_, _05293_, _06274_);
  or _71293_ (_20060_, _20059_, _19984_);
  or _71294_ (_20061_, _20060_, _05886_);
  and _71295_ (_20062_, _20061_, _07778_);
  and _71296_ (_20063_, _20062_, _20057_);
  and _71297_ (_20064_, _20063_, _20054_);
  or _71298_ (_20065_, _20064_, _19987_);
  and _71299_ (_20066_, _20065_, _07777_);
  nand _71300_ (_20067_, _20060_, _03622_);
  nor _71301_ (_20068_, _20067_, _19991_);
  or _71302_ (_20070_, _20068_, _20066_);
  and _71303_ (_20071_, _20070_, _06828_);
  or _71304_ (_20072_, _19984_, _05666_);
  and _71305_ (_20073_, _19997_, _03790_);
  and _71306_ (_20074_, _20073_, _20072_);
  or _71307_ (_20075_, _20074_, _03624_);
  or _71308_ (_20076_, _20075_, _20071_);
  nor _71309_ (_20077_, _12122_, _09236_);
  or _71310_ (_20078_, _19984_, _07795_);
  or _71311_ (_20079_, _20078_, _20077_);
  and _71312_ (_20081_, _20079_, _07793_);
  and _71313_ (_20082_, _20081_, _20076_);
  nor _71314_ (_20083_, _12003_, _09236_);
  or _71315_ (_20084_, _20083_, _19984_);
  and _71316_ (_20085_, _20084_, _03785_);
  or _71317_ (_20086_, _20085_, _03815_);
  or _71318_ (_20087_, _20086_, _20082_);
  or _71319_ (_20088_, _19993_, _04246_);
  and _71320_ (_20089_, _20088_, _03823_);
  and _71321_ (_20090_, _20089_, _20087_);
  and _71322_ (_20092_, _19984_, _03453_);
  or _71323_ (_20093_, _20092_, _03447_);
  or _71324_ (_20094_, _20093_, _20090_);
  or _71325_ (_20095_, _19993_, _03514_);
  and _71326_ (_20096_, _20095_, _43000_);
  and _71327_ (_20097_, _20096_, _20094_);
  or _71328_ (_43534_, _20097_, _19983_);
  or _71329_ (_20098_, _05293_, \oc8051_golden_model_1.P0 [1]);
  and _71330_ (_20099_, _12213_, _05293_);
  not _71331_ (_20100_, _20099_);
  and _71332_ (_20102_, _20100_, _20098_);
  or _71333_ (_20103_, _20102_, _04081_);
  nand _71334_ (_20104_, _05293_, _03274_);
  and _71335_ (_20105_, _20104_, _20098_);
  and _71336_ (_20106_, _20105_, _04409_);
  not _71337_ (_20107_, \oc8051_golden_model_1.P0 [1]);
  nor _71338_ (_20108_, _04409_, _20107_);
  or _71339_ (_20109_, _20108_, _03610_);
  or _71340_ (_20110_, _20109_, _20106_);
  and _71341_ (_20111_, _20110_, _04055_);
  and _71342_ (_20113_, _20111_, _20103_);
  and _71343_ (_20114_, _12224_, _05209_);
  nor _71344_ (_20115_, _05209_, _20107_);
  or _71345_ (_20116_, _20115_, _03723_);
  or _71346_ (_20117_, _20116_, _20114_);
  and _71347_ (_20118_, _20117_, _14265_);
  or _71348_ (_20119_, _20118_, _20113_);
  nor _71349_ (_20120_, _05293_, _20107_);
  and _71350_ (_20121_, _05293_, _06764_);
  or _71351_ (_20122_, _20121_, _20120_);
  or _71352_ (_20124_, _20122_, _03996_);
  and _71353_ (_20125_, _20124_, _20119_);
  or _71354_ (_20126_, _20125_, _03729_);
  or _71355_ (_20127_, _20105_, _03737_);
  and _71356_ (_20128_, _20127_, _03736_);
  and _71357_ (_20129_, _20128_, _20126_);
  and _71358_ (_20130_, _12211_, _05209_);
  or _71359_ (_20131_, _20130_, _20115_);
  and _71360_ (_20132_, _20131_, _03714_);
  or _71361_ (_20133_, _20132_, _03719_);
  or _71362_ (_20135_, _20133_, _20129_);
  and _71363_ (_20136_, _20114_, _12239_);
  or _71364_ (_20137_, _20115_, _06840_);
  or _71365_ (_20138_, _20137_, _20136_);
  and _71366_ (_20139_, _20138_, _20135_);
  and _71367_ (_20140_, _20139_, _03710_);
  or _71368_ (_20141_, _12255_, _12211_);
  and _71369_ (_20142_, _20141_, _05209_);
  or _71370_ (_20143_, _20115_, _20142_);
  and _71371_ (_20144_, _20143_, _03505_);
  or _71372_ (_20146_, _20144_, _07390_);
  or _71373_ (_20147_, _20146_, _20140_);
  or _71374_ (_20148_, _20122_, _06838_);
  and _71375_ (_20149_, _20148_, _20147_);
  or _71376_ (_20150_, _20149_, _04481_);
  and _71377_ (_20151_, _06501_, _05293_);
  or _71378_ (_20152_, _20120_, _07400_);
  or _71379_ (_20153_, _20152_, _20151_);
  and _71380_ (_20154_, _20153_, _03589_);
  and _71381_ (_20155_, _20154_, _20150_);
  and _71382_ (_20157_, _06340_, \oc8051_golden_model_1.P1 [1]);
  and _71383_ (_20158_, _06343_, \oc8051_golden_model_1.P0 [1]);
  and _71384_ (_20159_, _06346_, \oc8051_golden_model_1.P2 [1]);
  and _71385_ (_20160_, _06348_, \oc8051_golden_model_1.P3 [1]);
  or _71386_ (_20161_, _20160_, _20159_);
  or _71387_ (_20162_, _20161_, _20158_);
  nor _71388_ (_20163_, _20162_, _20157_);
  and _71389_ (_20164_, _20163_, _12280_);
  and _71390_ (_20165_, _20164_, _12294_);
  nand _71391_ (_20166_, _20165_, _12310_);
  or _71392_ (_20168_, _20166_, _12268_);
  and _71393_ (_20169_, _20168_, _05293_);
  or _71394_ (_20170_, _20169_, _20120_);
  and _71395_ (_20171_, _20170_, _03222_);
  or _71396_ (_20172_, _20171_, _20155_);
  and _71397_ (_20173_, _20172_, _03602_);
  or _71398_ (_20174_, _12327_, _09236_);
  and _71399_ (_20175_, _20174_, _03600_);
  nand _71400_ (_20176_, _05293_, _04303_);
  and _71401_ (_20177_, _20176_, _03601_);
  or _71402_ (_20179_, _20177_, _20175_);
  and _71403_ (_20180_, _20179_, _20098_);
  or _71404_ (_20181_, _20180_, _20173_);
  and _71405_ (_20182_, _20181_, _07778_);
  or _71406_ (_20183_, _12333_, _09236_);
  and _71407_ (_20184_, _20098_, _03780_);
  and _71408_ (_20185_, _20184_, _20183_);
  or _71409_ (_20186_, _20185_, _20182_);
  and _71410_ (_20187_, _20186_, _07777_);
  or _71411_ (_20188_, _12207_, _09236_);
  and _71412_ (_20190_, _20098_, _03622_);
  and _71413_ (_20191_, _20190_, _20188_);
  or _71414_ (_20192_, _20191_, _20187_);
  and _71415_ (_20193_, _20192_, _06828_);
  or _71416_ (_20194_, _20120_, _05618_);
  and _71417_ (_20195_, _20105_, _03790_);
  and _71418_ (_20196_, _20195_, _20194_);
  or _71419_ (_20197_, _20196_, _20193_);
  and _71420_ (_20198_, _20197_, _03786_);
  or _71421_ (_20199_, _20176_, _05618_);
  and _71422_ (_20201_, _20098_, _03624_);
  and _71423_ (_20202_, _20201_, _20199_);
  or _71424_ (_20203_, _20104_, _05618_);
  and _71425_ (_20204_, _20098_, _03785_);
  and _71426_ (_20205_, _20204_, _20203_);
  or _71427_ (_20206_, _20205_, _03815_);
  or _71428_ (_20207_, _20206_, _20202_);
  or _71429_ (_20208_, _20207_, _20198_);
  or _71430_ (_20209_, _20102_, _04246_);
  and _71431_ (_20210_, _20209_, _03823_);
  and _71432_ (_20212_, _20210_, _20208_);
  and _71433_ (_20213_, _20131_, _03453_);
  or _71434_ (_20214_, _20213_, _03447_);
  or _71435_ (_20215_, _20214_, _20212_);
  or _71436_ (_20216_, _20120_, _03514_);
  or _71437_ (_20217_, _20216_, _20099_);
  and _71438_ (_20218_, _20217_, _43000_);
  and _71439_ (_20219_, _20218_, _20215_);
  nor _71440_ (_20220_, _43000_, _20107_);
  or _71441_ (_20221_, _20220_, rst);
  or _71442_ (_43535_, _20221_, _20219_);
  not _71443_ (_20223_, \oc8051_golden_model_1.P0 [2]);
  nor _71444_ (_20224_, _05293_, _20223_);
  nor _71445_ (_20225_, _09236_, _04875_);
  or _71446_ (_20226_, _20225_, _20224_);
  or _71447_ (_20227_, _20226_, _06838_);
  and _71448_ (_20228_, _20226_, _03723_);
  nor _71449_ (_20229_, _05209_, _20223_);
  and _71450_ (_20230_, _12411_, _05209_);
  or _71451_ (_20231_, _20230_, _20229_);
  or _71452_ (_20233_, _20231_, _04055_);
  nor _71453_ (_20234_, _12416_, _09236_);
  or _71454_ (_20235_, _20234_, _20224_);
  and _71455_ (_20236_, _20235_, _03610_);
  nor _71456_ (_20237_, _04409_, _20223_);
  and _71457_ (_20238_, _05293_, \oc8051_golden_model_1.ACC [2]);
  or _71458_ (_20239_, _20238_, _20224_);
  and _71459_ (_20240_, _20239_, _04409_);
  or _71460_ (_20241_, _20240_, _20237_);
  and _71461_ (_20242_, _20241_, _04081_);
  or _71462_ (_20244_, _20242_, _03715_);
  or _71463_ (_20245_, _20244_, _20236_);
  and _71464_ (_20246_, _20245_, _20233_);
  and _71465_ (_20247_, _20246_, _03996_);
  or _71466_ (_20248_, _20247_, _20228_);
  or _71467_ (_20249_, _20248_, _03729_);
  or _71468_ (_20250_, _20239_, _03737_);
  and _71469_ (_20251_, _20250_, _03736_);
  and _71470_ (_20252_, _20251_, _20249_);
  and _71471_ (_20253_, _12409_, _05209_);
  or _71472_ (_20255_, _20253_, _20229_);
  and _71473_ (_20256_, _20255_, _03714_);
  or _71474_ (_20257_, _20256_, _03719_);
  or _71475_ (_20258_, _20257_, _20252_);
  or _71476_ (_20259_, _20229_, _12443_);
  and _71477_ (_20260_, _20259_, _20231_);
  or _71478_ (_20261_, _20260_, _06840_);
  and _71479_ (_20262_, _20261_, _03710_);
  and _71480_ (_20263_, _20262_, _20258_);
  or _71481_ (_20264_, _12460_, _12409_);
  and _71482_ (_20266_, _20264_, _05209_);
  or _71483_ (_20267_, _20266_, _20229_);
  and _71484_ (_20268_, _20267_, _03505_);
  or _71485_ (_20269_, _20268_, _07390_);
  or _71486_ (_20270_, _20269_, _20263_);
  and _71487_ (_20271_, _20270_, _20227_);
  or _71488_ (_20272_, _20271_, _04481_);
  and _71489_ (_20273_, _06637_, _05293_);
  or _71490_ (_20274_, _20224_, _07400_);
  or _71491_ (_20275_, _20274_, _20273_);
  and _71492_ (_20277_, _20275_, _03589_);
  and _71493_ (_20278_, _20277_, _20272_);
  and _71494_ (_20279_, _06340_, \oc8051_golden_model_1.P1 [2]);
  and _71495_ (_20280_, _06343_, \oc8051_golden_model_1.P0 [2]);
  and _71496_ (_20281_, _06346_, \oc8051_golden_model_1.P2 [2]);
  and _71497_ (_20282_, _06348_, \oc8051_golden_model_1.P3 [2]);
  or _71498_ (_20283_, _20282_, _20281_);
  or _71499_ (_20284_, _20283_, _20280_);
  nor _71500_ (_20285_, _20284_, _20279_);
  and _71501_ (_20286_, _20285_, _12486_);
  and _71502_ (_20288_, _20286_, _12496_);
  nand _71503_ (_20289_, _20288_, _12516_);
  or _71504_ (_20290_, _20289_, _12474_);
  and _71505_ (_20291_, _20290_, _05293_);
  or _71506_ (_20292_, _20224_, _20291_);
  and _71507_ (_20293_, _20292_, _03222_);
  or _71508_ (_20294_, _20293_, _20278_);
  or _71509_ (_20295_, _20294_, _08828_);
  and _71510_ (_20296_, _12533_, _05293_);
  or _71511_ (_20297_, _20224_, _07766_);
  or _71512_ (_20299_, _20297_, _20296_);
  and _71513_ (_20300_, _05293_, _06332_);
  or _71514_ (_20301_, _20300_, _20224_);
  or _71515_ (_20302_, _20301_, _05886_);
  and _71516_ (_20303_, _20302_, _07778_);
  and _71517_ (_20304_, _20303_, _20299_);
  and _71518_ (_20305_, _20304_, _20295_);
  and _71519_ (_20306_, _12539_, _05293_);
  or _71520_ (_20307_, _20306_, _20224_);
  and _71521_ (_20308_, _20307_, _03780_);
  or _71522_ (_20310_, _20308_, _20305_);
  and _71523_ (_20311_, _20310_, _07777_);
  or _71524_ (_20312_, _20224_, _05718_);
  and _71525_ (_20313_, _20301_, _03622_);
  and _71526_ (_20314_, _20313_, _20312_);
  or _71527_ (_20315_, _20314_, _20311_);
  and _71528_ (_20316_, _20315_, _06828_);
  and _71529_ (_20317_, _20239_, _03790_);
  and _71530_ (_20318_, _20317_, _20312_);
  or _71531_ (_20319_, _20318_, _03624_);
  or _71532_ (_20321_, _20319_, _20316_);
  nor _71533_ (_20322_, _12532_, _09236_);
  or _71534_ (_20323_, _20224_, _07795_);
  or _71535_ (_20324_, _20323_, _20322_);
  and _71536_ (_20325_, _20324_, _07793_);
  and _71537_ (_20326_, _20325_, _20321_);
  nor _71538_ (_20327_, _12538_, _09236_);
  or _71539_ (_20328_, _20327_, _20224_);
  and _71540_ (_20329_, _20328_, _03785_);
  or _71541_ (_20330_, _20329_, _03815_);
  or _71542_ (_20332_, _20330_, _20326_);
  or _71543_ (_20333_, _20235_, _04246_);
  and _71544_ (_20334_, _20333_, _03823_);
  and _71545_ (_20335_, _20334_, _20332_);
  and _71546_ (_20336_, _20255_, _03453_);
  or _71547_ (_20337_, _20336_, _03447_);
  or _71548_ (_20338_, _20337_, _20335_);
  and _71549_ (_20339_, _12592_, _05293_);
  or _71550_ (_20340_, _20224_, _03514_);
  or _71551_ (_20341_, _20340_, _20339_);
  and _71552_ (_20343_, _20341_, _43000_);
  and _71553_ (_20344_, _20343_, _20338_);
  nor _71554_ (_20345_, _43000_, _20223_);
  or _71555_ (_20346_, _20345_, rst);
  or _71556_ (_43536_, _20346_, _20344_);
  not _71557_ (_20347_, \oc8051_golden_model_1.P0 [3]);
  nor _71558_ (_20348_, _43000_, _20347_);
  or _71559_ (_20349_, _20348_, rst);
  nor _71560_ (_20350_, _05293_, _20347_);
  nor _71561_ (_20351_, _09236_, _05005_);
  or _71562_ (_20353_, _20351_, _20350_);
  or _71563_ (_20354_, _20353_, _06838_);
  nor _71564_ (_20355_, _12627_, _09236_);
  or _71565_ (_20356_, _20355_, _20350_);
  or _71566_ (_20357_, _20356_, _04081_);
  and _71567_ (_20358_, _05293_, \oc8051_golden_model_1.ACC [3]);
  or _71568_ (_20359_, _20358_, _20350_);
  and _71569_ (_20360_, _20359_, _04409_);
  nor _71570_ (_20361_, _04409_, _20347_);
  or _71571_ (_20362_, _20361_, _03610_);
  or _71572_ (_20364_, _20362_, _20360_);
  and _71573_ (_20365_, _20364_, _04055_);
  and _71574_ (_20366_, _20365_, _20357_);
  nor _71575_ (_20367_, _05209_, _20347_);
  and _71576_ (_20368_, _12631_, _05209_);
  or _71577_ (_20369_, _20368_, _20367_);
  and _71578_ (_20370_, _20369_, _03715_);
  or _71579_ (_20371_, _20370_, _03723_);
  or _71580_ (_20372_, _20371_, _20366_);
  or _71581_ (_20373_, _20353_, _03996_);
  and _71582_ (_20375_, _20373_, _20372_);
  or _71583_ (_20376_, _20375_, _03729_);
  or _71584_ (_20377_, _20359_, _03737_);
  and _71585_ (_20378_, _20377_, _03736_);
  and _71586_ (_20379_, _20378_, _20376_);
  and _71587_ (_20380_, _12641_, _05209_);
  or _71588_ (_20381_, _20380_, _20367_);
  and _71589_ (_20382_, _20381_, _03714_);
  or _71590_ (_20383_, _20382_, _03719_);
  or _71591_ (_20384_, _20383_, _20379_);
  or _71592_ (_20386_, _20367_, _12648_);
  and _71593_ (_20387_, _20386_, _20369_);
  or _71594_ (_20388_, _20387_, _06840_);
  and _71595_ (_20389_, _20388_, _03710_);
  and _71596_ (_20390_, _20389_, _20384_);
  or _71597_ (_20391_, _12641_, _12610_);
  and _71598_ (_20392_, _20391_, _05209_);
  or _71599_ (_20393_, _20392_, _20367_);
  and _71600_ (_20394_, _20393_, _03505_);
  or _71601_ (_20395_, _20394_, _07390_);
  or _71602_ (_20397_, _20395_, _20390_);
  and _71603_ (_20398_, _20397_, _20354_);
  or _71604_ (_20399_, _20398_, _04481_);
  and _71605_ (_20400_, _06592_, _05293_);
  or _71606_ (_20401_, _20350_, _07400_);
  or _71607_ (_20402_, _20401_, _20400_);
  and _71608_ (_20403_, _20402_, _03589_);
  and _71609_ (_20404_, _20403_, _20399_);
  and _71610_ (_20405_, _06343_, \oc8051_golden_model_1.P0 [3]);
  and _71611_ (_20406_, _06340_, \oc8051_golden_model_1.P1 [3]);
  and _71612_ (_20408_, _06346_, \oc8051_golden_model_1.P2 [3]);
  and _71613_ (_20409_, _06348_, \oc8051_golden_model_1.P3 [3]);
  or _71614_ (_20410_, _20409_, _20408_);
  or _71615_ (_20411_, _20410_, _20406_);
  nor _71616_ (_20412_, _20411_, _20405_);
  and _71617_ (_20413_, _20412_, _12713_);
  and _71618_ (_20414_, _20413_, _12700_);
  nand _71619_ (_20415_, _20414_, _12693_);
  or _71620_ (_20416_, _20415_, _12672_);
  and _71621_ (_20417_, _20416_, _05293_);
  or _71622_ (_20419_, _20350_, _20417_);
  and _71623_ (_20420_, _20419_, _03222_);
  or _71624_ (_20421_, _20420_, _20404_);
  or _71625_ (_20422_, _20421_, _08828_);
  and _71626_ (_20423_, _12733_, _05293_);
  or _71627_ (_20424_, _20350_, _07766_);
  or _71628_ (_20425_, _20424_, _20423_);
  and _71629_ (_20426_, _05293_, _06276_);
  or _71630_ (_20427_, _20426_, _20350_);
  or _71631_ (_20428_, _20427_, _05886_);
  and _71632_ (_20430_, _20428_, _07778_);
  and _71633_ (_20431_, _20430_, _20425_);
  and _71634_ (_20432_, _20431_, _20422_);
  and _71635_ (_20433_, _12739_, _05293_);
  or _71636_ (_20434_, _20433_, _20350_);
  and _71637_ (_20435_, _20434_, _03780_);
  or _71638_ (_20436_, _20435_, _20432_);
  and _71639_ (_20437_, _20436_, _07777_);
  or _71640_ (_20438_, _20350_, _05567_);
  and _71641_ (_20439_, _20427_, _03622_);
  and _71642_ (_20441_, _20439_, _20438_);
  or _71643_ (_20442_, _20441_, _20437_);
  and _71644_ (_20443_, _20442_, _06828_);
  and _71645_ (_20444_, _20359_, _03790_);
  and _71646_ (_20445_, _20444_, _20438_);
  or _71647_ (_20446_, _20445_, _03624_);
  or _71648_ (_20447_, _20446_, _20443_);
  nor _71649_ (_20448_, _12732_, _09236_);
  or _71650_ (_20449_, _20350_, _07795_);
  or _71651_ (_20450_, _20449_, _20448_);
  and _71652_ (_20452_, _20450_, _07793_);
  and _71653_ (_20453_, _20452_, _20447_);
  nor _71654_ (_20454_, _12738_, _09236_);
  or _71655_ (_20455_, _20454_, _20350_);
  and _71656_ (_20456_, _20455_, _03785_);
  or _71657_ (_20457_, _20456_, _03815_);
  or _71658_ (_20458_, _20457_, _20453_);
  or _71659_ (_20459_, _20356_, _04246_);
  and _71660_ (_20460_, _20459_, _03823_);
  and _71661_ (_20461_, _20460_, _20458_);
  and _71662_ (_20462_, _20381_, _03453_);
  or _71663_ (_20463_, _20462_, _03447_);
  or _71664_ (_20464_, _20463_, _20461_);
  and _71665_ (_20465_, _12794_, _05293_);
  or _71666_ (_20466_, _20350_, _03514_);
  or _71667_ (_20467_, _20466_, _20465_);
  and _71668_ (_20468_, _20467_, _43000_);
  and _71669_ (_20469_, _20468_, _20464_);
  or _71670_ (_43537_, _20469_, _20349_);
  and _71671_ (_20470_, _09236_, \oc8051_golden_model_1.P0 [4]);
  nor _71672_ (_20472_, _05777_, _09236_);
  or _71673_ (_20473_, _20472_, _20470_);
  or _71674_ (_20474_, _20473_, _06838_);
  not _71675_ (_20475_, \oc8051_golden_model_1.P0 [4]);
  nor _71676_ (_20476_, _05209_, _20475_);
  and _71677_ (_20477_, _12827_, _05209_);
  or _71678_ (_20478_, _20477_, _20476_);
  and _71679_ (_20479_, _20478_, _03714_);
  nor _71680_ (_20480_, _12841_, _09236_);
  or _71681_ (_20481_, _20480_, _20470_);
  or _71682_ (_20483_, _20481_, _04081_);
  and _71683_ (_20484_, _05293_, \oc8051_golden_model_1.ACC [4]);
  or _71684_ (_20485_, _20484_, _20470_);
  and _71685_ (_20486_, _20485_, _04409_);
  nor _71686_ (_20487_, _04409_, _20475_);
  or _71687_ (_20488_, _20487_, _03610_);
  or _71688_ (_20489_, _20488_, _20486_);
  and _71689_ (_20490_, _20489_, _04055_);
  and _71690_ (_20491_, _20490_, _20483_);
  and _71691_ (_20492_, _12845_, _05209_);
  or _71692_ (_20494_, _20492_, _20476_);
  and _71693_ (_20495_, _20494_, _03715_);
  or _71694_ (_20496_, _20495_, _03723_);
  or _71695_ (_20497_, _20496_, _20491_);
  or _71696_ (_20498_, _20473_, _03996_);
  and _71697_ (_20499_, _20498_, _20497_);
  or _71698_ (_20500_, _20499_, _03729_);
  or _71699_ (_20501_, _20485_, _03737_);
  and _71700_ (_20502_, _20501_, _03736_);
  and _71701_ (_20503_, _20502_, _20500_);
  or _71702_ (_20504_, _20503_, _20479_);
  and _71703_ (_20505_, _20504_, _06840_);
  and _71704_ (_20506_, _12861_, _05209_);
  or _71705_ (_20507_, _20506_, _20476_);
  and _71706_ (_20508_, _20507_, _03719_);
  or _71707_ (_20509_, _20508_, _20505_);
  and _71708_ (_20510_, _20509_, _03710_);
  or _71709_ (_20511_, _12827_, _12824_);
  and _71710_ (_20512_, _20511_, _05209_);
  or _71711_ (_20513_, _20512_, _20476_);
  and _71712_ (_20515_, _20513_, _03505_);
  or _71713_ (_20516_, _20515_, _07390_);
  or _71714_ (_20517_, _20516_, _20510_);
  and _71715_ (_20518_, _20517_, _20474_);
  or _71716_ (_20519_, _20518_, _04481_);
  and _71717_ (_20520_, _06730_, _05293_);
  or _71718_ (_20521_, _20470_, _07400_);
  or _71719_ (_20522_, _20521_, _20520_);
  and _71720_ (_20523_, _20522_, _03589_);
  and _71721_ (_20524_, _20523_, _20519_);
  and _71722_ (_20526_, _06343_, \oc8051_golden_model_1.P0 [4]);
  and _71723_ (_20527_, _06340_, \oc8051_golden_model_1.P1 [4]);
  and _71724_ (_20528_, _06346_, \oc8051_golden_model_1.P2 [4]);
  and _71725_ (_20529_, _06348_, \oc8051_golden_model_1.P3 [4]);
  or _71726_ (_20530_, _20529_, _20528_);
  or _71727_ (_20531_, _20530_, _20527_);
  nor _71728_ (_20532_, _20531_, _20526_);
  and _71729_ (_20533_, _20532_, _12899_);
  and _71730_ (_20534_, _20533_, _12913_);
  nand _71731_ (_20535_, _20534_, _12930_);
  or _71732_ (_20536_, _20535_, _12887_);
  and _71733_ (_20537_, _20536_, _05293_);
  or _71734_ (_20538_, _20537_, _20470_);
  and _71735_ (_20539_, _20538_, _03222_);
  or _71736_ (_20540_, _20539_, _08828_);
  or _71737_ (_20541_, _20540_, _20524_);
  and _71738_ (_20542_, _12821_, _05293_);
  or _71739_ (_20543_, _20470_, _07766_);
  or _71740_ (_20544_, _20543_, _20542_);
  and _71741_ (_20545_, _06298_, _05293_);
  or _71742_ (_20547_, _20545_, _20470_);
  or _71743_ (_20548_, _20547_, _05886_);
  and _71744_ (_20549_, _20548_, _07778_);
  and _71745_ (_20550_, _20549_, _20544_);
  and _71746_ (_20551_, _20550_, _20541_);
  and _71747_ (_20552_, _12817_, _05293_);
  or _71748_ (_20553_, _20552_, _20470_);
  and _71749_ (_20554_, _20553_, _03780_);
  or _71750_ (_20555_, _20554_, _20551_);
  and _71751_ (_20556_, _20555_, _07777_);
  or _71752_ (_20558_, _20470_, _05825_);
  and _71753_ (_20559_, _20547_, _03622_);
  and _71754_ (_20560_, _20559_, _20558_);
  or _71755_ (_20561_, _20560_, _20556_);
  and _71756_ (_20562_, _20561_, _06828_);
  and _71757_ (_20563_, _20485_, _03790_);
  and _71758_ (_20564_, _20563_, _20558_);
  or _71759_ (_20565_, _20564_, _03624_);
  or _71760_ (_20566_, _20565_, _20562_);
  nor _71761_ (_20567_, _12819_, _09236_);
  or _71762_ (_20568_, _20470_, _07795_);
  or _71763_ (_20569_, _20568_, _20567_);
  and _71764_ (_20570_, _20569_, _07793_);
  and _71765_ (_20571_, _20570_, _20566_);
  nor _71766_ (_20572_, _12816_, _09236_);
  or _71767_ (_20573_, _20572_, _20470_);
  and _71768_ (_20574_, _20573_, _03785_);
  or _71769_ (_20575_, _20574_, _03815_);
  or _71770_ (_20576_, _20575_, _20571_);
  or _71771_ (_20577_, _20481_, _04246_);
  and _71772_ (_20579_, _20577_, _03823_);
  and _71773_ (_20580_, _20579_, _20576_);
  and _71774_ (_20581_, _20478_, _03453_);
  or _71775_ (_20582_, _20581_, _03447_);
  or _71776_ (_20583_, _20582_, _20580_);
  and _71777_ (_20584_, _13003_, _05293_);
  or _71778_ (_20585_, _20470_, _03514_);
  or _71779_ (_20586_, _20585_, _20584_);
  and _71780_ (_20587_, _20586_, _43000_);
  and _71781_ (_20588_, _20587_, _20583_);
  nor _71782_ (_20590_, \oc8051_golden_model_1.P0 [4], rst);
  nor _71783_ (_20591_, _20590_, _04794_);
  or _71784_ (_43538_, _20591_, _20588_);
  not _71785_ (_20592_, \oc8051_golden_model_1.P0 [5]);
  nor _71786_ (_20593_, _43000_, _20592_);
  or _71787_ (_20594_, _20593_, rst);
  nor _71788_ (_20595_, _05293_, _20592_);
  nor _71789_ (_20596_, _13014_, _09236_);
  or _71790_ (_20597_, _20596_, _20595_);
  or _71791_ (_20598_, _20597_, _04081_);
  and _71792_ (_20599_, _05293_, \oc8051_golden_model_1.ACC [5]);
  or _71793_ (_20600_, _20599_, _20595_);
  and _71794_ (_20601_, _20600_, _04409_);
  nor _71795_ (_20602_, _04409_, _20592_);
  or _71796_ (_20603_, _20602_, _03610_);
  or _71797_ (_20604_, _20603_, _20601_);
  and _71798_ (_20605_, _20604_, _04055_);
  and _71799_ (_20606_, _20605_, _20598_);
  nor _71800_ (_20607_, _05209_, _20592_);
  and _71801_ (_20608_, _13037_, _05209_);
  or _71802_ (_20610_, _20608_, _20607_);
  and _71803_ (_20611_, _20610_, _03715_);
  or _71804_ (_20612_, _20611_, _03723_);
  or _71805_ (_20613_, _20612_, _20606_);
  nor _71806_ (_20614_, _05469_, _09236_);
  or _71807_ (_20615_, _20614_, _20595_);
  or _71808_ (_20616_, _20615_, _03996_);
  and _71809_ (_20617_, _20616_, _20613_);
  or _71810_ (_20618_, _20617_, _03729_);
  or _71811_ (_20619_, _20600_, _03737_);
  and _71812_ (_20621_, _20619_, _03736_);
  and _71813_ (_20622_, _20621_, _20618_);
  and _71814_ (_20623_, _13047_, _05209_);
  or _71815_ (_20624_, _20623_, _20607_);
  and _71816_ (_20625_, _20624_, _03714_);
  or _71817_ (_20626_, _20625_, _03719_);
  or _71818_ (_20627_, _20626_, _20622_);
  or _71819_ (_20628_, _20607_, _13054_);
  and _71820_ (_20629_, _20628_, _20610_);
  or _71821_ (_20630_, _20629_, _06840_);
  and _71822_ (_20631_, _20630_, _03710_);
  and _71823_ (_20632_, _20631_, _20627_);
  or _71824_ (_20633_, _13047_, _13019_);
  and _71825_ (_20634_, _20633_, _05209_);
  or _71826_ (_20635_, _20634_, _20607_);
  and _71827_ (_20636_, _20635_, _03505_);
  or _71828_ (_20637_, _20636_, _07390_);
  or _71829_ (_20638_, _20637_, _20632_);
  or _71830_ (_20639_, _20615_, _06838_);
  and _71831_ (_20640_, _20639_, _20638_);
  or _71832_ (_20642_, _20640_, _04481_);
  and _71833_ (_20643_, _06684_, _05293_);
  or _71834_ (_20644_, _20595_, _07400_);
  or _71835_ (_20645_, _20644_, _20643_);
  and _71836_ (_20646_, _20645_, _03589_);
  and _71837_ (_20647_, _20646_, _20642_);
  and _71838_ (_20648_, _06340_, \oc8051_golden_model_1.P1 [5]);
  and _71839_ (_20649_, _06343_, \oc8051_golden_model_1.P0 [5]);
  and _71840_ (_20650_, _06346_, \oc8051_golden_model_1.P2 [5]);
  and _71841_ (_20651_, _06348_, \oc8051_golden_model_1.P3 [5]);
  or _71842_ (_20653_, _20651_, _20650_);
  or _71843_ (_20654_, _20653_, _20649_);
  or _71844_ (_20655_, _20654_, _20648_);
  nor _71845_ (_20656_, _20655_, _13103_);
  and _71846_ (_20657_, _20656_, _13122_);
  and _71847_ (_20658_, _20657_, _13102_);
  nand _71848_ (_20659_, _20658_, _13095_);
  or _71849_ (_20660_, _20659_, _13081_);
  and _71850_ (_20661_, _20660_, _05293_);
  or _71851_ (_20662_, _20661_, _20595_);
  and _71852_ (_20663_, _20662_, _03222_);
  or _71853_ (_20664_, _20663_, _08828_);
  or _71854_ (_20665_, _20664_, _20647_);
  and _71855_ (_20666_, _13141_, _05293_);
  or _71856_ (_20667_, _20595_, _07766_);
  or _71857_ (_20668_, _20667_, _20666_);
  and _71858_ (_20669_, _06306_, _05293_);
  or _71859_ (_20670_, _20669_, _20595_);
  or _71860_ (_20671_, _20670_, _05886_);
  and _71861_ (_20672_, _20671_, _07778_);
  and _71862_ (_20674_, _20672_, _20668_);
  and _71863_ (_20675_, _20674_, _20665_);
  and _71864_ (_20676_, _13147_, _05293_);
  or _71865_ (_20677_, _20676_, _20595_);
  and _71866_ (_20678_, _20677_, _03780_);
  or _71867_ (_20679_, _20678_, _20675_);
  and _71868_ (_20680_, _20679_, _07777_);
  or _71869_ (_20681_, _20595_, _05518_);
  and _71870_ (_20682_, _20670_, _03622_);
  and _71871_ (_20683_, _20682_, _20681_);
  or _71872_ (_20685_, _20683_, _20680_);
  and _71873_ (_20686_, _20685_, _06828_);
  and _71874_ (_20687_, _20600_, _03790_);
  and _71875_ (_20688_, _20687_, _20681_);
  or _71876_ (_20689_, _20688_, _03624_);
  or _71877_ (_20690_, _20689_, _20686_);
  nor _71878_ (_20691_, _13140_, _09236_);
  or _71879_ (_20692_, _20595_, _07795_);
  or _71880_ (_20693_, _20692_, _20691_);
  and _71881_ (_20694_, _20693_, _07793_);
  and _71882_ (_20695_, _20694_, _20690_);
  nor _71883_ (_20696_, _13146_, _09236_);
  or _71884_ (_20697_, _20696_, _20595_);
  and _71885_ (_20698_, _20697_, _03785_);
  or _71886_ (_20699_, _20698_, _03815_);
  or _71887_ (_20700_, _20699_, _20695_);
  or _71888_ (_20701_, _20597_, _04246_);
  and _71889_ (_20702_, _20701_, _03823_);
  and _71890_ (_20703_, _20702_, _20700_);
  and _71891_ (_20704_, _20624_, _03453_);
  or _71892_ (_20706_, _20704_, _03447_);
  or _71893_ (_20707_, _20706_, _20703_);
  and _71894_ (_20708_, _13199_, _05293_);
  or _71895_ (_20709_, _20595_, _03514_);
  or _71896_ (_20710_, _20709_, _20708_);
  and _71897_ (_20711_, _20710_, _43000_);
  and _71898_ (_20712_, _20711_, _20707_);
  or _71899_ (_43539_, _20712_, _20594_);
  not _71900_ (_20713_, \oc8051_golden_model_1.P0 [6]);
  nor _71901_ (_20714_, _05293_, _20713_);
  nor _71902_ (_20716_, _13242_, _09236_);
  or _71903_ (_20717_, _20716_, _20714_);
  or _71904_ (_20718_, _20717_, _04081_);
  and _71905_ (_20719_, _05293_, \oc8051_golden_model_1.ACC [6]);
  or _71906_ (_20720_, _20719_, _20714_);
  and _71907_ (_20721_, _20720_, _04409_);
  nor _71908_ (_20722_, _04409_, _20713_);
  or _71909_ (_20723_, _20722_, _03610_);
  or _71910_ (_20724_, _20723_, _20721_);
  and _71911_ (_20725_, _20724_, _04055_);
  and _71912_ (_20726_, _20725_, _20718_);
  nor _71913_ (_20727_, _05209_, _20713_);
  and _71914_ (_20728_, _13229_, _05209_);
  or _71915_ (_20729_, _20728_, _20727_);
  and _71916_ (_20730_, _20729_, _03715_);
  or _71917_ (_20731_, _20730_, _03723_);
  or _71918_ (_20732_, _20731_, _20726_);
  nor _71919_ (_20733_, _05363_, _09236_);
  or _71920_ (_20734_, _20733_, _20714_);
  or _71921_ (_20735_, _20734_, _03996_);
  and _71922_ (_20737_, _20735_, _20732_);
  or _71923_ (_20738_, _20737_, _03729_);
  or _71924_ (_20739_, _20720_, _03737_);
  and _71925_ (_20740_, _20739_, _03736_);
  and _71926_ (_20741_, _20740_, _20738_);
  and _71927_ (_20742_, _13253_, _05209_);
  or _71928_ (_20743_, _20742_, _20727_);
  and _71929_ (_20744_, _20743_, _03714_);
  or _71930_ (_20745_, _20744_, _03719_);
  or _71931_ (_20746_, _20745_, _20741_);
  or _71932_ (_20748_, _20727_, _13260_);
  and _71933_ (_20749_, _20748_, _20729_);
  or _71934_ (_20750_, _20749_, _06840_);
  and _71935_ (_20751_, _20750_, _03710_);
  and _71936_ (_20752_, _20751_, _20746_);
  or _71937_ (_20753_, _13253_, _13225_);
  and _71938_ (_20754_, _20753_, _05209_);
  or _71939_ (_20755_, _20754_, _20727_);
  and _71940_ (_20756_, _20755_, _03505_);
  or _71941_ (_20757_, _20756_, _07390_);
  or _71942_ (_20758_, _20757_, _20752_);
  or _71943_ (_20759_, _20734_, _06838_);
  and _71944_ (_20760_, _20759_, _20758_);
  or _71945_ (_20761_, _20760_, _04481_);
  and _71946_ (_20762_, _06455_, _05293_);
  or _71947_ (_20763_, _20714_, _07400_);
  or _71948_ (_20764_, _20763_, _20762_);
  and _71949_ (_20765_, _20764_, _03589_);
  and _71950_ (_20766_, _20765_, _20761_);
  and _71951_ (_20767_, _06340_, \oc8051_golden_model_1.P1 [6]);
  and _71952_ (_20769_, _06343_, \oc8051_golden_model_1.P0 [6]);
  and _71953_ (_20770_, _06346_, \oc8051_golden_model_1.P2 [6]);
  and _71954_ (_20771_, _06348_, \oc8051_golden_model_1.P3 [6]);
  or _71955_ (_20772_, _20771_, _20770_);
  or _71956_ (_20773_, _20772_, _20769_);
  nor _71957_ (_20774_, _20773_, _20767_);
  and _71958_ (_20775_, _20774_, _13290_);
  and _71959_ (_20776_, _20775_, _13313_);
  nand _71960_ (_20777_, _20776_, _13329_);
  or _71961_ (_20778_, _20777_, _13287_);
  and _71962_ (_20780_, _20778_, _05293_);
  or _71963_ (_20781_, _20780_, _20714_);
  and _71964_ (_20782_, _20781_, _03222_);
  or _71965_ (_20783_, _20782_, _08828_);
  or _71966_ (_20784_, _20783_, _20766_);
  and _71967_ (_20785_, _13347_, _05293_);
  or _71968_ (_20786_, _20714_, _07766_);
  or _71969_ (_20787_, _20786_, _20785_);
  and _71970_ (_20788_, _13339_, _05293_);
  or _71971_ (_20789_, _20788_, _20714_);
  or _71972_ (_20790_, _20789_, _05886_);
  and _71973_ (_20791_, _20790_, _07778_);
  and _71974_ (_20792_, _20791_, _20787_);
  and _71975_ (_20793_, _20792_, _20784_);
  and _71976_ (_20794_, _13353_, _05293_);
  or _71977_ (_20795_, _20794_, _20714_);
  and _71978_ (_20796_, _20795_, _03780_);
  or _71979_ (_20797_, _20796_, _20793_);
  and _71980_ (_20798_, _20797_, _07777_);
  or _71981_ (_20799_, _20714_, _05412_);
  and _71982_ (_20801_, _20789_, _03622_);
  and _71983_ (_20802_, _20801_, _20799_);
  or _71984_ (_20803_, _20802_, _20798_);
  and _71985_ (_20804_, _20803_, _06828_);
  and _71986_ (_20805_, _20720_, _03790_);
  and _71987_ (_20806_, _20805_, _20799_);
  or _71988_ (_20807_, _20806_, _03624_);
  or _71989_ (_20808_, _20807_, _20804_);
  nor _71990_ (_20809_, _13346_, _09236_);
  or _71991_ (_20810_, _20714_, _07795_);
  or _71992_ (_20812_, _20810_, _20809_);
  and _71993_ (_20813_, _20812_, _07793_);
  and _71994_ (_20814_, _20813_, _20808_);
  nor _71995_ (_20815_, _13352_, _09236_);
  or _71996_ (_20816_, _20815_, _20714_);
  and _71997_ (_20817_, _20816_, _03785_);
  or _71998_ (_20818_, _20817_, _03815_);
  or _71999_ (_20819_, _20818_, _20814_);
  or _72000_ (_20820_, _20717_, _04246_);
  and _72001_ (_20821_, _20820_, _03823_);
  and _72002_ (_20822_, _20821_, _20819_);
  and _72003_ (_20823_, _20743_, _03453_);
  or _72004_ (_20824_, _20823_, _03447_);
  or _72005_ (_20825_, _20824_, _20822_);
  and _72006_ (_20826_, _13402_, _05293_);
  or _72007_ (_20827_, _20714_, _03514_);
  or _72008_ (_20828_, _20827_, _20826_);
  and _72009_ (_20829_, _20828_, _43000_);
  and _72010_ (_20830_, _20829_, _20825_);
  nor _72011_ (_20831_, _43000_, _20713_);
  or _72012_ (_20833_, _20831_, rst);
  or _72013_ (_43540_, _20833_, _20830_);
  not _72014_ (_20834_, \oc8051_golden_model_1.P1 [0]);
  nor _72015_ (_20835_, _43000_, _20834_);
  or _72016_ (_20836_, _20835_, rst);
  nor _72017_ (_20837_, _05266_, _20834_);
  and _72018_ (_20838_, _12128_, _05266_);
  or _72019_ (_20839_, _20838_, _20837_);
  and _72020_ (_20840_, _20839_, _03780_);
  and _72021_ (_20841_, _05266_, _04620_);
  or _72022_ (_20843_, _20841_, _20837_);
  or _72023_ (_20844_, _20843_, _06838_);
  nor _72024_ (_20845_, _05666_, _09352_);
  or _72025_ (_20846_, _20845_, _20837_);
  and _72026_ (_20847_, _20846_, _03610_);
  nor _72027_ (_20848_, _04409_, _20834_);
  and _72028_ (_20849_, _05266_, \oc8051_golden_model_1.ACC [0]);
  or _72029_ (_20850_, _20849_, _20837_);
  and _72030_ (_20851_, _20850_, _04409_);
  or _72031_ (_20852_, _20851_, _20848_);
  and _72032_ (_20853_, _20852_, _04081_);
  or _72033_ (_20854_, _20853_, _03715_);
  or _72034_ (_20855_, _20854_, _20847_);
  and _72035_ (_20856_, _12021_, _05916_);
  nor _72036_ (_20857_, _05916_, _20834_);
  or _72037_ (_20858_, _20857_, _04055_);
  or _72038_ (_20859_, _20858_, _20856_);
  and _72039_ (_20860_, _20859_, _03996_);
  and _72040_ (_20861_, _20860_, _20855_);
  and _72041_ (_20862_, _20843_, _03723_);
  or _72042_ (_20864_, _20862_, _03729_);
  or _72043_ (_20865_, _20864_, _20861_);
  or _72044_ (_20866_, _20850_, _03737_);
  and _72045_ (_20867_, _20866_, _03736_);
  and _72046_ (_20868_, _20867_, _20865_);
  and _72047_ (_20869_, _20837_, _03714_);
  or _72048_ (_20870_, _20869_, _03719_);
  or _72049_ (_20871_, _20870_, _20868_);
  or _72050_ (_20872_, _20846_, _06840_);
  and _72051_ (_20873_, _20872_, _03710_);
  and _72052_ (_20875_, _20873_, _20871_);
  and _72053_ (_20876_, _20023_, _05916_);
  or _72054_ (_20877_, _20876_, _20857_);
  and _72055_ (_20878_, _20877_, _03505_);
  or _72056_ (_20879_, _20878_, _07390_);
  or _72057_ (_20880_, _20879_, _20875_);
  and _72058_ (_20881_, _20880_, _20844_);
  or _72059_ (_20882_, _20881_, _04481_);
  and _72060_ (_20883_, _06546_, _05266_);
  or _72061_ (_20884_, _20837_, _07400_);
  or _72062_ (_20886_, _20884_, _20883_);
  and _72063_ (_20887_, _20886_, _03589_);
  and _72064_ (_20888_, _20887_, _20882_);
  and _72065_ (_20889_, _20049_, _05266_);
  or _72066_ (_20890_, _20889_, _20837_);
  and _72067_ (_20891_, _20890_, _03222_);
  or _72068_ (_20892_, _20891_, _20888_);
  or _72069_ (_20893_, _20892_, _08828_);
  and _72070_ (_20894_, _12124_, _05266_);
  or _72071_ (_20895_, _20837_, _07766_);
  or _72072_ (_20896_, _20895_, _20894_);
  and _72073_ (_20897_, _05266_, _06274_);
  or _72074_ (_20898_, _20897_, _20837_);
  or _72075_ (_20899_, _20898_, _05886_);
  and _72076_ (_20900_, _20899_, _07778_);
  and _72077_ (_20901_, _20900_, _20896_);
  and _72078_ (_20902_, _20901_, _20893_);
  or _72079_ (_20903_, _20902_, _20840_);
  and _72080_ (_20904_, _20903_, _07777_);
  nand _72081_ (_20905_, _20898_, _03622_);
  nor _72082_ (_20907_, _20905_, _20845_);
  or _72083_ (_20908_, _20907_, _20904_);
  and _72084_ (_20909_, _20908_, _06828_);
  or _72085_ (_20910_, _20837_, _05666_);
  and _72086_ (_20911_, _20850_, _03790_);
  and _72087_ (_20912_, _20911_, _20910_);
  or _72088_ (_20913_, _20912_, _03624_);
  or _72089_ (_20914_, _20913_, _20909_);
  nor _72090_ (_20915_, _12122_, _09352_);
  or _72091_ (_20916_, _20837_, _07795_);
  or _72092_ (_20918_, _20916_, _20915_);
  and _72093_ (_20919_, _20918_, _07793_);
  and _72094_ (_20920_, _20919_, _20914_);
  nor _72095_ (_20921_, _12003_, _09352_);
  or _72096_ (_20922_, _20921_, _20837_);
  and _72097_ (_20923_, _20922_, _03785_);
  or _72098_ (_20924_, _20923_, _03815_);
  or _72099_ (_20925_, _20924_, _20920_);
  or _72100_ (_20926_, _20846_, _04246_);
  and _72101_ (_20927_, _20926_, _03823_);
  and _72102_ (_20928_, _20927_, _20925_);
  and _72103_ (_20929_, _20837_, _03453_);
  or _72104_ (_20930_, _20929_, _03447_);
  or _72105_ (_20931_, _20930_, _20928_);
  or _72106_ (_20932_, _20846_, _03514_);
  and _72107_ (_20933_, _20932_, _43000_);
  and _72108_ (_20934_, _20933_, _20931_);
  or _72109_ (_43543_, _20934_, _20836_);
  or _72110_ (_20935_, _05266_, \oc8051_golden_model_1.P1 [1]);
  and _72111_ (_20936_, _12213_, _05266_);
  not _72112_ (_20938_, _20936_);
  and _72113_ (_20939_, _20938_, _20935_);
  or _72114_ (_20940_, _20939_, _04081_);
  nand _72115_ (_20941_, _05266_, _03274_);
  and _72116_ (_20942_, _20941_, _20935_);
  and _72117_ (_20943_, _20942_, _04409_);
  not _72118_ (_20944_, \oc8051_golden_model_1.P1 [1]);
  nor _72119_ (_20945_, _04409_, _20944_);
  or _72120_ (_20946_, _20945_, _03610_);
  or _72121_ (_20947_, _20946_, _20943_);
  and _72122_ (_20949_, _20947_, _04055_);
  and _72123_ (_20950_, _20949_, _20940_);
  and _72124_ (_20951_, _12224_, _05916_);
  nor _72125_ (_20952_, _05916_, _20944_);
  or _72126_ (_20953_, _20952_, _03723_);
  or _72127_ (_20954_, _20953_, _20951_);
  and _72128_ (_20955_, _20954_, _14265_);
  or _72129_ (_20956_, _20955_, _20950_);
  nor _72130_ (_20957_, _05266_, _20944_);
  and _72131_ (_20958_, _05266_, _06764_);
  or _72132_ (_20960_, _20958_, _20957_);
  or _72133_ (_20961_, _20960_, _03996_);
  and _72134_ (_20962_, _20961_, _20956_);
  or _72135_ (_20963_, _20962_, _03729_);
  or _72136_ (_20964_, _20942_, _03737_);
  and _72137_ (_20965_, _20964_, _03736_);
  and _72138_ (_20966_, _20965_, _20963_);
  and _72139_ (_20967_, _12211_, _05916_);
  or _72140_ (_20968_, _20967_, _20952_);
  and _72141_ (_20969_, _20968_, _03714_);
  or _72142_ (_20970_, _20969_, _03719_);
  or _72143_ (_20971_, _20970_, _20966_);
  and _72144_ (_20972_, _20951_, _12239_);
  or _72145_ (_20973_, _20952_, _06840_);
  or _72146_ (_20974_, _20973_, _20972_);
  and _72147_ (_20975_, _20974_, _20971_);
  and _72148_ (_20976_, _20975_, _03710_);
  and _72149_ (_20977_, _20141_, _05916_);
  or _72150_ (_20978_, _20952_, _20977_);
  and _72151_ (_20979_, _20978_, _03505_);
  or _72152_ (_20981_, _20979_, _07390_);
  or _72153_ (_20982_, _20981_, _20976_);
  or _72154_ (_20983_, _20960_, _06838_);
  and _72155_ (_20984_, _20983_, _20982_);
  or _72156_ (_20985_, _20984_, _04481_);
  and _72157_ (_20986_, _06501_, _05266_);
  or _72158_ (_20987_, _20957_, _07400_);
  or _72159_ (_20988_, _20987_, _20986_);
  and _72160_ (_20989_, _20988_, _03589_);
  and _72161_ (_20990_, _20989_, _20985_);
  and _72162_ (_20992_, _20168_, _05266_);
  or _72163_ (_20993_, _20992_, _20957_);
  and _72164_ (_20994_, _20993_, _03222_);
  or _72165_ (_20995_, _20994_, _20990_);
  and _72166_ (_20996_, _20995_, _03602_);
  or _72167_ (_20997_, _12327_, _09352_);
  and _72168_ (_20998_, _20997_, _03600_);
  nand _72169_ (_20999_, _05266_, _04303_);
  and _72170_ (_21000_, _20999_, _03601_);
  or _72171_ (_21001_, _21000_, _20998_);
  and _72172_ (_21002_, _21001_, _20935_);
  or _72173_ (_21003_, _21002_, _20996_);
  and _72174_ (_21004_, _21003_, _07778_);
  or _72175_ (_21005_, _12333_, _09352_);
  and _72176_ (_21006_, _20935_, _03780_);
  and _72177_ (_21007_, _21006_, _21005_);
  or _72178_ (_21008_, _21007_, _21004_);
  and _72179_ (_21009_, _21008_, _07777_);
  or _72180_ (_21010_, _12207_, _09352_);
  and _72181_ (_21011_, _20935_, _03622_);
  and _72182_ (_21013_, _21011_, _21010_);
  or _72183_ (_21014_, _21013_, _21009_);
  and _72184_ (_21015_, _21014_, _06828_);
  or _72185_ (_21016_, _20957_, _05618_);
  and _72186_ (_21017_, _20942_, _03790_);
  and _72187_ (_21018_, _21017_, _21016_);
  or _72188_ (_21019_, _21018_, _21015_);
  and _72189_ (_21020_, _21019_, _03786_);
  or _72190_ (_21021_, _20999_, _05618_);
  and _72191_ (_21022_, _20935_, _03624_);
  and _72192_ (_21024_, _21022_, _21021_);
  or _72193_ (_21025_, _20941_, _05618_);
  and _72194_ (_21026_, _20935_, _03785_);
  and _72195_ (_21027_, _21026_, _21025_);
  or _72196_ (_21028_, _21027_, _03815_);
  or _72197_ (_21029_, _21028_, _21024_);
  or _72198_ (_21030_, _21029_, _21020_);
  or _72199_ (_21031_, _20939_, _04246_);
  and _72200_ (_21032_, _21031_, _03823_);
  and _72201_ (_21033_, _21032_, _21030_);
  and _72202_ (_21035_, _20968_, _03453_);
  or _72203_ (_21036_, _21035_, _03447_);
  or _72204_ (_21037_, _21036_, _21033_);
  or _72205_ (_21038_, _20957_, _03514_);
  or _72206_ (_21039_, _21038_, _20936_);
  and _72207_ (_21040_, _21039_, _43000_);
  and _72208_ (_21041_, _21040_, _21037_);
  nor _72209_ (_21042_, _43000_, _20944_);
  or _72210_ (_21043_, _21042_, rst);
  or _72211_ (_43544_, _21043_, _21041_);
  not _72212_ (_21045_, \oc8051_golden_model_1.P1 [2]);
  nor _72213_ (_21046_, _43000_, _21045_);
  or _72214_ (_21047_, _21046_, rst);
  nor _72215_ (_21048_, _05266_, _21045_);
  nor _72216_ (_21049_, _09352_, _04875_);
  or _72217_ (_21050_, _21049_, _21048_);
  or _72218_ (_21051_, _21050_, _06838_);
  or _72219_ (_21052_, _21050_, _03996_);
  nor _72220_ (_21053_, _12416_, _09352_);
  or _72221_ (_21054_, _21053_, _21048_);
  or _72222_ (_21056_, _21054_, _04081_);
  and _72223_ (_21057_, _05266_, \oc8051_golden_model_1.ACC [2]);
  or _72224_ (_21058_, _21057_, _21048_);
  and _72225_ (_21059_, _21058_, _04409_);
  nor _72226_ (_21060_, _04409_, _21045_);
  or _72227_ (_21061_, _21060_, _03610_);
  or _72228_ (_21062_, _21061_, _21059_);
  and _72229_ (_21063_, _21062_, _04055_);
  and _72230_ (_21064_, _21063_, _21056_);
  nor _72231_ (_21065_, _05916_, _21045_);
  and _72232_ (_21067_, _12411_, _05916_);
  or _72233_ (_21068_, _21067_, _21065_);
  and _72234_ (_21069_, _21068_, _03715_);
  or _72235_ (_21070_, _21069_, _03723_);
  or _72236_ (_21071_, _21070_, _21064_);
  and _72237_ (_21072_, _21071_, _21052_);
  or _72238_ (_21073_, _21072_, _03729_);
  or _72239_ (_21074_, _21058_, _03737_);
  and _72240_ (_21075_, _21074_, _03736_);
  and _72241_ (_21076_, _21075_, _21073_);
  and _72242_ (_21078_, _12409_, _05916_);
  or _72243_ (_21079_, _21078_, _21065_);
  and _72244_ (_21080_, _21079_, _03714_);
  or _72245_ (_21081_, _21080_, _03719_);
  or _72246_ (_21082_, _21081_, _21076_);
  and _72247_ (_21083_, _21067_, _12443_);
  or _72248_ (_21084_, _21065_, _06840_);
  or _72249_ (_21085_, _21084_, _21083_);
  and _72250_ (_21086_, _21085_, _03710_);
  and _72251_ (_21087_, _21086_, _21082_);
  and _72252_ (_21089_, _20264_, _05916_);
  or _72253_ (_21090_, _21089_, _21065_);
  and _72254_ (_21091_, _21090_, _03505_);
  or _72255_ (_21092_, _21091_, _07390_);
  or _72256_ (_21093_, _21092_, _21087_);
  and _72257_ (_21094_, _21093_, _21051_);
  or _72258_ (_21095_, _21094_, _04481_);
  and _72259_ (_21096_, _06637_, _05266_);
  or _72260_ (_21097_, _21048_, _07400_);
  or _72261_ (_21098_, _21097_, _21096_);
  and _72262_ (_21100_, _21098_, _03589_);
  and _72263_ (_21101_, _21100_, _21095_);
  and _72264_ (_21102_, _20290_, _05266_);
  or _72265_ (_21103_, _21048_, _21102_);
  and _72266_ (_21104_, _21103_, _03222_);
  or _72267_ (_21105_, _21104_, _21101_);
  or _72268_ (_21106_, _21105_, _08828_);
  and _72269_ (_21107_, _12533_, _05266_);
  or _72270_ (_21108_, _21048_, _07766_);
  or _72271_ (_21109_, _21108_, _21107_);
  and _72272_ (_21110_, _05266_, _06332_);
  or _72273_ (_21111_, _21110_, _21048_);
  or _72274_ (_21112_, _21111_, _05886_);
  and _72275_ (_21113_, _21112_, _07778_);
  and _72276_ (_21114_, _21113_, _21109_);
  and _72277_ (_21115_, _21114_, _21106_);
  and _72278_ (_21116_, _12539_, _05266_);
  or _72279_ (_21117_, _21116_, _21048_);
  and _72280_ (_21118_, _21117_, _03780_);
  or _72281_ (_21119_, _21118_, _21115_);
  and _72282_ (_21120_, _21119_, _07777_);
  or _72283_ (_21121_, _21048_, _05718_);
  and _72284_ (_21122_, _21111_, _03622_);
  and _72285_ (_21123_, _21122_, _21121_);
  or _72286_ (_21124_, _21123_, _21120_);
  and _72287_ (_21125_, _21124_, _06828_);
  and _72288_ (_21126_, _21058_, _03790_);
  and _72289_ (_21127_, _21126_, _21121_);
  or _72290_ (_21128_, _21127_, _03624_);
  or _72291_ (_21129_, _21128_, _21125_);
  nor _72292_ (_21131_, _12532_, _09352_);
  or _72293_ (_21132_, _21048_, _07795_);
  or _72294_ (_21133_, _21132_, _21131_);
  and _72295_ (_21134_, _21133_, _07793_);
  and _72296_ (_21135_, _21134_, _21129_);
  nor _72297_ (_21136_, _12538_, _09352_);
  or _72298_ (_21137_, _21136_, _21048_);
  and _72299_ (_21138_, _21137_, _03785_);
  or _72300_ (_21139_, _21138_, _03815_);
  or _72301_ (_21140_, _21139_, _21135_);
  or _72302_ (_21142_, _21054_, _04246_);
  and _72303_ (_21143_, _21142_, _03823_);
  and _72304_ (_21144_, _21143_, _21140_);
  and _72305_ (_21145_, _21079_, _03453_);
  or _72306_ (_21146_, _21145_, _03447_);
  or _72307_ (_21147_, _21146_, _21144_);
  and _72308_ (_21148_, _12592_, _05266_);
  or _72309_ (_21149_, _21048_, _03514_);
  or _72310_ (_21150_, _21149_, _21148_);
  and _72311_ (_21151_, _21150_, _43000_);
  and _72312_ (_21153_, _21151_, _21147_);
  or _72313_ (_43545_, _21153_, _21047_);
  and _72314_ (_21154_, _09352_, \oc8051_golden_model_1.P1 [3]);
  nor _72315_ (_21155_, _09352_, _05005_);
  or _72316_ (_21156_, _21155_, _21154_);
  or _72317_ (_21157_, _21156_, _06838_);
  nor _72318_ (_21158_, _12627_, _09352_);
  or _72319_ (_21159_, _21158_, _21154_);
  or _72320_ (_21160_, _21159_, _04081_);
  and _72321_ (_21161_, _05266_, \oc8051_golden_model_1.ACC [3]);
  or _72322_ (_21163_, _21161_, _21154_);
  and _72323_ (_21164_, _21163_, _04409_);
  and _72324_ (_21165_, _09029_, \oc8051_golden_model_1.P1 [3]);
  or _72325_ (_21166_, _21165_, _03610_);
  or _72326_ (_21167_, _21166_, _21164_);
  and _72327_ (_21168_, _21167_, _04055_);
  and _72328_ (_21169_, _21168_, _21160_);
  not _72329_ (_21170_, _05916_);
  and _72330_ (_21171_, _21170_, \oc8051_golden_model_1.P1 [3]);
  and _72331_ (_21172_, _12631_, _05916_);
  or _72332_ (_21174_, _21172_, _21171_);
  and _72333_ (_21175_, _21174_, _03715_);
  or _72334_ (_21176_, _21175_, _03723_);
  or _72335_ (_21177_, _21176_, _21169_);
  or _72336_ (_21178_, _21156_, _03996_);
  and _72337_ (_21179_, _21178_, _21177_);
  or _72338_ (_21180_, _21179_, _03729_);
  or _72339_ (_21181_, _21163_, _03737_);
  and _72340_ (_21182_, _21181_, _03736_);
  and _72341_ (_21183_, _21182_, _21180_);
  and _72342_ (_21185_, _12641_, _05916_);
  or _72343_ (_21186_, _21185_, _21171_);
  and _72344_ (_21187_, _21186_, _03714_);
  or _72345_ (_21188_, _21187_, _03719_);
  or _72346_ (_21189_, _21188_, _21183_);
  or _72347_ (_21190_, _21171_, _12648_);
  and _72348_ (_21191_, _21190_, _21174_);
  or _72349_ (_21192_, _21191_, _06840_);
  and _72350_ (_21193_, _21192_, _03710_);
  and _72351_ (_21194_, _21193_, _21189_);
  and _72352_ (_21196_, _20391_, _05916_);
  or _72353_ (_21197_, _21196_, _21171_);
  and _72354_ (_21198_, _21197_, _03505_);
  or _72355_ (_21199_, _21198_, _07390_);
  or _72356_ (_21200_, _21199_, _21194_);
  and _72357_ (_21201_, _21200_, _21157_);
  or _72358_ (_21202_, _21201_, _04481_);
  and _72359_ (_21203_, _06592_, _05266_);
  or _72360_ (_21204_, _21154_, _07400_);
  or _72361_ (_21205_, _21204_, _21203_);
  and _72362_ (_21207_, _21205_, _03589_);
  and _72363_ (_21208_, _21207_, _21202_);
  and _72364_ (_21209_, _20416_, _05266_);
  or _72365_ (_21210_, _21154_, _21209_);
  and _72366_ (_21211_, _21210_, _03222_);
  or _72367_ (_21212_, _21211_, _21208_);
  or _72368_ (_21213_, _21212_, _08828_);
  and _72369_ (_21214_, _12733_, _05266_);
  or _72370_ (_21215_, _21154_, _07766_);
  or _72371_ (_21216_, _21215_, _21214_);
  and _72372_ (_21218_, _05266_, _06276_);
  or _72373_ (_21219_, _21218_, _21154_);
  or _72374_ (_21220_, _21219_, _05886_);
  and _72375_ (_21221_, _21220_, _07778_);
  and _72376_ (_21222_, _21221_, _21216_);
  and _72377_ (_21223_, _21222_, _21213_);
  and _72378_ (_21224_, _12739_, _05266_);
  or _72379_ (_21225_, _21224_, _21154_);
  and _72380_ (_21226_, _21225_, _03780_);
  or _72381_ (_21227_, _21226_, _21223_);
  and _72382_ (_21229_, _21227_, _07777_);
  or _72383_ (_21230_, _21154_, _05567_);
  and _72384_ (_21231_, _21219_, _03622_);
  and _72385_ (_21232_, _21231_, _21230_);
  or _72386_ (_21233_, _21232_, _21229_);
  and _72387_ (_21234_, _21233_, _06828_);
  and _72388_ (_21235_, _21163_, _03790_);
  and _72389_ (_21236_, _21235_, _21230_);
  or _72390_ (_21237_, _21236_, _03624_);
  or _72391_ (_21238_, _21237_, _21234_);
  nor _72392_ (_21240_, _12732_, _09352_);
  or _72393_ (_21241_, _21154_, _07795_);
  or _72394_ (_21242_, _21241_, _21240_);
  and _72395_ (_21243_, _21242_, _07793_);
  and _72396_ (_21244_, _21243_, _21238_);
  nor _72397_ (_21245_, _12738_, _09352_);
  or _72398_ (_21246_, _21245_, _21154_);
  and _72399_ (_21247_, _21246_, _03785_);
  or _72400_ (_21248_, _21247_, _03815_);
  or _72401_ (_21249_, _21248_, _21244_);
  or _72402_ (_21251_, _21159_, _04246_);
  and _72403_ (_21252_, _21251_, _03823_);
  and _72404_ (_21253_, _21252_, _21249_);
  and _72405_ (_21254_, _21186_, _03453_);
  or _72406_ (_21255_, _21254_, _03447_);
  or _72407_ (_21256_, _21255_, _21253_);
  and _72408_ (_21257_, _12794_, _05266_);
  or _72409_ (_21258_, _21154_, _03514_);
  or _72410_ (_21259_, _21258_, _21257_);
  and _72411_ (_21260_, _21259_, _43000_);
  and _72412_ (_21262_, _21260_, _21256_);
  nor _72413_ (_21263_, \oc8051_golden_model_1.P1 [3], rst);
  nor _72414_ (_21264_, _21263_, _04794_);
  or _72415_ (_43546_, _21264_, _21262_);
  nor _72416_ (_21265_, \oc8051_golden_model_1.P1 [4], rst);
  nor _72417_ (_21266_, _21265_, _04794_);
  and _72418_ (_21267_, _09352_, \oc8051_golden_model_1.P1 [4]);
  nor _72419_ (_21268_, _05777_, _09352_);
  or _72420_ (_21269_, _21268_, _21267_);
  or _72421_ (_21270_, _21269_, _06838_);
  and _72422_ (_21272_, _21170_, \oc8051_golden_model_1.P1 [4]);
  and _72423_ (_21273_, _12827_, _05916_);
  or _72424_ (_21274_, _21273_, _21272_);
  and _72425_ (_21275_, _21274_, _03714_);
  nor _72426_ (_21276_, _12841_, _09352_);
  or _72427_ (_21277_, _21276_, _21267_);
  or _72428_ (_21278_, _21277_, _04081_);
  and _72429_ (_21279_, _05266_, \oc8051_golden_model_1.ACC [4]);
  or _72430_ (_21280_, _21279_, _21267_);
  and _72431_ (_21281_, _21280_, _04409_);
  and _72432_ (_21283_, _09029_, \oc8051_golden_model_1.P1 [4]);
  or _72433_ (_21284_, _21283_, _03610_);
  or _72434_ (_21285_, _21284_, _21281_);
  and _72435_ (_21286_, _21285_, _04055_);
  and _72436_ (_21287_, _21286_, _21278_);
  and _72437_ (_21288_, _12845_, _05916_);
  or _72438_ (_21289_, _21288_, _21272_);
  and _72439_ (_21290_, _21289_, _03715_);
  or _72440_ (_21291_, _21290_, _03723_);
  or _72441_ (_21292_, _21291_, _21287_);
  or _72442_ (_21294_, _21269_, _03996_);
  and _72443_ (_21295_, _21294_, _21292_);
  or _72444_ (_21296_, _21295_, _03729_);
  or _72445_ (_21297_, _21280_, _03737_);
  and _72446_ (_21298_, _21297_, _03736_);
  and _72447_ (_21299_, _21298_, _21296_);
  or _72448_ (_21300_, _21299_, _21275_);
  and _72449_ (_21301_, _21300_, _06840_);
  and _72450_ (_21302_, _12861_, _05916_);
  or _72451_ (_21303_, _21302_, _21272_);
  and _72452_ (_21305_, _21303_, _03719_);
  or _72453_ (_21306_, _21305_, _21301_);
  and _72454_ (_21307_, _21306_, _03710_);
  and _72455_ (_21308_, _20511_, _05916_);
  or _72456_ (_21309_, _21308_, _21272_);
  and _72457_ (_21310_, _21309_, _03505_);
  or _72458_ (_21311_, _21310_, _07390_);
  or _72459_ (_21312_, _21311_, _21307_);
  and _72460_ (_21313_, _21312_, _21270_);
  or _72461_ (_21314_, _21313_, _04481_);
  and _72462_ (_21316_, _06730_, _05266_);
  or _72463_ (_21317_, _21267_, _07400_);
  or _72464_ (_21318_, _21317_, _21316_);
  and _72465_ (_21319_, _21318_, _03589_);
  and _72466_ (_21320_, _21319_, _21314_);
  and _72467_ (_21321_, _20536_, _05266_);
  or _72468_ (_21322_, _21321_, _21267_);
  and _72469_ (_21323_, _21322_, _03222_);
  or _72470_ (_21324_, _21323_, _08828_);
  or _72471_ (_21325_, _21324_, _21320_);
  and _72472_ (_21327_, _12821_, _05266_);
  or _72473_ (_21328_, _21267_, _07766_);
  or _72474_ (_21329_, _21328_, _21327_);
  and _72475_ (_21330_, _06298_, _05266_);
  or _72476_ (_21331_, _21330_, _21267_);
  or _72477_ (_21332_, _21331_, _05886_);
  and _72478_ (_21333_, _21332_, _07778_);
  and _72479_ (_21334_, _21333_, _21329_);
  and _72480_ (_21335_, _21334_, _21325_);
  and _72481_ (_21336_, _12817_, _05266_);
  or _72482_ (_21338_, _21336_, _21267_);
  and _72483_ (_21339_, _21338_, _03780_);
  or _72484_ (_21340_, _21339_, _21335_);
  and _72485_ (_21341_, _21340_, _07777_);
  or _72486_ (_21342_, _21267_, _05825_);
  and _72487_ (_21343_, _21331_, _03622_);
  and _72488_ (_21344_, _21343_, _21342_);
  or _72489_ (_21345_, _21344_, _21341_);
  and _72490_ (_21346_, _21345_, _06828_);
  and _72491_ (_21347_, _21280_, _03790_);
  and _72492_ (_21349_, _21347_, _21342_);
  or _72493_ (_21350_, _21349_, _03624_);
  or _72494_ (_21351_, _21350_, _21346_);
  nor _72495_ (_21352_, _12819_, _09352_);
  or _72496_ (_21353_, _21267_, _07795_);
  or _72497_ (_21354_, _21353_, _21352_);
  and _72498_ (_21355_, _21354_, _07793_);
  and _72499_ (_21356_, _21355_, _21351_);
  nor _72500_ (_21357_, _12816_, _09352_);
  or _72501_ (_21358_, _21357_, _21267_);
  and _72502_ (_21360_, _21358_, _03785_);
  or _72503_ (_21361_, _21360_, _03815_);
  or _72504_ (_21362_, _21361_, _21356_);
  or _72505_ (_21363_, _21277_, _04246_);
  and _72506_ (_21364_, _21363_, _03823_);
  and _72507_ (_21365_, _21364_, _21362_);
  and _72508_ (_21366_, _21274_, _03453_);
  or _72509_ (_21367_, _21366_, _03447_);
  or _72510_ (_21368_, _21367_, _21365_);
  and _72511_ (_21369_, _13003_, _05266_);
  or _72512_ (_21371_, _21267_, _03514_);
  or _72513_ (_21372_, _21371_, _21369_);
  and _72514_ (_21373_, _21372_, _43000_);
  and _72515_ (_21374_, _21373_, _21368_);
  or _72516_ (_43547_, _21374_, _21266_);
  nor _72517_ (_21375_, \oc8051_golden_model_1.P1 [5], rst);
  nor _72518_ (_21376_, _21375_, _04794_);
  and _72519_ (_21377_, _09352_, \oc8051_golden_model_1.P1 [5]);
  nor _72520_ (_21378_, _13014_, _09352_);
  or _72521_ (_21379_, _21378_, _21377_);
  or _72522_ (_21381_, _21379_, _04081_);
  and _72523_ (_21382_, _05266_, \oc8051_golden_model_1.ACC [5]);
  or _72524_ (_21383_, _21382_, _21377_);
  and _72525_ (_21384_, _21383_, _04409_);
  and _72526_ (_21385_, _09029_, \oc8051_golden_model_1.P1 [5]);
  or _72527_ (_21386_, _21385_, _03610_);
  or _72528_ (_21387_, _21386_, _21384_);
  and _72529_ (_21388_, _21387_, _04055_);
  and _72530_ (_21389_, _21388_, _21381_);
  and _72531_ (_21390_, _21170_, \oc8051_golden_model_1.P1 [5]);
  and _72532_ (_21392_, _13037_, _05916_);
  or _72533_ (_21393_, _21392_, _21390_);
  and _72534_ (_21394_, _21393_, _03715_);
  or _72535_ (_21395_, _21394_, _03723_);
  or _72536_ (_21396_, _21395_, _21389_);
  nor _72537_ (_21397_, _05469_, _09352_);
  or _72538_ (_21398_, _21397_, _21377_);
  or _72539_ (_21399_, _21398_, _03996_);
  and _72540_ (_21400_, _21399_, _21396_);
  or _72541_ (_21401_, _21400_, _03729_);
  or _72542_ (_21403_, _21383_, _03737_);
  and _72543_ (_21404_, _21403_, _03736_);
  and _72544_ (_21405_, _21404_, _21401_);
  and _72545_ (_21406_, _13047_, _05916_);
  or _72546_ (_21407_, _21406_, _21390_);
  and _72547_ (_21408_, _21407_, _03714_);
  or _72548_ (_21409_, _21408_, _03719_);
  or _72549_ (_21410_, _21409_, _21405_);
  or _72550_ (_21411_, _21390_, _13054_);
  and _72551_ (_21412_, _21411_, _21393_);
  or _72552_ (_21414_, _21412_, _06840_);
  and _72553_ (_21415_, _21414_, _03710_);
  and _72554_ (_21416_, _21415_, _21410_);
  and _72555_ (_21417_, _20633_, _05916_);
  or _72556_ (_21418_, _21417_, _21390_);
  and _72557_ (_21419_, _21418_, _03505_);
  or _72558_ (_21420_, _21419_, _07390_);
  or _72559_ (_21421_, _21420_, _21416_);
  or _72560_ (_21422_, _21398_, _06838_);
  and _72561_ (_21423_, _21422_, _21421_);
  or _72562_ (_21425_, _21423_, _04481_);
  and _72563_ (_21426_, _06684_, _05266_);
  or _72564_ (_21427_, _21377_, _07400_);
  or _72565_ (_21428_, _21427_, _21426_);
  and _72566_ (_21429_, _21428_, _03589_);
  and _72567_ (_21430_, _21429_, _21425_);
  and _72568_ (_21431_, _20660_, _05266_);
  or _72569_ (_21432_, _21431_, _21377_);
  and _72570_ (_21433_, _21432_, _03222_);
  or _72571_ (_21434_, _21433_, _08828_);
  or _72572_ (_21436_, _21434_, _21430_);
  and _72573_ (_21437_, _13141_, _05266_);
  or _72574_ (_21438_, _21377_, _07766_);
  or _72575_ (_21439_, _21438_, _21437_);
  and _72576_ (_21440_, _06306_, _05266_);
  or _72577_ (_21441_, _21440_, _21377_);
  or _72578_ (_21442_, _21441_, _05886_);
  and _72579_ (_21443_, _21442_, _07778_);
  and _72580_ (_21444_, _21443_, _21439_);
  and _72581_ (_21445_, _21444_, _21436_);
  and _72582_ (_21447_, _13147_, _05266_);
  or _72583_ (_21448_, _21447_, _21377_);
  and _72584_ (_21449_, _21448_, _03780_);
  or _72585_ (_21450_, _21449_, _21445_);
  and _72586_ (_21451_, _21450_, _07777_);
  or _72587_ (_21452_, _21377_, _05518_);
  and _72588_ (_21453_, _21441_, _03622_);
  and _72589_ (_21454_, _21453_, _21452_);
  or _72590_ (_21455_, _21454_, _21451_);
  and _72591_ (_21456_, _21455_, _06828_);
  and _72592_ (_21458_, _21383_, _03790_);
  and _72593_ (_21459_, _21458_, _21452_);
  or _72594_ (_21460_, _21459_, _03624_);
  or _72595_ (_21461_, _21460_, _21456_);
  nor _72596_ (_21462_, _13140_, _09352_);
  or _72597_ (_21463_, _21377_, _07795_);
  or _72598_ (_21464_, _21463_, _21462_);
  and _72599_ (_21465_, _21464_, _07793_);
  and _72600_ (_21466_, _21465_, _21461_);
  nor _72601_ (_21467_, _13146_, _09352_);
  or _72602_ (_21469_, _21467_, _21377_);
  and _72603_ (_21470_, _21469_, _03785_);
  or _72604_ (_21471_, _21470_, _03815_);
  or _72605_ (_21472_, _21471_, _21466_);
  or _72606_ (_21473_, _21379_, _04246_);
  and _72607_ (_21474_, _21473_, _03823_);
  and _72608_ (_21475_, _21474_, _21472_);
  and _72609_ (_21476_, _21407_, _03453_);
  or _72610_ (_21477_, _21476_, _03447_);
  or _72611_ (_21478_, _21477_, _21475_);
  and _72612_ (_21480_, _13199_, _05266_);
  or _72613_ (_21481_, _21377_, _03514_);
  or _72614_ (_21482_, _21481_, _21480_);
  and _72615_ (_21483_, _21482_, _43000_);
  and _72616_ (_21484_, _21483_, _21478_);
  or _72617_ (_43550_, _21484_, _21376_);
  not _72618_ (_21485_, \oc8051_golden_model_1.P1 [6]);
  nor _72619_ (_21486_, _05266_, _21485_);
  nor _72620_ (_21487_, _13242_, _09352_);
  or _72621_ (_21488_, _21487_, _21486_);
  or _72622_ (_21491_, _21488_, _04081_);
  and _72623_ (_21492_, _05266_, \oc8051_golden_model_1.ACC [6]);
  or _72624_ (_21493_, _21492_, _21486_);
  and _72625_ (_21494_, _21493_, _04409_);
  nor _72626_ (_21495_, _04409_, _21485_);
  or _72627_ (_21496_, _21495_, _03610_);
  or _72628_ (_21497_, _21496_, _21494_);
  and _72629_ (_21498_, _21497_, _04055_);
  and _72630_ (_21499_, _21498_, _21491_);
  nor _72631_ (_21500_, _05916_, _21485_);
  and _72632_ (_21503_, _13229_, _05916_);
  or _72633_ (_21504_, _21503_, _21500_);
  and _72634_ (_21505_, _21504_, _03715_);
  or _72635_ (_21506_, _21505_, _03723_);
  or _72636_ (_21507_, _21506_, _21499_);
  nor _72637_ (_21508_, _05363_, _09352_);
  or _72638_ (_21509_, _21508_, _21486_);
  or _72639_ (_21510_, _21509_, _03996_);
  and _72640_ (_21511_, _21510_, _21507_);
  or _72641_ (_21512_, _21511_, _03729_);
  or _72642_ (_21515_, _21493_, _03737_);
  and _72643_ (_21516_, _21515_, _03736_);
  and _72644_ (_21517_, _21516_, _21512_);
  and _72645_ (_21518_, _13253_, _05916_);
  or _72646_ (_21519_, _21518_, _21500_);
  and _72647_ (_21520_, _21519_, _03714_);
  or _72648_ (_21521_, _21520_, _03719_);
  or _72649_ (_21522_, _21521_, _21517_);
  or _72650_ (_21523_, _21500_, _13260_);
  and _72651_ (_21524_, _21523_, _21504_);
  or _72652_ (_21527_, _21524_, _06840_);
  and _72653_ (_21528_, _21527_, _03710_);
  and _72654_ (_21529_, _21528_, _21522_);
  and _72655_ (_21530_, _20753_, _05916_);
  or _72656_ (_21531_, _21530_, _21500_);
  and _72657_ (_21532_, _21531_, _03505_);
  or _72658_ (_21533_, _21532_, _07390_);
  or _72659_ (_21534_, _21533_, _21529_);
  or _72660_ (_21535_, _21509_, _06838_);
  and _72661_ (_21536_, _21535_, _21534_);
  or _72662_ (_21539_, _21536_, _04481_);
  and _72663_ (_21540_, _06455_, _05266_);
  or _72664_ (_21541_, _21486_, _07400_);
  or _72665_ (_21542_, _21541_, _21540_);
  and _72666_ (_21543_, _21542_, _03589_);
  and _72667_ (_21544_, _21543_, _21539_);
  and _72668_ (_21545_, _20778_, _05266_);
  or _72669_ (_21546_, _21545_, _21486_);
  and _72670_ (_21547_, _21546_, _03222_);
  or _72671_ (_21548_, _21547_, _08828_);
  or _72672_ (_21551_, _21548_, _21544_);
  and _72673_ (_21552_, _13347_, _05266_);
  or _72674_ (_21553_, _21486_, _07766_);
  or _72675_ (_21554_, _21553_, _21552_);
  and _72676_ (_21555_, _13339_, _05266_);
  or _72677_ (_21556_, _21555_, _21486_);
  or _72678_ (_21557_, _21556_, _05886_);
  and _72679_ (_21558_, _21557_, _07778_);
  and _72680_ (_21559_, _21558_, _21554_);
  and _72681_ (_21560_, _21559_, _21551_);
  and _72682_ (_21562_, _13353_, _05266_);
  or _72683_ (_21563_, _21562_, _21486_);
  and _72684_ (_21564_, _21563_, _03780_);
  or _72685_ (_21565_, _21564_, _21560_);
  and _72686_ (_21566_, _21565_, _07777_);
  or _72687_ (_21567_, _21486_, _05412_);
  and _72688_ (_21568_, _21556_, _03622_);
  and _72689_ (_21569_, _21568_, _21567_);
  or _72690_ (_21570_, _21569_, _21566_);
  and _72691_ (_21571_, _21570_, _06828_);
  and _72692_ (_21573_, _21493_, _03790_);
  and _72693_ (_21574_, _21573_, _21567_);
  or _72694_ (_21575_, _21574_, _03624_);
  or _72695_ (_21576_, _21575_, _21571_);
  nor _72696_ (_21577_, _13346_, _09352_);
  or _72697_ (_21578_, _21486_, _07795_);
  or _72698_ (_21579_, _21578_, _21577_);
  and _72699_ (_21580_, _21579_, _07793_);
  and _72700_ (_21581_, _21580_, _21576_);
  nor _72701_ (_21582_, _13352_, _09352_);
  or _72702_ (_21584_, _21582_, _21486_);
  and _72703_ (_21585_, _21584_, _03785_);
  or _72704_ (_21586_, _21585_, _03815_);
  or _72705_ (_21587_, _21586_, _21581_);
  or _72706_ (_21588_, _21488_, _04246_);
  and _72707_ (_21589_, _21588_, _03823_);
  and _72708_ (_21590_, _21589_, _21587_);
  and _72709_ (_21591_, _21519_, _03453_);
  or _72710_ (_21592_, _21591_, _03447_);
  or _72711_ (_21593_, _21592_, _21590_);
  and _72712_ (_21595_, _13402_, _05266_);
  or _72713_ (_21596_, _21486_, _03514_);
  or _72714_ (_21597_, _21596_, _21595_);
  and _72715_ (_21598_, _21597_, _43000_);
  and _72716_ (_21599_, _21598_, _21593_);
  nor _72717_ (_21600_, _43000_, _21485_);
  or _72718_ (_21601_, _21600_, rst);
  or _72719_ (_43551_, _21601_, _21599_);
  not _72720_ (_21602_, \oc8051_golden_model_1.P2 [0]);
  nor _72721_ (_21603_, _43000_, _21602_);
  or _72722_ (_21605_, _21603_, rst);
  nor _72723_ (_21606_, _05235_, _21602_);
  and _72724_ (_21607_, _12128_, _05235_);
  or _72725_ (_21608_, _21607_, _21606_);
  and _72726_ (_21609_, _21608_, _03780_);
  and _72727_ (_21610_, _05235_, _04620_);
  or _72728_ (_21611_, _21610_, _21606_);
  or _72729_ (_21612_, _21611_, _06838_);
  nor _72730_ (_21613_, _05666_, _09454_);
  or _72731_ (_21614_, _21613_, _21606_);
  and _72732_ (_21616_, _21614_, _03610_);
  nor _72733_ (_21617_, _04409_, _21602_);
  and _72734_ (_21618_, _05235_, \oc8051_golden_model_1.ACC [0]);
  or _72735_ (_21619_, _21618_, _21606_);
  and _72736_ (_21620_, _21619_, _04409_);
  or _72737_ (_21621_, _21620_, _21617_);
  and _72738_ (_21622_, _21621_, _04081_);
  or _72739_ (_21623_, _21622_, _03715_);
  or _72740_ (_21624_, _21623_, _21616_);
  and _72741_ (_21625_, _12021_, _05918_);
  nor _72742_ (_21627_, _05918_, _21602_);
  or _72743_ (_21628_, _21627_, _04055_);
  or _72744_ (_21629_, _21628_, _21625_);
  and _72745_ (_21630_, _21629_, _03996_);
  and _72746_ (_21631_, _21630_, _21624_);
  and _72747_ (_21632_, _21611_, _03723_);
  or _72748_ (_21633_, _21632_, _03729_);
  or _72749_ (_21634_, _21633_, _21631_);
  or _72750_ (_21635_, _21619_, _03737_);
  and _72751_ (_21636_, _21635_, _03736_);
  and _72752_ (_21638_, _21636_, _21634_);
  and _72753_ (_21639_, _21606_, _03714_);
  or _72754_ (_21640_, _21639_, _03719_);
  or _72755_ (_21641_, _21640_, _21638_);
  or _72756_ (_21642_, _21614_, _06840_);
  and _72757_ (_21643_, _21642_, _03710_);
  and _72758_ (_21644_, _21643_, _21641_);
  and _72759_ (_21645_, _20023_, _05918_);
  or _72760_ (_21646_, _21645_, _21627_);
  and _72761_ (_21647_, _21646_, _03505_);
  or _72762_ (_21649_, _21647_, _07390_);
  or _72763_ (_21650_, _21649_, _21644_);
  and _72764_ (_21651_, _21650_, _21612_);
  or _72765_ (_21652_, _21651_, _04481_);
  and _72766_ (_21653_, _06546_, _05235_);
  or _72767_ (_21654_, _21606_, _07400_);
  or _72768_ (_21655_, _21654_, _21653_);
  and _72769_ (_21656_, _21655_, _03589_);
  and _72770_ (_21657_, _21656_, _21652_);
  and _72771_ (_21658_, _20049_, _05235_);
  or _72772_ (_21660_, _21658_, _21606_);
  and _72773_ (_21661_, _21660_, _03222_);
  or _72774_ (_21662_, _21661_, _21657_);
  or _72775_ (_21663_, _21662_, _08828_);
  and _72776_ (_21664_, _12124_, _05235_);
  or _72777_ (_21665_, _21606_, _07766_);
  or _72778_ (_21666_, _21665_, _21664_);
  and _72779_ (_21667_, _05235_, _06274_);
  or _72780_ (_21668_, _21667_, _21606_);
  or _72781_ (_21669_, _21668_, _05886_);
  and _72782_ (_21671_, _21669_, _07778_);
  and _72783_ (_21672_, _21671_, _21666_);
  and _72784_ (_21673_, _21672_, _21663_);
  or _72785_ (_21674_, _21673_, _21609_);
  and _72786_ (_21675_, _21674_, _07777_);
  nand _72787_ (_21676_, _21668_, _03622_);
  nor _72788_ (_21677_, _21676_, _21613_);
  or _72789_ (_21678_, _21677_, _21675_);
  and _72790_ (_21679_, _21678_, _06828_);
  or _72791_ (_21680_, _21606_, _05666_);
  and _72792_ (_21682_, _21619_, _03790_);
  and _72793_ (_21683_, _21682_, _21680_);
  or _72794_ (_21684_, _21683_, _03624_);
  or _72795_ (_21685_, _21684_, _21679_);
  nor _72796_ (_21686_, _12122_, _09454_);
  or _72797_ (_21687_, _21606_, _07795_);
  or _72798_ (_21688_, _21687_, _21686_);
  and _72799_ (_21689_, _21688_, _07793_);
  and _72800_ (_21690_, _21689_, _21685_);
  nor _72801_ (_21691_, _12003_, _09454_);
  or _72802_ (_21693_, _21691_, _21606_);
  and _72803_ (_21694_, _21693_, _03785_);
  or _72804_ (_21695_, _21694_, _03815_);
  or _72805_ (_21696_, _21695_, _21690_);
  or _72806_ (_21697_, _21614_, _04246_);
  and _72807_ (_21698_, _21697_, _03823_);
  and _72808_ (_21699_, _21698_, _21696_);
  and _72809_ (_21700_, _21606_, _03453_);
  or _72810_ (_21701_, _21700_, _03447_);
  or _72811_ (_21702_, _21701_, _21699_);
  or _72812_ (_21704_, _21614_, _03514_);
  and _72813_ (_21705_, _21704_, _43000_);
  and _72814_ (_21706_, _21705_, _21702_);
  or _72815_ (_43552_, _21706_, _21605_);
  or _72816_ (_21707_, _05235_, \oc8051_golden_model_1.P2 [1]);
  and _72817_ (_21708_, _12213_, _05235_);
  not _72818_ (_21709_, _21708_);
  and _72819_ (_21710_, _21709_, _21707_);
  or _72820_ (_21711_, _21710_, _04081_);
  nand _72821_ (_21712_, _05235_, _03274_);
  and _72822_ (_21714_, _21712_, _21707_);
  and _72823_ (_21715_, _21714_, _04409_);
  not _72824_ (_21716_, \oc8051_golden_model_1.P2 [1]);
  nor _72825_ (_21717_, _04409_, _21716_);
  or _72826_ (_21718_, _21717_, _03610_);
  or _72827_ (_21719_, _21718_, _21715_);
  and _72828_ (_21720_, _21719_, _04055_);
  and _72829_ (_21721_, _21720_, _21711_);
  and _72830_ (_21722_, _12224_, _05918_);
  nor _72831_ (_21723_, _05918_, _21716_);
  or _72832_ (_21725_, _21723_, _03723_);
  or _72833_ (_21726_, _21725_, _21722_);
  and _72834_ (_21727_, _21726_, _14265_);
  or _72835_ (_21728_, _21727_, _21721_);
  nor _72836_ (_21729_, _05235_, _21716_);
  and _72837_ (_21730_, _05235_, _06764_);
  or _72838_ (_21731_, _21730_, _21729_);
  or _72839_ (_21732_, _21731_, _03996_);
  and _72840_ (_21733_, _21732_, _21728_);
  or _72841_ (_21734_, _21733_, _03729_);
  or _72842_ (_21736_, _21714_, _03737_);
  and _72843_ (_21737_, _21736_, _03736_);
  and _72844_ (_21738_, _21737_, _21734_);
  and _72845_ (_21739_, _12211_, _05918_);
  or _72846_ (_21740_, _21739_, _21723_);
  and _72847_ (_21741_, _21740_, _03714_);
  or _72848_ (_21742_, _21741_, _03719_);
  or _72849_ (_21743_, _21742_, _21738_);
  and _72850_ (_21744_, _21722_, _12239_);
  or _72851_ (_21745_, _21723_, _06840_);
  or _72852_ (_21747_, _21745_, _21744_);
  and _72853_ (_21748_, _21747_, _21743_);
  and _72854_ (_21749_, _21748_, _03710_);
  and _72855_ (_21750_, _20141_, _05918_);
  or _72856_ (_21751_, _21723_, _21750_);
  and _72857_ (_21752_, _21751_, _03505_);
  or _72858_ (_21753_, _21752_, _07390_);
  or _72859_ (_21754_, _21753_, _21749_);
  or _72860_ (_21755_, _21731_, _06838_);
  and _72861_ (_21756_, _21755_, _21754_);
  or _72862_ (_21758_, _21756_, _04481_);
  and _72863_ (_21759_, _06501_, _05235_);
  or _72864_ (_21760_, _21729_, _07400_);
  or _72865_ (_21761_, _21760_, _21759_);
  and _72866_ (_21762_, _21761_, _03589_);
  and _72867_ (_21763_, _21762_, _21758_);
  and _72868_ (_21764_, _20168_, _05235_);
  or _72869_ (_21765_, _21764_, _21729_);
  and _72870_ (_21766_, _21765_, _03222_);
  or _72871_ (_21767_, _21766_, _21763_);
  and _72872_ (_21769_, _21767_, _03602_);
  or _72873_ (_21770_, _12327_, _09454_);
  and _72874_ (_21771_, _21770_, _03600_);
  nand _72875_ (_21772_, _05235_, _04303_);
  and _72876_ (_21773_, _21772_, _03601_);
  or _72877_ (_21774_, _21773_, _21771_);
  and _72878_ (_21775_, _21774_, _21707_);
  or _72879_ (_21776_, _21775_, _21769_);
  and _72880_ (_21777_, _21776_, _07778_);
  or _72881_ (_21778_, _12333_, _09454_);
  and _72882_ (_21780_, _21707_, _03780_);
  and _72883_ (_21781_, _21780_, _21778_);
  or _72884_ (_21782_, _21781_, _21777_);
  and _72885_ (_21783_, _21782_, _07777_);
  or _72886_ (_21784_, _12207_, _09454_);
  and _72887_ (_21785_, _21707_, _03622_);
  and _72888_ (_21786_, _21785_, _21784_);
  or _72889_ (_21787_, _21786_, _21783_);
  and _72890_ (_21788_, _21787_, _06828_);
  or _72891_ (_21789_, _21729_, _05618_);
  and _72892_ (_21791_, _21714_, _03790_);
  and _72893_ (_21792_, _21791_, _21789_);
  or _72894_ (_21793_, _21792_, _21788_);
  and _72895_ (_21794_, _21793_, _03786_);
  or _72896_ (_21795_, _21772_, _05618_);
  and _72897_ (_21796_, _21707_, _03624_);
  and _72898_ (_21797_, _21796_, _21795_);
  or _72899_ (_21798_, _21712_, _05618_);
  and _72900_ (_21799_, _21707_, _03785_);
  and _72901_ (_21800_, _21799_, _21798_);
  or _72902_ (_21802_, _21800_, _03815_);
  or _72903_ (_21803_, _21802_, _21797_);
  or _72904_ (_21804_, _21803_, _21794_);
  or _72905_ (_21805_, _21710_, _04246_);
  and _72906_ (_21806_, _21805_, _03823_);
  and _72907_ (_21807_, _21806_, _21804_);
  and _72908_ (_21808_, _21740_, _03453_);
  or _72909_ (_21809_, _21808_, _03447_);
  or _72910_ (_21810_, _21809_, _21807_);
  or _72911_ (_21811_, _21729_, _03514_);
  or _72912_ (_21813_, _21811_, _21708_);
  and _72913_ (_21814_, _21813_, _43000_);
  and _72914_ (_21815_, _21814_, _21810_);
  nor _72915_ (_21816_, _43000_, _21716_);
  or _72916_ (_21817_, _21816_, rst);
  or _72917_ (_43553_, _21817_, _21815_);
  not _72918_ (_21818_, \oc8051_golden_model_1.P2 [2]);
  nor _72919_ (_21819_, _43000_, _21818_);
  or _72920_ (_21820_, _21819_, rst);
  nor _72921_ (_21821_, _05235_, _21818_);
  nor _72922_ (_21823_, _09454_, _04875_);
  or _72923_ (_21824_, _21823_, _21821_);
  or _72924_ (_21825_, _21824_, _06838_);
  or _72925_ (_21826_, _21824_, _03996_);
  nor _72926_ (_21827_, _12416_, _09454_);
  or _72927_ (_21828_, _21827_, _21821_);
  or _72928_ (_21829_, _21828_, _04081_);
  and _72929_ (_21830_, _05235_, \oc8051_golden_model_1.ACC [2]);
  or _72930_ (_21831_, _21830_, _21821_);
  and _72931_ (_21832_, _21831_, _04409_);
  nor _72932_ (_21834_, _04409_, _21818_);
  or _72933_ (_21835_, _21834_, _03610_);
  or _72934_ (_21836_, _21835_, _21832_);
  and _72935_ (_21837_, _21836_, _04055_);
  and _72936_ (_21838_, _21837_, _21829_);
  nor _72937_ (_21839_, _05918_, _21818_);
  and _72938_ (_21840_, _12411_, _05918_);
  or _72939_ (_21841_, _21840_, _21839_);
  and _72940_ (_21842_, _21841_, _03715_);
  or _72941_ (_21843_, _21842_, _03723_);
  or _72942_ (_21845_, _21843_, _21838_);
  and _72943_ (_21846_, _21845_, _21826_);
  or _72944_ (_21847_, _21846_, _03729_);
  or _72945_ (_21848_, _21831_, _03737_);
  and _72946_ (_21849_, _21848_, _03736_);
  and _72947_ (_21850_, _21849_, _21847_);
  and _72948_ (_21851_, _12409_, _05918_);
  or _72949_ (_21852_, _21851_, _21839_);
  and _72950_ (_21853_, _21852_, _03714_);
  or _72951_ (_21854_, _21853_, _03719_);
  or _72952_ (_21856_, _21854_, _21850_);
  and _72953_ (_21857_, _21840_, _12443_);
  or _72954_ (_21858_, _21839_, _06840_);
  or _72955_ (_21859_, _21858_, _21857_);
  and _72956_ (_21860_, _21859_, _03710_);
  and _72957_ (_21861_, _21860_, _21856_);
  and _72958_ (_21862_, _20264_, _05918_);
  or _72959_ (_21863_, _21862_, _21839_);
  and _72960_ (_21864_, _21863_, _03505_);
  or _72961_ (_21865_, _21864_, _07390_);
  or _72962_ (_21867_, _21865_, _21861_);
  and _72963_ (_21868_, _21867_, _21825_);
  or _72964_ (_21869_, _21868_, _04481_);
  and _72965_ (_21870_, _06637_, _05235_);
  or _72966_ (_21871_, _21821_, _07400_);
  or _72967_ (_21872_, _21871_, _21870_);
  and _72968_ (_21873_, _21872_, _03589_);
  and _72969_ (_21874_, _21873_, _21869_);
  and _72970_ (_21875_, _20290_, _05235_);
  or _72971_ (_21876_, _21821_, _21875_);
  and _72972_ (_21878_, _21876_, _03222_);
  or _72973_ (_21879_, _21878_, _21874_);
  or _72974_ (_21880_, _21879_, _08828_);
  and _72975_ (_21881_, _12533_, _05235_);
  or _72976_ (_21882_, _21821_, _07766_);
  or _72977_ (_21883_, _21882_, _21881_);
  and _72978_ (_21884_, _05235_, _06332_);
  or _72979_ (_21885_, _21884_, _21821_);
  or _72980_ (_21886_, _21885_, _05886_);
  and _72981_ (_21887_, _21886_, _07778_);
  and _72982_ (_21889_, _21887_, _21883_);
  and _72983_ (_21890_, _21889_, _21880_);
  and _72984_ (_21891_, _12539_, _05235_);
  or _72985_ (_21892_, _21891_, _21821_);
  and _72986_ (_21893_, _21892_, _03780_);
  or _72987_ (_21894_, _21893_, _21890_);
  and _72988_ (_21895_, _21894_, _07777_);
  or _72989_ (_21896_, _21821_, _05718_);
  and _72990_ (_21897_, _21885_, _03622_);
  and _72991_ (_21898_, _21897_, _21896_);
  or _72992_ (_21900_, _21898_, _21895_);
  and _72993_ (_21901_, _21900_, _06828_);
  and _72994_ (_21902_, _21831_, _03790_);
  and _72995_ (_21903_, _21902_, _21896_);
  or _72996_ (_21904_, _21903_, _03624_);
  or _72997_ (_21905_, _21904_, _21901_);
  nor _72998_ (_21906_, _12532_, _09454_);
  or _72999_ (_21907_, _21821_, _07795_);
  or _73000_ (_21908_, _21907_, _21906_);
  and _73001_ (_21909_, _21908_, _07793_);
  and _73002_ (_21911_, _21909_, _21905_);
  nor _73003_ (_21912_, _12538_, _09454_);
  or _73004_ (_21913_, _21912_, _21821_);
  and _73005_ (_21914_, _21913_, _03785_);
  or _73006_ (_21915_, _21914_, _03815_);
  or _73007_ (_21916_, _21915_, _21911_);
  or _73008_ (_21917_, _21828_, _04246_);
  and _73009_ (_21918_, _21917_, _03823_);
  and _73010_ (_21919_, _21918_, _21916_);
  and _73011_ (_21920_, _21852_, _03453_);
  or _73012_ (_21922_, _21920_, _03447_);
  or _73013_ (_21923_, _21922_, _21919_);
  and _73014_ (_21924_, _12592_, _05235_);
  or _73015_ (_21925_, _21821_, _03514_);
  or _73016_ (_21926_, _21925_, _21924_);
  and _73017_ (_21927_, _21926_, _43000_);
  and _73018_ (_21928_, _21927_, _21923_);
  or _73019_ (_43554_, _21928_, _21820_);
  and _73020_ (_21929_, _09454_, \oc8051_golden_model_1.P2 [3]);
  nor _73021_ (_21930_, _09454_, _05005_);
  or _73022_ (_21932_, _21930_, _21929_);
  or _73023_ (_21933_, _21932_, _06838_);
  nor _73024_ (_21934_, _12627_, _09454_);
  or _73025_ (_21935_, _21934_, _21929_);
  or _73026_ (_21936_, _21935_, _04081_);
  and _73027_ (_21937_, _05235_, \oc8051_golden_model_1.ACC [3]);
  or _73028_ (_21938_, _21937_, _21929_);
  and _73029_ (_21939_, _21938_, _04409_);
  and _73030_ (_21940_, _09029_, \oc8051_golden_model_1.P2 [3]);
  or _73031_ (_21941_, _21940_, _03610_);
  or _73032_ (_21943_, _21941_, _21939_);
  and _73033_ (_21944_, _21943_, _04055_);
  and _73034_ (_21945_, _21944_, _21936_);
  not _73035_ (_21946_, _05918_);
  and _73036_ (_21947_, _21946_, \oc8051_golden_model_1.P2 [3]);
  and _73037_ (_21948_, _12631_, _05918_);
  or _73038_ (_21949_, _21948_, _21947_);
  and _73039_ (_21950_, _21949_, _03715_);
  or _73040_ (_21951_, _21950_, _03723_);
  or _73041_ (_21952_, _21951_, _21945_);
  or _73042_ (_21954_, _21932_, _03996_);
  and _73043_ (_21955_, _21954_, _21952_);
  or _73044_ (_21956_, _21955_, _03729_);
  or _73045_ (_21957_, _21938_, _03737_);
  and _73046_ (_21958_, _21957_, _03736_);
  and _73047_ (_21959_, _21958_, _21956_);
  and _73048_ (_21960_, _12641_, _05918_);
  or _73049_ (_21961_, _21960_, _21947_);
  and _73050_ (_21962_, _21961_, _03714_);
  or _73051_ (_21963_, _21962_, _03719_);
  or _73052_ (_21965_, _21963_, _21959_);
  or _73053_ (_21966_, _21947_, _12648_);
  and _73054_ (_21967_, _21966_, _21949_);
  or _73055_ (_21968_, _21967_, _06840_);
  and _73056_ (_21969_, _21968_, _03710_);
  and _73057_ (_21970_, _21969_, _21965_);
  and _73058_ (_21971_, _20391_, _05918_);
  or _73059_ (_21972_, _21971_, _21947_);
  and _73060_ (_21973_, _21972_, _03505_);
  or _73061_ (_21974_, _21973_, _07390_);
  or _73062_ (_21976_, _21974_, _21970_);
  and _73063_ (_21977_, _21976_, _21933_);
  or _73064_ (_21978_, _21977_, _04481_);
  and _73065_ (_21979_, _06592_, _05235_);
  or _73066_ (_21980_, _21929_, _07400_);
  or _73067_ (_21981_, _21980_, _21979_);
  and _73068_ (_21982_, _21981_, _03589_);
  and _73069_ (_21983_, _21982_, _21978_);
  and _73070_ (_21984_, _20416_, _05235_);
  or _73071_ (_21985_, _21929_, _21984_);
  and _73072_ (_21987_, _21985_, _03222_);
  or _73073_ (_21988_, _21987_, _21983_);
  or _73074_ (_21989_, _21988_, _08828_);
  and _73075_ (_21990_, _12733_, _05235_);
  or _73076_ (_21991_, _21929_, _07766_);
  or _73077_ (_21992_, _21991_, _21990_);
  and _73078_ (_21993_, _05235_, _06276_);
  or _73079_ (_21994_, _21993_, _21929_);
  or _73080_ (_21995_, _21994_, _05886_);
  and _73081_ (_21996_, _21995_, _07778_);
  and _73082_ (_21998_, _21996_, _21992_);
  and _73083_ (_21999_, _21998_, _21989_);
  and _73084_ (_22000_, _12739_, _05235_);
  or _73085_ (_22001_, _22000_, _21929_);
  and _73086_ (_22002_, _22001_, _03780_);
  or _73087_ (_22003_, _22002_, _21999_);
  and _73088_ (_22004_, _22003_, _07777_);
  or _73089_ (_22005_, _21929_, _05567_);
  and _73090_ (_22006_, _21994_, _03622_);
  and _73091_ (_22007_, _22006_, _22005_);
  or _73092_ (_22009_, _22007_, _22004_);
  and _73093_ (_22010_, _22009_, _06828_);
  and _73094_ (_22011_, _21938_, _03790_);
  and _73095_ (_22012_, _22011_, _22005_);
  or _73096_ (_22013_, _22012_, _03624_);
  or _73097_ (_22014_, _22013_, _22010_);
  nor _73098_ (_22015_, _12732_, _09454_);
  or _73099_ (_22016_, _21929_, _07795_);
  or _73100_ (_22017_, _22016_, _22015_);
  and _73101_ (_22018_, _22017_, _07793_);
  and _73102_ (_22020_, _22018_, _22014_);
  nor _73103_ (_22021_, _12738_, _09454_);
  or _73104_ (_22022_, _22021_, _21929_);
  and _73105_ (_22023_, _22022_, _03785_);
  or _73106_ (_22024_, _22023_, _03815_);
  or _73107_ (_22025_, _22024_, _22020_);
  or _73108_ (_22026_, _21935_, _04246_);
  and _73109_ (_22027_, _22026_, _03823_);
  and _73110_ (_22028_, _22027_, _22025_);
  and _73111_ (_22029_, _21961_, _03453_);
  or _73112_ (_22031_, _22029_, _03447_);
  or _73113_ (_22032_, _22031_, _22028_);
  and _73114_ (_22033_, _12794_, _05235_);
  or _73115_ (_22034_, _21929_, _03514_);
  or _73116_ (_22035_, _22034_, _22033_);
  and _73117_ (_22036_, _22035_, _43000_);
  and _73118_ (_22037_, _22036_, _22032_);
  nor _73119_ (_22038_, \oc8051_golden_model_1.P2 [3], rst);
  nor _73120_ (_22039_, _22038_, _04794_);
  or _73121_ (_43555_, _22039_, _22037_);
  nor _73122_ (_22041_, \oc8051_golden_model_1.P2 [4], rst);
  nor _73123_ (_22042_, _22041_, _04794_);
  and _73124_ (_22043_, _09454_, \oc8051_golden_model_1.P2 [4]);
  nor _73125_ (_22044_, _05777_, _09454_);
  or _73126_ (_22045_, _22044_, _22043_);
  or _73127_ (_22046_, _22045_, _06838_);
  and _73128_ (_22047_, _21946_, \oc8051_golden_model_1.P2 [4]);
  and _73129_ (_22048_, _12827_, _05918_);
  or _73130_ (_22049_, _22048_, _22047_);
  and _73131_ (_22050_, _22049_, _03714_);
  nor _73132_ (_22051_, _12841_, _09454_);
  or _73133_ (_22052_, _22051_, _22043_);
  or _73134_ (_22053_, _22052_, _04081_);
  and _73135_ (_22054_, _05235_, \oc8051_golden_model_1.ACC [4]);
  or _73136_ (_22055_, _22054_, _22043_);
  and _73137_ (_22056_, _22055_, _04409_);
  and _73138_ (_22057_, _09029_, \oc8051_golden_model_1.P2 [4]);
  or _73139_ (_22058_, _22057_, _03610_);
  or _73140_ (_22059_, _22058_, _22056_);
  and _73141_ (_22060_, _22059_, _04055_);
  and _73142_ (_22063_, _22060_, _22053_);
  and _73143_ (_22064_, _12845_, _05918_);
  or _73144_ (_22065_, _22064_, _22047_);
  and _73145_ (_22066_, _22065_, _03715_);
  or _73146_ (_22067_, _22066_, _03723_);
  or _73147_ (_22068_, _22067_, _22063_);
  or _73148_ (_22069_, _22045_, _03996_);
  and _73149_ (_22070_, _22069_, _22068_);
  or _73150_ (_22071_, _22070_, _03729_);
  or _73151_ (_22072_, _22055_, _03737_);
  and _73152_ (_22074_, _22072_, _03736_);
  and _73153_ (_22075_, _22074_, _22071_);
  or _73154_ (_22076_, _22075_, _22050_);
  and _73155_ (_22077_, _22076_, _06840_);
  and _73156_ (_22078_, _12861_, _05918_);
  or _73157_ (_22079_, _22078_, _22047_);
  and _73158_ (_22080_, _22079_, _03719_);
  or _73159_ (_22081_, _22080_, _22077_);
  and _73160_ (_22082_, _22081_, _03710_);
  and _73161_ (_22083_, _20511_, _05918_);
  or _73162_ (_22085_, _22083_, _22047_);
  and _73163_ (_22086_, _22085_, _03505_);
  or _73164_ (_22087_, _22086_, _07390_);
  or _73165_ (_22088_, _22087_, _22082_);
  and _73166_ (_22089_, _22088_, _22046_);
  or _73167_ (_22090_, _22089_, _04481_);
  and _73168_ (_22091_, _06730_, _05235_);
  or _73169_ (_22092_, _22043_, _07400_);
  or _73170_ (_22093_, _22092_, _22091_);
  and _73171_ (_22094_, _22093_, _03589_);
  and _73172_ (_22096_, _22094_, _22090_);
  and _73173_ (_22097_, _20536_, _05235_);
  or _73174_ (_22098_, _22097_, _22043_);
  and _73175_ (_22099_, _22098_, _03222_);
  or _73176_ (_22100_, _22099_, _08828_);
  or _73177_ (_22101_, _22100_, _22096_);
  and _73178_ (_22102_, _12821_, _05235_);
  or _73179_ (_22103_, _22043_, _07766_);
  or _73180_ (_22104_, _22103_, _22102_);
  and _73181_ (_22105_, _06298_, _05235_);
  or _73182_ (_22107_, _22105_, _22043_);
  or _73183_ (_22108_, _22107_, _05886_);
  and _73184_ (_22109_, _22108_, _07778_);
  and _73185_ (_22110_, _22109_, _22104_);
  and _73186_ (_22111_, _22110_, _22101_);
  and _73187_ (_22112_, _12817_, _05235_);
  or _73188_ (_22113_, _22112_, _22043_);
  and _73189_ (_22114_, _22113_, _03780_);
  or _73190_ (_22115_, _22114_, _22111_);
  and _73191_ (_22116_, _22115_, _07777_);
  or _73192_ (_22118_, _22043_, _05825_);
  and _73193_ (_22119_, _22107_, _03622_);
  and _73194_ (_22120_, _22119_, _22118_);
  or _73195_ (_22121_, _22120_, _22116_);
  and _73196_ (_22122_, _22121_, _06828_);
  and _73197_ (_22123_, _22055_, _03790_);
  and _73198_ (_22124_, _22123_, _22118_);
  or _73199_ (_22125_, _22124_, _03624_);
  or _73200_ (_22126_, _22125_, _22122_);
  nor _73201_ (_22127_, _12819_, _09454_);
  or _73202_ (_22129_, _22043_, _07795_);
  or _73203_ (_22130_, _22129_, _22127_);
  and _73204_ (_22131_, _22130_, _07793_);
  and _73205_ (_22132_, _22131_, _22126_);
  nor _73206_ (_22133_, _12816_, _09454_);
  or _73207_ (_22134_, _22133_, _22043_);
  and _73208_ (_22135_, _22134_, _03785_);
  or _73209_ (_22136_, _22135_, _03815_);
  or _73210_ (_22137_, _22136_, _22132_);
  or _73211_ (_22138_, _22052_, _04246_);
  and _73212_ (_22140_, _22138_, _03823_);
  and _73213_ (_22141_, _22140_, _22137_);
  and _73214_ (_22142_, _22049_, _03453_);
  or _73215_ (_22143_, _22142_, _03447_);
  or _73216_ (_22144_, _22143_, _22141_);
  and _73217_ (_22145_, _13003_, _05235_);
  or _73218_ (_22146_, _22043_, _03514_);
  or _73219_ (_22147_, _22146_, _22145_);
  and _73220_ (_22148_, _22147_, _43000_);
  and _73221_ (_22149_, _22148_, _22144_);
  or _73222_ (_43556_, _22149_, _22042_);
  and _73223_ (_22151_, _09454_, \oc8051_golden_model_1.P2 [5]);
  nor _73224_ (_22152_, _13014_, _09454_);
  or _73225_ (_22153_, _22152_, _22151_);
  or _73226_ (_22154_, _22153_, _04081_);
  and _73227_ (_22155_, _05235_, \oc8051_golden_model_1.ACC [5]);
  or _73228_ (_22156_, _22155_, _22151_);
  and _73229_ (_22157_, _22156_, _04409_);
  and _73230_ (_22158_, _09029_, \oc8051_golden_model_1.P2 [5]);
  or _73231_ (_22159_, _22158_, _03610_);
  or _73232_ (_22161_, _22159_, _22157_);
  and _73233_ (_22162_, _22161_, _04055_);
  and _73234_ (_22163_, _22162_, _22154_);
  and _73235_ (_22164_, _21946_, \oc8051_golden_model_1.P2 [5]);
  and _73236_ (_22165_, _13037_, _05918_);
  or _73237_ (_22166_, _22165_, _22164_);
  and _73238_ (_22167_, _22166_, _03715_);
  or _73239_ (_22168_, _22167_, _03723_);
  or _73240_ (_22169_, _22168_, _22163_);
  nor _73241_ (_22170_, _05469_, _09454_);
  or _73242_ (_22172_, _22170_, _22151_);
  or _73243_ (_22173_, _22172_, _03996_);
  and _73244_ (_22174_, _22173_, _22169_);
  or _73245_ (_22175_, _22174_, _03729_);
  or _73246_ (_22176_, _22156_, _03737_);
  and _73247_ (_22177_, _22176_, _03736_);
  and _73248_ (_22178_, _22177_, _22175_);
  and _73249_ (_22179_, _13047_, _05918_);
  or _73250_ (_22180_, _22179_, _22164_);
  and _73251_ (_22181_, _22180_, _03714_);
  or _73252_ (_22183_, _22181_, _03719_);
  or _73253_ (_22184_, _22183_, _22178_);
  or _73254_ (_22185_, _22164_, _13054_);
  and _73255_ (_22186_, _22185_, _22166_);
  or _73256_ (_22187_, _22186_, _06840_);
  and _73257_ (_22188_, _22187_, _03710_);
  and _73258_ (_22189_, _22188_, _22184_);
  and _73259_ (_22190_, _20633_, _05918_);
  or _73260_ (_22191_, _22190_, _22164_);
  and _73261_ (_22192_, _22191_, _03505_);
  or _73262_ (_22194_, _22192_, _07390_);
  or _73263_ (_22195_, _22194_, _22189_);
  or _73264_ (_22196_, _22172_, _06838_);
  and _73265_ (_22197_, _22196_, _22195_);
  or _73266_ (_22198_, _22197_, _04481_);
  and _73267_ (_22199_, _06684_, _05235_);
  or _73268_ (_22200_, _22151_, _07400_);
  or _73269_ (_22201_, _22200_, _22199_);
  and _73270_ (_22202_, _22201_, _03589_);
  and _73271_ (_22203_, _22202_, _22198_);
  and _73272_ (_22205_, _20660_, _05235_);
  or _73273_ (_22206_, _22205_, _22151_);
  and _73274_ (_22207_, _22206_, _03222_);
  or _73275_ (_22208_, _22207_, _08828_);
  or _73276_ (_22209_, _22208_, _22203_);
  and _73277_ (_22210_, _13141_, _05235_);
  or _73278_ (_22211_, _22151_, _07766_);
  or _73279_ (_22212_, _22211_, _22210_);
  and _73280_ (_22213_, _06306_, _05235_);
  or _73281_ (_22214_, _22213_, _22151_);
  or _73282_ (_22216_, _22214_, _05886_);
  and _73283_ (_22217_, _22216_, _07778_);
  and _73284_ (_22218_, _22217_, _22212_);
  and _73285_ (_22219_, _22218_, _22209_);
  and _73286_ (_22220_, _13147_, _05235_);
  or _73287_ (_22221_, _22220_, _22151_);
  and _73288_ (_22222_, _22221_, _03780_);
  or _73289_ (_22223_, _22222_, _22219_);
  and _73290_ (_22224_, _22223_, _07777_);
  or _73291_ (_22225_, _22151_, _05518_);
  and _73292_ (_22227_, _22214_, _03622_);
  and _73293_ (_22228_, _22227_, _22225_);
  or _73294_ (_22229_, _22228_, _22224_);
  and _73295_ (_22230_, _22229_, _06828_);
  and _73296_ (_22231_, _22156_, _03790_);
  and _73297_ (_22232_, _22231_, _22225_);
  or _73298_ (_22233_, _22232_, _03624_);
  or _73299_ (_22234_, _22233_, _22230_);
  nor _73300_ (_22235_, _13140_, _09454_);
  or _73301_ (_22236_, _22151_, _07795_);
  or _73302_ (_22238_, _22236_, _22235_);
  and _73303_ (_22239_, _22238_, _07793_);
  and _73304_ (_22240_, _22239_, _22234_);
  nor _73305_ (_22241_, _13146_, _09454_);
  or _73306_ (_22242_, _22241_, _22151_);
  and _73307_ (_22243_, _22242_, _03785_);
  or _73308_ (_22244_, _22243_, _03815_);
  or _73309_ (_22245_, _22244_, _22240_);
  or _73310_ (_22246_, _22153_, _04246_);
  and _73311_ (_22247_, _22246_, _03823_);
  and _73312_ (_22249_, _22247_, _22245_);
  and _73313_ (_22250_, _22180_, _03453_);
  or _73314_ (_22251_, _22250_, _03447_);
  or _73315_ (_22252_, _22251_, _22249_);
  and _73316_ (_22253_, _13199_, _05235_);
  or _73317_ (_22254_, _22151_, _03514_);
  or _73318_ (_22255_, _22254_, _22253_);
  and _73319_ (_22256_, _22255_, _43000_);
  and _73320_ (_22257_, _22256_, _22252_);
  nor _73321_ (_22258_, \oc8051_golden_model_1.P2 [5], rst);
  nor _73322_ (_22260_, _22258_, _04794_);
  or _73323_ (_43557_, _22260_, _22257_);
  not _73324_ (_22261_, \oc8051_golden_model_1.P2 [6]);
  nor _73325_ (_22262_, _43000_, _22261_);
  or _73326_ (_22263_, _22262_, rst);
  nor _73327_ (_22264_, _05235_, _22261_);
  nor _73328_ (_22265_, _13242_, _09454_);
  or _73329_ (_22266_, _22265_, _22264_);
  or _73330_ (_22267_, _22266_, _04081_);
  and _73331_ (_22268_, _05235_, \oc8051_golden_model_1.ACC [6]);
  or _73332_ (_22270_, _22268_, _22264_);
  and _73333_ (_22271_, _22270_, _04409_);
  nor _73334_ (_22272_, _04409_, _22261_);
  or _73335_ (_22273_, _22272_, _03610_);
  or _73336_ (_22274_, _22273_, _22271_);
  and _73337_ (_22275_, _22274_, _04055_);
  and _73338_ (_22276_, _22275_, _22267_);
  nor _73339_ (_22277_, _05918_, _22261_);
  and _73340_ (_22278_, _13229_, _05918_);
  or _73341_ (_22279_, _22278_, _22277_);
  and _73342_ (_22281_, _22279_, _03715_);
  or _73343_ (_22282_, _22281_, _03723_);
  or _73344_ (_22283_, _22282_, _22276_);
  nor _73345_ (_22284_, _05363_, _09454_);
  or _73346_ (_22285_, _22284_, _22264_);
  or _73347_ (_22286_, _22285_, _03996_);
  and _73348_ (_22287_, _22286_, _22283_);
  or _73349_ (_22288_, _22287_, _03729_);
  or _73350_ (_22289_, _22270_, _03737_);
  and _73351_ (_22290_, _22289_, _03736_);
  and _73352_ (_22292_, _22290_, _22288_);
  and _73353_ (_22293_, _13253_, _05918_);
  or _73354_ (_22294_, _22293_, _22277_);
  and _73355_ (_22295_, _22294_, _03714_);
  or _73356_ (_22296_, _22295_, _03719_);
  or _73357_ (_22297_, _22296_, _22292_);
  or _73358_ (_22298_, _22277_, _13260_);
  and _73359_ (_22299_, _22298_, _22279_);
  or _73360_ (_22300_, _22299_, _06840_);
  and _73361_ (_22301_, _22300_, _03710_);
  and _73362_ (_22303_, _22301_, _22297_);
  and _73363_ (_22304_, _20753_, _05918_);
  or _73364_ (_22305_, _22304_, _22277_);
  and _73365_ (_22306_, _22305_, _03505_);
  or _73366_ (_22307_, _22306_, _07390_);
  or _73367_ (_22308_, _22307_, _22303_);
  or _73368_ (_22309_, _22285_, _06838_);
  and _73369_ (_22310_, _22309_, _22308_);
  or _73370_ (_22311_, _22310_, _04481_);
  and _73371_ (_22312_, _06455_, _05235_);
  or _73372_ (_22314_, _22264_, _07400_);
  or _73373_ (_22315_, _22314_, _22312_);
  and _73374_ (_22316_, _22315_, _03589_);
  and _73375_ (_22317_, _22316_, _22311_);
  and _73376_ (_22318_, _20778_, _05235_);
  or _73377_ (_22319_, _22318_, _22264_);
  and _73378_ (_22320_, _22319_, _03222_);
  or _73379_ (_22321_, _22320_, _08828_);
  or _73380_ (_22322_, _22321_, _22317_);
  and _73381_ (_22323_, _13347_, _05235_);
  or _73382_ (_22326_, _22264_, _07766_);
  or _73383_ (_22327_, _22326_, _22323_);
  and _73384_ (_22328_, _13339_, _05235_);
  or _73385_ (_22329_, _22328_, _22264_);
  or _73386_ (_22330_, _22329_, _05886_);
  and _73387_ (_22331_, _22330_, _07778_);
  and _73388_ (_22332_, _22331_, _22327_);
  and _73389_ (_22333_, _22332_, _22322_);
  and _73390_ (_22334_, _13353_, _05235_);
  or _73391_ (_22335_, _22334_, _22264_);
  and _73392_ (_22337_, _22335_, _03780_);
  or _73393_ (_22338_, _22337_, _22333_);
  and _73394_ (_22339_, _22338_, _07777_);
  or _73395_ (_22340_, _22264_, _05412_);
  and _73396_ (_22341_, _22329_, _03622_);
  and _73397_ (_22342_, _22341_, _22340_);
  or _73398_ (_22343_, _22342_, _22339_);
  and _73399_ (_22344_, _22343_, _06828_);
  and _73400_ (_22345_, _22270_, _03790_);
  and _73401_ (_22346_, _22345_, _22340_);
  or _73402_ (_22348_, _22346_, _03624_);
  or _73403_ (_22349_, _22348_, _22344_);
  nor _73404_ (_22350_, _13346_, _09454_);
  or _73405_ (_22351_, _22264_, _07795_);
  or _73406_ (_22352_, _22351_, _22350_);
  and _73407_ (_22353_, _22352_, _07793_);
  and _73408_ (_22354_, _22353_, _22349_);
  nor _73409_ (_22355_, _13352_, _09454_);
  or _73410_ (_22356_, _22355_, _22264_);
  and _73411_ (_22357_, _22356_, _03785_);
  or _73412_ (_22359_, _22357_, _03815_);
  or _73413_ (_22360_, _22359_, _22354_);
  or _73414_ (_22361_, _22266_, _04246_);
  and _73415_ (_22362_, _22361_, _03823_);
  and _73416_ (_22363_, _22362_, _22360_);
  and _73417_ (_22364_, _22294_, _03453_);
  or _73418_ (_22365_, _22364_, _03447_);
  or _73419_ (_22366_, _22365_, _22363_);
  and _73420_ (_22367_, _13402_, _05235_);
  or _73421_ (_22368_, _22264_, _03514_);
  or _73422_ (_22370_, _22368_, _22367_);
  and _73423_ (_22371_, _22370_, _43000_);
  and _73424_ (_22372_, _22371_, _22366_);
  or _73425_ (_43558_, _22372_, _22263_);
  not _73426_ (_22373_, \oc8051_golden_model_1.P3 [0]);
  nor _73427_ (_22374_, _05239_, _22373_);
  and _73428_ (_22375_, _12128_, _05239_);
  or _73429_ (_22376_, _22375_, _22374_);
  and _73430_ (_22377_, _22376_, _03780_);
  and _73431_ (_22378_, _05239_, _04620_);
  or _73432_ (_22380_, _22378_, _22374_);
  or _73433_ (_22381_, _22380_, _06838_);
  nor _73434_ (_22382_, _05666_, _09557_);
  or _73435_ (_22383_, _22382_, _22374_);
  or _73436_ (_22384_, _22383_, _04081_);
  and _73437_ (_22385_, _05239_, \oc8051_golden_model_1.ACC [0]);
  or _73438_ (_22386_, _22385_, _22374_);
  and _73439_ (_22387_, _22386_, _04409_);
  nor _73440_ (_22388_, _04409_, _22373_);
  or _73441_ (_22389_, _22388_, _03610_);
  or _73442_ (_22391_, _22389_, _22387_);
  and _73443_ (_22392_, _22391_, _04055_);
  and _73444_ (_22393_, _22392_, _22384_);
  nor _73445_ (_22394_, _05929_, _22373_);
  and _73446_ (_22395_, _12021_, _05929_);
  or _73447_ (_22396_, _22395_, _22394_);
  and _73448_ (_22397_, _22396_, _03715_);
  or _73449_ (_22398_, _22397_, _22393_);
  and _73450_ (_22399_, _22398_, _03996_);
  and _73451_ (_22400_, _22380_, _03723_);
  or _73452_ (_22402_, _22400_, _03729_);
  or _73453_ (_22403_, _22402_, _22399_);
  or _73454_ (_22404_, _22386_, _03737_);
  and _73455_ (_22405_, _22404_, _03736_);
  and _73456_ (_22406_, _22405_, _22403_);
  and _73457_ (_22407_, _22374_, _03714_);
  or _73458_ (_22408_, _22407_, _03719_);
  or _73459_ (_22409_, _22408_, _22406_);
  or _73460_ (_22410_, _22383_, _06840_);
  and _73461_ (_22411_, _22410_, _03710_);
  and _73462_ (_22413_, _22411_, _22409_);
  and _73463_ (_22414_, _20023_, _05929_);
  or _73464_ (_22415_, _22414_, _22394_);
  and _73465_ (_22416_, _22415_, _03505_);
  or _73466_ (_22417_, _22416_, _07390_);
  or _73467_ (_22418_, _22417_, _22413_);
  and _73468_ (_22419_, _22418_, _22381_);
  or _73469_ (_22420_, _22419_, _04481_);
  and _73470_ (_22421_, _06546_, _05239_);
  or _73471_ (_22422_, _22374_, _07400_);
  or _73472_ (_22424_, _22422_, _22421_);
  and _73473_ (_22425_, _22424_, _03589_);
  and _73474_ (_22426_, _22425_, _22420_);
  and _73475_ (_22427_, _20049_, _05239_);
  or _73476_ (_22428_, _22427_, _22374_);
  and _73477_ (_22429_, _22428_, _03222_);
  or _73478_ (_22430_, _22429_, _22426_);
  or _73479_ (_22431_, _22430_, _08828_);
  and _73480_ (_22432_, _12124_, _05239_);
  or _73481_ (_22433_, _22374_, _07766_);
  or _73482_ (_22436_, _22433_, _22432_);
  and _73483_ (_22437_, _05239_, _06274_);
  or _73484_ (_22438_, _22437_, _22374_);
  or _73485_ (_22439_, _22438_, _05886_);
  and _73486_ (_22440_, _22439_, _07778_);
  and _73487_ (_22441_, _22440_, _22436_);
  and _73488_ (_22442_, _22441_, _22431_);
  or _73489_ (_22443_, _22442_, _22377_);
  and _73490_ (_22444_, _22443_, _07777_);
  nand _73491_ (_22445_, _22438_, _03622_);
  nor _73492_ (_22447_, _22445_, _22382_);
  or _73493_ (_22448_, _22447_, _22444_);
  and _73494_ (_22449_, _22448_, _06828_);
  or _73495_ (_22450_, _22374_, _05666_);
  and _73496_ (_22451_, _22386_, _03790_);
  and _73497_ (_22452_, _22451_, _22450_);
  or _73498_ (_22453_, _22452_, _03624_);
  or _73499_ (_22454_, _22453_, _22449_);
  nor _73500_ (_22455_, _12122_, _09557_);
  or _73501_ (_22456_, _22374_, _07795_);
  or _73502_ (_22458_, _22456_, _22455_);
  and _73503_ (_22459_, _22458_, _07793_);
  and _73504_ (_22460_, _22459_, _22454_);
  nor _73505_ (_22461_, _12003_, _09557_);
  or _73506_ (_22462_, _22461_, _22374_);
  and _73507_ (_22463_, _22462_, _03785_);
  or _73508_ (_22464_, _22463_, _03815_);
  or _73509_ (_22465_, _22464_, _22460_);
  or _73510_ (_22466_, _22383_, _04246_);
  and _73511_ (_22467_, _22466_, _03823_);
  and _73512_ (_22469_, _22467_, _22465_);
  and _73513_ (_22470_, _22374_, _03453_);
  or _73514_ (_22471_, _22470_, _03447_);
  or _73515_ (_22472_, _22471_, _22469_);
  or _73516_ (_22473_, _22383_, _03514_);
  and _73517_ (_22474_, _22473_, _43000_);
  and _73518_ (_22475_, _22474_, _22472_);
  nor _73519_ (_22476_, _43000_, _22373_);
  or _73520_ (_22477_, _22476_, rst);
  or _73521_ (_43561_, _22477_, _22475_);
  or _73522_ (_22479_, _05239_, \oc8051_golden_model_1.P3 [1]);
  and _73523_ (_22480_, _12213_, _05239_);
  not _73524_ (_22481_, _22480_);
  and _73525_ (_22482_, _22481_, _22479_);
  or _73526_ (_22483_, _22482_, _04081_);
  nand _73527_ (_22484_, _05239_, _03274_);
  and _73528_ (_22485_, _22484_, _22479_);
  and _73529_ (_22486_, _22485_, _04409_);
  not _73530_ (_22487_, \oc8051_golden_model_1.P3 [1]);
  nor _73531_ (_22488_, _04409_, _22487_);
  or _73532_ (_22490_, _22488_, _03610_);
  or _73533_ (_22491_, _22490_, _22486_);
  and _73534_ (_22492_, _22491_, _04055_);
  and _73535_ (_22493_, _22492_, _22483_);
  and _73536_ (_22494_, _12224_, _05929_);
  nor _73537_ (_22495_, _05929_, _22487_);
  or _73538_ (_22496_, _22495_, _03723_);
  or _73539_ (_22497_, _22496_, _22494_);
  and _73540_ (_22498_, _22497_, _14265_);
  or _73541_ (_22499_, _22498_, _22493_);
  nor _73542_ (_22501_, _05239_, _22487_);
  and _73543_ (_22502_, _05239_, _06764_);
  or _73544_ (_22503_, _22502_, _22501_);
  or _73545_ (_22504_, _22503_, _03996_);
  and _73546_ (_22505_, _22504_, _22499_);
  or _73547_ (_22506_, _22505_, _03729_);
  or _73548_ (_22507_, _22485_, _03737_);
  and _73549_ (_22508_, _22507_, _03736_);
  and _73550_ (_22509_, _22508_, _22506_);
  and _73551_ (_22510_, _12211_, _05929_);
  or _73552_ (_22512_, _22510_, _22495_);
  and _73553_ (_22513_, _22512_, _03714_);
  or _73554_ (_22514_, _22513_, _03719_);
  or _73555_ (_22515_, _22514_, _22509_);
  and _73556_ (_22516_, _22494_, _12239_);
  or _73557_ (_22517_, _22495_, _06840_);
  or _73558_ (_22518_, _22517_, _22516_);
  and _73559_ (_22519_, _22518_, _22515_);
  and _73560_ (_22520_, _22519_, _03710_);
  and _73561_ (_22521_, _20141_, _05929_);
  or _73562_ (_22523_, _22495_, _22521_);
  and _73563_ (_22524_, _22523_, _03505_);
  or _73564_ (_22525_, _22524_, _07390_);
  or _73565_ (_22526_, _22525_, _22520_);
  or _73566_ (_22527_, _22503_, _06838_);
  and _73567_ (_22528_, _22527_, _22526_);
  or _73568_ (_22529_, _22528_, _04481_);
  and _73569_ (_22530_, _06501_, _05239_);
  or _73570_ (_22531_, _22501_, _07400_);
  or _73571_ (_22532_, _22531_, _22530_);
  and _73572_ (_22534_, _22532_, _03589_);
  and _73573_ (_22535_, _22534_, _22529_);
  and _73574_ (_22536_, _20168_, _05239_);
  or _73575_ (_22537_, _22536_, _22501_);
  and _73576_ (_22538_, _22537_, _03222_);
  or _73577_ (_22539_, _22538_, _22535_);
  and _73578_ (_22540_, _22539_, _03602_);
  or _73579_ (_22541_, _12327_, _09557_);
  and _73580_ (_22542_, _22541_, _03600_);
  nand _73581_ (_22543_, _05239_, _04303_);
  and _73582_ (_22545_, _22543_, _03601_);
  or _73583_ (_22546_, _22545_, _22542_);
  and _73584_ (_22547_, _22546_, _22479_);
  or _73585_ (_22548_, _22547_, _22540_);
  and _73586_ (_22549_, _22548_, _07778_);
  or _73587_ (_22550_, _12333_, _09557_);
  and _73588_ (_22551_, _22479_, _03780_);
  and _73589_ (_22552_, _22551_, _22550_);
  or _73590_ (_22553_, _22552_, _22549_);
  and _73591_ (_22554_, _22553_, _07777_);
  or _73592_ (_22556_, _12207_, _09557_);
  and _73593_ (_22557_, _22479_, _03622_);
  and _73594_ (_22558_, _22557_, _22556_);
  or _73595_ (_22559_, _22558_, _22554_);
  and _73596_ (_22560_, _22559_, _06828_);
  or _73597_ (_22561_, _22501_, _05618_);
  and _73598_ (_22562_, _22485_, _03790_);
  and _73599_ (_22563_, _22562_, _22561_);
  or _73600_ (_22564_, _22563_, _22560_);
  and _73601_ (_22565_, _22564_, _03786_);
  or _73602_ (_22567_, _22543_, _05618_);
  and _73603_ (_22568_, _22479_, _03624_);
  and _73604_ (_22569_, _22568_, _22567_);
  or _73605_ (_22570_, _22484_, _05618_);
  and _73606_ (_22571_, _22479_, _03785_);
  and _73607_ (_22572_, _22571_, _22570_);
  or _73608_ (_22573_, _22572_, _03815_);
  or _73609_ (_22574_, _22573_, _22569_);
  or _73610_ (_22575_, _22574_, _22565_);
  or _73611_ (_22576_, _22482_, _04246_);
  and _73612_ (_22578_, _22576_, _03823_);
  and _73613_ (_22579_, _22578_, _22575_);
  and _73614_ (_22580_, _22512_, _03453_);
  or _73615_ (_22581_, _22580_, _03447_);
  or _73616_ (_22582_, _22581_, _22579_);
  or _73617_ (_22583_, _22501_, _03514_);
  or _73618_ (_22584_, _22583_, _22480_);
  and _73619_ (_22585_, _22584_, _43000_);
  and _73620_ (_22586_, _22585_, _22582_);
  nor _73621_ (_22587_, _43000_, _22487_);
  or _73622_ (_22589_, _22587_, rst);
  or _73623_ (_43562_, _22589_, _22586_);
  not _73624_ (_22590_, \oc8051_golden_model_1.P3 [2]);
  nor _73625_ (_22591_, _05239_, _22590_);
  nor _73626_ (_22592_, _09557_, _04875_);
  or _73627_ (_22593_, _22592_, _22591_);
  or _73628_ (_22594_, _22593_, _06838_);
  and _73629_ (_22595_, _22593_, _03723_);
  nor _73630_ (_22596_, _05929_, _22590_);
  and _73631_ (_22597_, _12411_, _05929_);
  or _73632_ (_22599_, _22597_, _22596_);
  or _73633_ (_22600_, _22599_, _04055_);
  nor _73634_ (_22601_, _12416_, _09557_);
  or _73635_ (_22602_, _22601_, _22591_);
  and _73636_ (_22603_, _22602_, _03610_);
  nor _73637_ (_22604_, _04409_, _22590_);
  and _73638_ (_22605_, _05239_, \oc8051_golden_model_1.ACC [2]);
  or _73639_ (_22606_, _22605_, _22591_);
  and _73640_ (_22607_, _22606_, _04409_);
  or _73641_ (_22608_, _22607_, _22604_);
  and _73642_ (_22610_, _22608_, _04081_);
  or _73643_ (_22611_, _22610_, _03715_);
  or _73644_ (_22612_, _22611_, _22603_);
  and _73645_ (_22613_, _22612_, _22600_);
  and _73646_ (_22614_, _22613_, _03996_);
  or _73647_ (_22615_, _22614_, _22595_);
  or _73648_ (_22616_, _22615_, _03729_);
  or _73649_ (_22617_, _22606_, _03737_);
  and _73650_ (_22618_, _22617_, _03736_);
  and _73651_ (_22619_, _22618_, _22616_);
  and _73652_ (_22621_, _12409_, _05929_);
  or _73653_ (_22622_, _22621_, _22596_);
  and _73654_ (_22623_, _22622_, _03714_);
  or _73655_ (_22624_, _22623_, _03719_);
  or _73656_ (_22625_, _22624_, _22619_);
  or _73657_ (_22626_, _22596_, _12443_);
  and _73658_ (_22627_, _22626_, _22599_);
  or _73659_ (_22628_, _22627_, _06840_);
  and _73660_ (_22629_, _22628_, _03710_);
  and _73661_ (_22630_, _22629_, _22625_);
  and _73662_ (_22632_, _20264_, _05929_);
  or _73663_ (_22633_, _22632_, _22596_);
  and _73664_ (_22634_, _22633_, _03505_);
  or _73665_ (_22635_, _22634_, _07390_);
  or _73666_ (_22636_, _22635_, _22630_);
  and _73667_ (_22637_, _22636_, _22594_);
  or _73668_ (_22638_, _22637_, _04481_);
  and _73669_ (_22639_, _06637_, _05239_);
  or _73670_ (_22640_, _22591_, _07400_);
  or _73671_ (_22641_, _22640_, _22639_);
  and _73672_ (_22643_, _22641_, _03589_);
  and _73673_ (_22644_, _22643_, _22638_);
  and _73674_ (_22645_, _20290_, _05239_);
  or _73675_ (_22646_, _22591_, _22645_);
  and _73676_ (_22647_, _22646_, _03222_);
  or _73677_ (_22648_, _22647_, _22644_);
  or _73678_ (_22649_, _22648_, _08828_);
  and _73679_ (_22650_, _12533_, _05239_);
  or _73680_ (_22651_, _22591_, _07766_);
  or _73681_ (_22652_, _22651_, _22650_);
  and _73682_ (_22654_, _05239_, _06332_);
  or _73683_ (_22655_, _22654_, _22591_);
  or _73684_ (_22656_, _22655_, _05886_);
  and _73685_ (_22657_, _22656_, _07778_);
  and _73686_ (_22658_, _22657_, _22652_);
  and _73687_ (_22659_, _22658_, _22649_);
  and _73688_ (_22660_, _12539_, _05239_);
  or _73689_ (_22661_, _22660_, _22591_);
  and _73690_ (_22662_, _22661_, _03780_);
  or _73691_ (_22663_, _22662_, _22659_);
  and _73692_ (_22665_, _22663_, _07777_);
  or _73693_ (_22666_, _22591_, _05718_);
  and _73694_ (_22667_, _22655_, _03622_);
  and _73695_ (_22668_, _22667_, _22666_);
  or _73696_ (_22669_, _22668_, _22665_);
  and _73697_ (_22670_, _22669_, _06828_);
  and _73698_ (_22671_, _22606_, _03790_);
  and _73699_ (_22672_, _22671_, _22666_);
  or _73700_ (_22673_, _22672_, _03624_);
  or _73701_ (_22674_, _22673_, _22670_);
  nor _73702_ (_22676_, _12532_, _09557_);
  or _73703_ (_22677_, _22591_, _07795_);
  or _73704_ (_22678_, _22677_, _22676_);
  and _73705_ (_22679_, _22678_, _07793_);
  and _73706_ (_22680_, _22679_, _22674_);
  nor _73707_ (_22681_, _12538_, _09557_);
  or _73708_ (_22682_, _22681_, _22591_);
  and _73709_ (_22683_, _22682_, _03785_);
  or _73710_ (_22684_, _22683_, _03815_);
  or _73711_ (_22685_, _22684_, _22680_);
  or _73712_ (_22687_, _22602_, _04246_);
  and _73713_ (_22688_, _22687_, _03823_);
  and _73714_ (_22689_, _22688_, _22685_);
  and _73715_ (_22690_, _22622_, _03453_);
  or _73716_ (_22691_, _22690_, _03447_);
  or _73717_ (_22692_, _22691_, _22689_);
  and _73718_ (_22693_, _12592_, _05239_);
  or _73719_ (_22694_, _22591_, _03514_);
  or _73720_ (_22695_, _22694_, _22693_);
  and _73721_ (_22696_, _22695_, _43000_);
  and _73722_ (_22698_, _22696_, _22692_);
  nor _73723_ (_22699_, _43000_, _22590_);
  or _73724_ (_22700_, _22699_, rst);
  or _73725_ (_43563_, _22700_, _22698_);
  and _73726_ (_22701_, _09557_, \oc8051_golden_model_1.P3 [3]);
  nor _73727_ (_22702_, _09557_, _05005_);
  or _73728_ (_22703_, _22702_, _22701_);
  or _73729_ (_22704_, _22703_, _06838_);
  nor _73730_ (_22705_, _12627_, _09557_);
  or _73731_ (_22706_, _22705_, _22701_);
  or _73732_ (_22708_, _22706_, _04081_);
  and _73733_ (_22709_, _05239_, \oc8051_golden_model_1.ACC [3]);
  or _73734_ (_22710_, _22709_, _22701_);
  and _73735_ (_22711_, _22710_, _04409_);
  and _73736_ (_22712_, _09029_, \oc8051_golden_model_1.P3 [3]);
  or _73737_ (_22713_, _22712_, _03610_);
  or _73738_ (_22714_, _22713_, _22711_);
  and _73739_ (_22715_, _22714_, _04055_);
  and _73740_ (_22716_, _22715_, _22708_);
  not _73741_ (_22717_, _05929_);
  and _73742_ (_22719_, _22717_, \oc8051_golden_model_1.P3 [3]);
  and _73743_ (_22720_, _12631_, _05929_);
  or _73744_ (_22721_, _22720_, _22719_);
  and _73745_ (_22722_, _22721_, _03715_);
  or _73746_ (_22723_, _22722_, _03723_);
  or _73747_ (_22724_, _22723_, _22716_);
  or _73748_ (_22725_, _22703_, _03996_);
  and _73749_ (_22726_, _22725_, _22724_);
  or _73750_ (_22727_, _22726_, _03729_);
  or _73751_ (_22728_, _22710_, _03737_);
  and _73752_ (_22730_, _22728_, _03736_);
  and _73753_ (_22731_, _22730_, _22727_);
  and _73754_ (_22732_, _12641_, _05929_);
  or _73755_ (_22733_, _22732_, _22719_);
  and _73756_ (_22734_, _22733_, _03714_);
  or _73757_ (_22735_, _22734_, _03719_);
  or _73758_ (_22736_, _22735_, _22731_);
  or _73759_ (_22737_, _22719_, _12648_);
  and _73760_ (_22738_, _22737_, _22721_);
  or _73761_ (_22739_, _22738_, _06840_);
  and _73762_ (_22741_, _22739_, _03710_);
  and _73763_ (_22742_, _22741_, _22736_);
  and _73764_ (_22743_, _20391_, _05929_);
  or _73765_ (_22744_, _22743_, _22719_);
  and _73766_ (_22745_, _22744_, _03505_);
  or _73767_ (_22746_, _22745_, _07390_);
  or _73768_ (_22747_, _22746_, _22742_);
  and _73769_ (_22748_, _22747_, _22704_);
  or _73770_ (_22749_, _22748_, _04481_);
  and _73771_ (_22750_, _06592_, _05239_);
  or _73772_ (_22752_, _22701_, _07400_);
  or _73773_ (_22753_, _22752_, _22750_);
  and _73774_ (_22754_, _22753_, _03589_);
  and _73775_ (_22755_, _22754_, _22749_);
  and _73776_ (_22756_, _20416_, _05239_);
  or _73777_ (_22757_, _22701_, _22756_);
  and _73778_ (_22758_, _22757_, _03222_);
  or _73779_ (_22759_, _22758_, _22755_);
  or _73780_ (_22760_, _22759_, _08828_);
  and _73781_ (_22761_, _12733_, _05239_);
  or _73782_ (_22763_, _22701_, _07766_);
  or _73783_ (_22764_, _22763_, _22761_);
  and _73784_ (_22765_, _05239_, _06276_);
  or _73785_ (_22766_, _22765_, _22701_);
  or _73786_ (_22767_, _22766_, _05886_);
  and _73787_ (_22768_, _22767_, _07778_);
  and _73788_ (_22769_, _22768_, _22764_);
  and _73789_ (_22770_, _22769_, _22760_);
  and _73790_ (_22771_, _12739_, _05239_);
  or _73791_ (_22772_, _22771_, _22701_);
  and _73792_ (_22774_, _22772_, _03780_);
  or _73793_ (_22775_, _22774_, _22770_);
  and _73794_ (_22776_, _22775_, _07777_);
  or _73795_ (_22777_, _22701_, _05567_);
  and _73796_ (_22778_, _22766_, _03622_);
  and _73797_ (_22779_, _22778_, _22777_);
  or _73798_ (_22780_, _22779_, _22776_);
  and _73799_ (_22781_, _22780_, _06828_);
  and _73800_ (_22782_, _22710_, _03790_);
  and _73801_ (_22783_, _22782_, _22777_);
  or _73802_ (_22785_, _22783_, _03624_);
  or _73803_ (_22786_, _22785_, _22781_);
  nor _73804_ (_22787_, _12732_, _09557_);
  or _73805_ (_22788_, _22701_, _07795_);
  or _73806_ (_22789_, _22788_, _22787_);
  and _73807_ (_22790_, _22789_, _07793_);
  and _73808_ (_22791_, _22790_, _22786_);
  nor _73809_ (_22792_, _12738_, _09557_);
  or _73810_ (_22793_, _22792_, _22701_);
  and _73811_ (_22794_, _22793_, _03785_);
  or _73812_ (_22796_, _22794_, _03815_);
  or _73813_ (_22797_, _22796_, _22791_);
  or _73814_ (_22798_, _22706_, _04246_);
  and _73815_ (_22799_, _22798_, _03823_);
  and _73816_ (_22800_, _22799_, _22797_);
  and _73817_ (_22801_, _22733_, _03453_);
  or _73818_ (_22802_, _22801_, _03447_);
  or _73819_ (_22803_, _22802_, _22800_);
  and _73820_ (_22804_, _12794_, _05239_);
  or _73821_ (_22805_, _22701_, _03514_);
  or _73822_ (_22807_, _22805_, _22804_);
  and _73823_ (_22808_, _22807_, _43000_);
  and _73824_ (_22809_, _22808_, _22803_);
  nor _73825_ (_22810_, \oc8051_golden_model_1.P3 [3], rst);
  nor _73826_ (_22811_, _22810_, _04794_);
  or _73827_ (_43564_, _22811_, _22809_);
  and _73828_ (_22812_, _09557_, \oc8051_golden_model_1.P3 [4]);
  nor _73829_ (_22813_, _05777_, _09557_);
  or _73830_ (_22814_, _22813_, _22812_);
  or _73831_ (_22815_, _22814_, _06838_);
  and _73832_ (_22817_, _22717_, \oc8051_golden_model_1.P3 [4]);
  and _73833_ (_22818_, _12827_, _05929_);
  or _73834_ (_22819_, _22818_, _22817_);
  and _73835_ (_22820_, _22819_, _03714_);
  nor _73836_ (_22821_, _12841_, _09557_);
  or _73837_ (_22822_, _22821_, _22812_);
  or _73838_ (_22823_, _22822_, _04081_);
  and _73839_ (_22824_, _05239_, \oc8051_golden_model_1.ACC [4]);
  or _73840_ (_22825_, _22824_, _22812_);
  and _73841_ (_22826_, _22825_, _04409_);
  and _73842_ (_22828_, _09029_, \oc8051_golden_model_1.P3 [4]);
  or _73843_ (_22829_, _22828_, _03610_);
  or _73844_ (_22830_, _22829_, _22826_);
  and _73845_ (_22831_, _22830_, _04055_);
  and _73846_ (_22832_, _22831_, _22823_);
  and _73847_ (_22833_, _12845_, _05929_);
  or _73848_ (_22834_, _22833_, _22817_);
  and _73849_ (_22835_, _22834_, _03715_);
  or _73850_ (_22836_, _22835_, _03723_);
  or _73851_ (_22837_, _22836_, _22832_);
  or _73852_ (_22839_, _22814_, _03996_);
  and _73853_ (_22840_, _22839_, _22837_);
  or _73854_ (_22841_, _22840_, _03729_);
  or _73855_ (_22842_, _22825_, _03737_);
  and _73856_ (_22843_, _22842_, _03736_);
  and _73857_ (_22844_, _22843_, _22841_);
  or _73858_ (_22845_, _22844_, _22820_);
  and _73859_ (_22846_, _22845_, _06840_);
  or _73860_ (_22847_, _22817_, _12860_);
  and _73861_ (_22848_, _22847_, _03719_);
  and _73862_ (_22850_, _22848_, _22834_);
  or _73863_ (_22851_, _22850_, _22846_);
  and _73864_ (_22852_, _22851_, _03710_);
  and _73865_ (_22853_, _20511_, _05929_);
  or _73866_ (_22854_, _22853_, _22817_);
  and _73867_ (_22855_, _22854_, _03505_);
  or _73868_ (_22856_, _22855_, _07390_);
  or _73869_ (_22857_, _22856_, _22852_);
  and _73870_ (_22858_, _22857_, _22815_);
  or _73871_ (_22859_, _22858_, _04481_);
  and _73872_ (_22861_, _06730_, _05239_);
  or _73873_ (_22862_, _22812_, _07400_);
  or _73874_ (_22863_, _22862_, _22861_);
  and _73875_ (_22864_, _22863_, _03589_);
  and _73876_ (_22865_, _22864_, _22859_);
  and _73877_ (_22866_, _20536_, _05239_);
  or _73878_ (_22867_, _22866_, _22812_);
  and _73879_ (_22868_, _22867_, _03222_);
  or _73880_ (_22869_, _22868_, _08828_);
  or _73881_ (_22870_, _22869_, _22865_);
  and _73882_ (_22872_, _12821_, _05239_);
  or _73883_ (_22873_, _22812_, _07766_);
  or _73884_ (_22874_, _22873_, _22872_);
  and _73885_ (_22875_, _06298_, _05239_);
  or _73886_ (_22876_, _22875_, _22812_);
  or _73887_ (_22877_, _22876_, _05886_);
  and _73888_ (_22878_, _22877_, _07778_);
  and _73889_ (_22879_, _22878_, _22874_);
  and _73890_ (_22880_, _22879_, _22870_);
  and _73891_ (_22881_, _12817_, _05239_);
  or _73892_ (_22883_, _22881_, _22812_);
  and _73893_ (_22884_, _22883_, _03780_);
  or _73894_ (_22885_, _22884_, _22880_);
  and _73895_ (_22886_, _22885_, _07777_);
  or _73896_ (_22887_, _22812_, _05825_);
  and _73897_ (_22888_, _22876_, _03622_);
  and _73898_ (_22889_, _22888_, _22887_);
  or _73899_ (_22890_, _22889_, _22886_);
  and _73900_ (_22891_, _22890_, _06828_);
  and _73901_ (_22892_, _22825_, _03790_);
  and _73902_ (_22894_, _22892_, _22887_);
  or _73903_ (_22895_, _22894_, _03624_);
  or _73904_ (_22896_, _22895_, _22891_);
  nor _73905_ (_22897_, _12819_, _09557_);
  or _73906_ (_22898_, _22812_, _07795_);
  or _73907_ (_22899_, _22898_, _22897_);
  and _73908_ (_22900_, _22899_, _07793_);
  and _73909_ (_22901_, _22900_, _22896_);
  nor _73910_ (_22902_, _12816_, _09557_);
  or _73911_ (_22903_, _22902_, _22812_);
  and _73912_ (_22905_, _22903_, _03785_);
  or _73913_ (_22906_, _22905_, _03815_);
  or _73914_ (_22907_, _22906_, _22901_);
  or _73915_ (_22908_, _22822_, _04246_);
  and _73916_ (_22909_, _22908_, _03823_);
  and _73917_ (_22910_, _22909_, _22907_);
  and _73918_ (_22911_, _22819_, _03453_);
  or _73919_ (_22912_, _22911_, _03447_);
  or _73920_ (_22913_, _22912_, _22910_);
  and _73921_ (_22914_, _13003_, _05239_);
  or _73922_ (_22916_, _22812_, _03514_);
  or _73923_ (_22917_, _22916_, _22914_);
  and _73924_ (_22918_, _22917_, _43000_);
  and _73925_ (_22919_, _22918_, _22913_);
  nor _73926_ (_22920_, \oc8051_golden_model_1.P3 [4], rst);
  nor _73927_ (_22921_, _22920_, _04794_);
  or _73928_ (_43565_, _22921_, _22919_);
  nor _73929_ (_22922_, \oc8051_golden_model_1.P3 [5], rst);
  nor _73930_ (_22923_, _22922_, _04794_);
  and _73931_ (_22924_, _09557_, \oc8051_golden_model_1.P3 [5]);
  nor _73932_ (_22926_, _13014_, _09557_);
  or _73933_ (_22927_, _22926_, _22924_);
  or _73934_ (_22928_, _22927_, _04081_);
  and _73935_ (_22929_, _05239_, \oc8051_golden_model_1.ACC [5]);
  or _73936_ (_22930_, _22929_, _22924_);
  and _73937_ (_22931_, _22930_, _04409_);
  and _73938_ (_22932_, _09029_, \oc8051_golden_model_1.P3 [5]);
  or _73939_ (_22933_, _22932_, _03610_);
  or _73940_ (_22934_, _22933_, _22931_);
  and _73941_ (_22935_, _22934_, _04055_);
  and _73942_ (_22937_, _22935_, _22928_);
  and _73943_ (_22938_, _22717_, \oc8051_golden_model_1.P3 [5]);
  and _73944_ (_22939_, _13037_, _05929_);
  or _73945_ (_22940_, _22939_, _22938_);
  and _73946_ (_22941_, _22940_, _03715_);
  or _73947_ (_22942_, _22941_, _03723_);
  or _73948_ (_22943_, _22942_, _22937_);
  nor _73949_ (_22944_, _05469_, _09557_);
  or _73950_ (_22945_, _22944_, _22924_);
  or _73951_ (_22946_, _22945_, _03996_);
  and _73952_ (_22948_, _22946_, _22943_);
  or _73953_ (_22949_, _22948_, _03729_);
  or _73954_ (_22950_, _22930_, _03737_);
  and _73955_ (_22951_, _22950_, _03736_);
  and _73956_ (_22952_, _22951_, _22949_);
  and _73957_ (_22953_, _13047_, _05929_);
  or _73958_ (_22954_, _22953_, _22938_);
  and _73959_ (_22955_, _22954_, _03714_);
  or _73960_ (_22956_, _22955_, _03719_);
  or _73961_ (_22957_, _22956_, _22952_);
  or _73962_ (_22959_, _22938_, _13054_);
  and _73963_ (_22960_, _22959_, _22940_);
  or _73964_ (_22961_, _22960_, _06840_);
  and _73965_ (_22962_, _22961_, _03710_);
  and _73966_ (_22963_, _22962_, _22957_);
  and _73967_ (_22964_, _20633_, _05929_);
  or _73968_ (_22965_, _22964_, _22938_);
  and _73969_ (_22966_, _22965_, _03505_);
  or _73970_ (_22967_, _22966_, _07390_);
  or _73971_ (_22968_, _22967_, _22963_);
  or _73972_ (_22970_, _22945_, _06838_);
  and _73973_ (_22971_, _22970_, _22968_);
  or _73974_ (_22972_, _22971_, _04481_);
  and _73975_ (_22973_, _06684_, _05239_);
  or _73976_ (_22974_, _22924_, _07400_);
  or _73977_ (_22975_, _22974_, _22973_);
  and _73978_ (_22976_, _22975_, _03589_);
  and _73979_ (_22977_, _22976_, _22972_);
  and _73980_ (_22978_, _20660_, _05239_);
  or _73981_ (_22979_, _22978_, _22924_);
  and _73982_ (_22981_, _22979_, _03222_);
  or _73983_ (_22982_, _22981_, _08828_);
  or _73984_ (_22983_, _22982_, _22977_);
  and _73985_ (_22984_, _13141_, _05239_);
  or _73986_ (_22985_, _22924_, _07766_);
  or _73987_ (_22986_, _22985_, _22984_);
  and _73988_ (_22987_, _06306_, _05239_);
  or _73989_ (_22988_, _22987_, _22924_);
  or _73990_ (_22989_, _22988_, _05886_);
  and _73991_ (_22990_, _22989_, _07778_);
  and _73992_ (_22991_, _22990_, _22986_);
  and _73993_ (_22992_, _22991_, _22983_);
  and _73994_ (_22993_, _13147_, _05239_);
  or _73995_ (_22994_, _22993_, _22924_);
  and _73996_ (_22995_, _22994_, _03780_);
  or _73997_ (_22996_, _22995_, _22992_);
  and _73998_ (_22997_, _22996_, _07777_);
  or _73999_ (_22998_, _22924_, _05518_);
  and _74000_ (_22999_, _22988_, _03622_);
  and _74001_ (_23000_, _22999_, _22998_);
  or _74002_ (_23003_, _23000_, _22997_);
  and _74003_ (_23004_, _23003_, _06828_);
  and _74004_ (_23005_, _22930_, _03790_);
  and _74005_ (_23006_, _23005_, _22998_);
  or _74006_ (_23007_, _23006_, _03624_);
  or _74007_ (_23008_, _23007_, _23004_);
  nor _74008_ (_23009_, _13140_, _09557_);
  or _74009_ (_23010_, _22924_, _07795_);
  or _74010_ (_23011_, _23010_, _23009_);
  and _74011_ (_23012_, _23011_, _07793_);
  and _74012_ (_23014_, _23012_, _23008_);
  nor _74013_ (_23015_, _13146_, _09557_);
  or _74014_ (_23016_, _23015_, _22924_);
  and _74015_ (_23017_, _23016_, _03785_);
  or _74016_ (_23018_, _23017_, _03815_);
  or _74017_ (_23019_, _23018_, _23014_);
  or _74018_ (_23020_, _22927_, _04246_);
  and _74019_ (_23021_, _23020_, _03823_);
  and _74020_ (_23022_, _23021_, _23019_);
  and _74021_ (_23023_, _22954_, _03453_);
  or _74022_ (_23024_, _23023_, _03447_);
  or _74023_ (_23025_, _23024_, _23022_);
  and _74024_ (_23026_, _13199_, _05239_);
  or _74025_ (_23027_, _22924_, _03514_);
  or _74026_ (_23028_, _23027_, _23026_);
  and _74027_ (_23029_, _23028_, _43000_);
  and _74028_ (_23030_, _23029_, _23025_);
  or _74029_ (_43566_, _23030_, _22923_);
  not _74030_ (_23031_, \oc8051_golden_model_1.P3 [6]);
  nor _74031_ (_23032_, _05239_, _23031_);
  nor _74032_ (_23035_, _13242_, _09557_);
  or _74033_ (_23036_, _23035_, _23032_);
  or _74034_ (_23037_, _23036_, _04081_);
  and _74035_ (_23038_, _05239_, \oc8051_golden_model_1.ACC [6]);
  or _74036_ (_23039_, _23038_, _23032_);
  and _74037_ (_23040_, _23039_, _04409_);
  nor _74038_ (_23041_, _04409_, _23031_);
  or _74039_ (_23042_, _23041_, _03610_);
  or _74040_ (_23043_, _23042_, _23040_);
  and _74041_ (_23044_, _23043_, _04055_);
  and _74042_ (_23046_, _23044_, _23037_);
  nor _74043_ (_23047_, _05929_, _23031_);
  and _74044_ (_23048_, _13229_, _05929_);
  or _74045_ (_23049_, _23048_, _23047_);
  and _74046_ (_23050_, _23049_, _03715_);
  or _74047_ (_23051_, _23050_, _03723_);
  or _74048_ (_23052_, _23051_, _23046_);
  nor _74049_ (_23053_, _05363_, _09557_);
  or _74050_ (_23054_, _23053_, _23032_);
  or _74051_ (_23055_, _23054_, _03996_);
  and _74052_ (_23056_, _23055_, _23052_);
  or _74053_ (_23057_, _23056_, _03729_);
  or _74054_ (_23058_, _23039_, _03737_);
  and _74055_ (_23059_, _23058_, _03736_);
  and _74056_ (_23060_, _23059_, _23057_);
  and _74057_ (_23061_, _13253_, _05929_);
  or _74058_ (_23062_, _23061_, _23047_);
  and _74059_ (_23063_, _23062_, _03714_);
  or _74060_ (_23064_, _23063_, _03719_);
  or _74061_ (_23065_, _23064_, _23060_);
  or _74062_ (_23068_, _23047_, _13260_);
  and _74063_ (_23069_, _23068_, _23049_);
  or _74064_ (_23070_, _23069_, _06840_);
  and _74065_ (_23071_, _23070_, _03710_);
  and _74066_ (_23072_, _23071_, _23065_);
  and _74067_ (_23073_, _20753_, _05929_);
  or _74068_ (_23074_, _23073_, _23047_);
  and _74069_ (_23075_, _23074_, _03505_);
  or _74070_ (_23076_, _23075_, _07390_);
  or _74071_ (_23077_, _23076_, _23072_);
  or _74072_ (_23079_, _23054_, _06838_);
  and _74073_ (_23080_, _23079_, _23077_);
  or _74074_ (_23081_, _23080_, _04481_);
  and _74075_ (_23082_, _06455_, _05239_);
  or _74076_ (_23083_, _23032_, _07400_);
  or _74077_ (_23084_, _23083_, _23082_);
  and _74078_ (_23085_, _23084_, _03589_);
  and _74079_ (_23086_, _23085_, _23081_);
  and _74080_ (_23087_, _20778_, _05239_);
  or _74081_ (_23088_, _23087_, _23032_);
  and _74082_ (_23089_, _23088_, _03222_);
  or _74083_ (_23090_, _23089_, _08828_);
  or _74084_ (_23091_, _23090_, _23086_);
  and _74085_ (_23092_, _13347_, _05239_);
  or _74086_ (_23093_, _23032_, _07766_);
  or _74087_ (_23094_, _23093_, _23092_);
  and _74088_ (_23095_, _13339_, _05239_);
  or _74089_ (_23096_, _23095_, _23032_);
  or _74090_ (_23097_, _23096_, _05886_);
  and _74091_ (_23098_, _23097_, _07778_);
  and _74092_ (_23101_, _23098_, _23094_);
  and _74093_ (_23102_, _23101_, _23091_);
  and _74094_ (_23103_, _13353_, _05239_);
  or _74095_ (_23104_, _23103_, _23032_);
  and _74096_ (_23105_, _23104_, _03780_);
  or _74097_ (_23106_, _23105_, _23102_);
  and _74098_ (_23107_, _23106_, _07777_);
  or _74099_ (_23108_, _23032_, _05412_);
  and _74100_ (_23109_, _23096_, _03622_);
  and _74101_ (_23110_, _23109_, _23108_);
  or _74102_ (_23112_, _23110_, _23107_);
  and _74103_ (_23113_, _23112_, _06828_);
  and _74104_ (_23114_, _23039_, _03790_);
  and _74105_ (_23115_, _23114_, _23108_);
  or _74106_ (_23116_, _23115_, _03624_);
  or _74107_ (_23117_, _23116_, _23113_);
  nor _74108_ (_23118_, _13346_, _09557_);
  or _74109_ (_23119_, _23032_, _07795_);
  or _74110_ (_23120_, _23119_, _23118_);
  and _74111_ (_23121_, _23120_, _07793_);
  and _74112_ (_23122_, _23121_, _23117_);
  nor _74113_ (_23123_, _13352_, _09557_);
  or _74114_ (_23124_, _23123_, _23032_);
  and _74115_ (_23125_, _23124_, _03785_);
  or _74116_ (_23126_, _23125_, _03815_);
  or _74117_ (_23127_, _23126_, _23122_);
  or _74118_ (_23128_, _23036_, _04246_);
  and _74119_ (_23129_, _23128_, _03823_);
  and _74120_ (_23130_, _23129_, _23127_);
  and _74121_ (_23131_, _23062_, _03453_);
  or _74122_ (_23134_, _23131_, _03447_);
  or _74123_ (_23135_, _23134_, _23130_);
  and _74124_ (_23136_, _13402_, _05239_);
  or _74125_ (_23137_, _23032_, _03514_);
  or _74126_ (_23138_, _23137_, _23136_);
  and _74127_ (_23139_, _23138_, _43000_);
  and _74128_ (_23140_, _23139_, _23135_);
  nor _74129_ (_23141_, _43000_, _23031_);
  or _74130_ (_23142_, _23141_, rst);
  or _74131_ (_43567_, _23142_, _23140_);
  and _74132_ (_23144_, _43004_, \oc8051_golden_model_1.PSW [0]);
  not _74133_ (_23145_, _15783_);
  nor _74134_ (_23146_, _16424_, _23145_);
  and _74135_ (_23147_, _16424_, _23145_);
  nor _74136_ (_23148_, _23147_, _23146_);
  nor _74137_ (_23149_, _23148_, _17075_);
  and _74138_ (_23150_, _23148_, _17075_);
  nor _74139_ (_23151_, _23150_, _23149_);
  not _74140_ (_23152_, _23151_);
  nor _74141_ (_23153_, _15460_, _14988_);
  and _74142_ (_23154_, _15460_, _14988_);
  nor _74143_ (_23155_, _23154_, _23153_);
  and _74144_ (_23156_, _23155_, _16105_);
  nor _74145_ (_23157_, _23155_, _16105_);
  nor _74146_ (_23158_, _23157_, _23156_);
  and _74147_ (_23159_, _23158_, _16761_);
  nor _74148_ (_23160_, _23158_, _16761_);
  or _74149_ (_23161_, _23160_, _23159_);
  and _74150_ (_23162_, _23161_, _08801_);
  nor _74151_ (_23163_, _23161_, _08801_);
  or _74152_ (_23166_, _23163_, _23162_);
  nand _74153_ (_23167_, _23166_, _23152_);
  or _74154_ (_23168_, _23166_, _23152_);
  and _74155_ (_23169_, _23168_, _03447_);
  and _74156_ (_23170_, _23169_, _23167_);
  not _74157_ (_23171_, _15529_);
  nor _74158_ (_23172_, _15263_, _14957_);
  and _74159_ (_23173_, _15263_, _14957_);
  nor _74160_ (_23174_, _23173_, _23172_);
  nor _74161_ (_23175_, _23174_, _23171_);
  and _74162_ (_23177_, _23174_, _23171_);
  or _74163_ (_23178_, _23177_, _23175_);
  and _74164_ (_23179_, _23178_, _15888_);
  nor _74165_ (_23180_, _23178_, _15888_);
  or _74166_ (_23181_, _23180_, _23179_);
  and _74167_ (_23182_, _23181_, _16199_);
  nor _74168_ (_23183_, _23181_, _16199_);
  or _74169_ (_23184_, _23183_, _23182_);
  and _74170_ (_23185_, _23184_, _16529_);
  nor _74171_ (_23186_, _23184_, _16529_);
  or _74172_ (_23187_, _23186_, _23185_);
  and _74173_ (_23188_, _23187_, _16862_);
  nor _74174_ (_23189_, _23187_, _16862_);
  or _74175_ (_23190_, _23189_, _23188_);
  and _74176_ (_23191_, _23190_, _08140_);
  nor _74177_ (_23192_, _23190_, _08140_);
  or _74178_ (_23193_, _23192_, _23191_);
  and _74179_ (_23194_, _23193_, _03453_);
  nor _74180_ (_23195_, _07525_, _07524_);
  nor _74181_ (_23196_, _23195_, _07433_);
  and _74182_ (_23199_, _23195_, _07433_);
  nor _74183_ (_23200_, _23199_, _23196_);
  nor _74184_ (_23201_, _07449_, _07448_);
  nor _74185_ (_23202_, _23201_, _15450_);
  and _74186_ (_23203_, _23201_, _15450_);
  nor _74187_ (_23204_, _23203_, _23202_);
  and _74188_ (_23205_, _23204_, _23200_);
  nor _74189_ (_23206_, _23204_, _23200_);
  nor _74190_ (_23207_, _23206_, _23205_);
  or _74191_ (_23208_, _23207_, _06075_);
  nand _74192_ (_23210_, _23207_, _06075_);
  and _74193_ (_23211_, _23210_, _23208_);
  nor _74194_ (_23212_, _03628_, _03203_);
  and _74195_ (_23213_, _23212_, _08733_);
  nor _74196_ (_23214_, _03972_, _03515_);
  and _74197_ (_23215_, _23214_, _23213_);
  nor _74198_ (_23216_, _04803_, _03491_);
  and _74199_ (_23217_, _23216_, _06409_);
  and _74200_ (_23218_, _23217_, _23215_);
  or _74201_ (_23219_, _23218_, _23211_);
  nor _74202_ (_23221_, _15279_, _15278_);
  nor _74203_ (_23222_, _15503_, \oc8051_golden_model_1.ACC [3]);
  and _74204_ (_23223_, _15503_, \oc8051_golden_model_1.ACC [3]);
  nor _74205_ (_23224_, _23223_, _23222_);
  nor _74206_ (_23225_, _23201_, \oc8051_golden_model_1.ACC [6]);
  and _74207_ (_23226_, _23201_, \oc8051_golden_model_1.ACC [6]);
  nor _74208_ (_23227_, _23226_, _23225_);
  and _74209_ (_23228_, _23227_, _23224_);
  nor _74210_ (_23229_, _23227_, _23224_);
  nor _74211_ (_23230_, _23229_, _23228_);
  nor _74212_ (_23232_, _23230_, _23221_);
  and _74213_ (_23233_, _23230_, _23221_);
  or _74214_ (_23234_, _23233_, _23232_);
  and _74215_ (_23235_, _23234_, _08587_);
  not _74216_ (_23236_, _06377_);
  nor _74217_ (_23237_, _12332_, _12003_);
  and _74218_ (_23238_, _12332_, _12003_);
  nor _74219_ (_23239_, _23238_, _23237_);
  and _74220_ (_23240_, _23239_, _12538_);
  nor _74221_ (_23241_, _23239_, _12538_);
  or _74222_ (_23243_, _23241_, _23240_);
  nand _74223_ (_23244_, _23243_, _12738_);
  or _74224_ (_23245_, _23243_, _12738_);
  and _74225_ (_23246_, _23245_, _23244_);
  nor _74226_ (_23247_, _13146_, _12816_);
  and _74227_ (_23248_, _13146_, _12816_);
  nor _74228_ (_23249_, _23248_, _23247_);
  nor _74229_ (_23250_, _23249_, _13352_);
  and _74230_ (_23251_, _23249_, _13352_);
  nor _74231_ (_23252_, _23251_, _23250_);
  not _74232_ (_23254_, _23252_);
  nor _74233_ (_23255_, _23254_, _23246_);
  and _74234_ (_23256_, _23254_, _23246_);
  nor _74235_ (_23257_, _23256_, _23255_);
  nor _74236_ (_23258_, _23257_, _23236_);
  and _74237_ (_23259_, _23257_, _23236_);
  or _74238_ (_23260_, _23259_, _23258_);
  and _74239_ (_23261_, _23260_, _03783_);
  nor _74240_ (_23262_, _04749_, _04722_);
  and _74241_ (_23263_, _23262_, _11707_);
  or _74242_ (_23265_, _23263_, _23211_);
  not _74243_ (_23266_, _03613_);
  and _74244_ (_23267_, _11671_, _23266_);
  and _74245_ (_23268_, _23267_, _03598_);
  or _74246_ (_23269_, _23268_, _23211_);
  nor _74247_ (_23270_, _06787_, _06638_);
  not _74248_ (_23271_, _23270_);
  nand _74249_ (_23272_, _23271_, _12203_);
  or _74250_ (_23273_, _23271_, _12203_);
  and _74251_ (_23274_, _23273_, _23272_);
  nor _74252_ (_23276_, _06789_, _06731_);
  nand _74253_ (_23277_, _23276_, _06456_);
  or _74254_ (_23278_, _23276_, _06456_);
  and _74255_ (_23279_, _23278_, _23277_);
  and _74256_ (_23280_, _23279_, _23274_);
  nor _74257_ (_23281_, _23279_, _23274_);
  or _74258_ (_23282_, _23281_, _23280_);
  nor _74259_ (_23283_, _23282_, _06069_);
  and _74260_ (_23284_, _23282_, _06069_);
  or _74261_ (_23285_, _23284_, _23283_);
  or _74262_ (_23287_, _23285_, _08067_);
  and _74263_ (_23288_, _06772_, _05469_);
  nor _74264_ (_23289_, _06772_, _05469_);
  nor _74265_ (_23290_, _23289_, _23288_);
  and _74266_ (_23291_, _12205_, _05777_);
  nor _74267_ (_23292_, _12205_, _05777_);
  nor _74268_ (_23293_, _23292_, _23291_);
  nor _74269_ (_23294_, _06766_, _05836_);
  nor _74270_ (_23295_, _23294_, _23293_);
  and _74271_ (_23296_, _23294_, _23293_);
  nor _74272_ (_23298_, _23296_, _23295_);
  or _74273_ (_23299_, _23298_, _23290_);
  nand _74274_ (_23300_, _23298_, _23290_);
  and _74275_ (_23301_, _23300_, _23299_);
  and _74276_ (_23302_, _23301_, _08079_);
  nor _74277_ (_23303_, _04729_, _03981_);
  and _74278_ (_23304_, _23303_, \oc8051_golden_model_1.PSW [0]);
  not _74279_ (_23305_, _23303_);
  and _74280_ (_23306_, _23305_, _23211_);
  or _74281_ (_23307_, _23306_, _23304_);
  and _74282_ (_23309_, _23307_, _08078_);
  or _74283_ (_23310_, _23309_, _08066_);
  or _74284_ (_23311_, _23310_, _23302_);
  and _74285_ (_23312_, _06072_, _03235_);
  and _74286_ (_23313_, _23312_, _23311_);
  and _74287_ (_23314_, _23313_, _23287_);
  and _74288_ (_23315_, _23211_, _06073_);
  or _74289_ (_23316_, _23315_, _04422_);
  or _74290_ (_23317_, _23316_, _23314_);
  nor _74291_ (_23318_, _23227_, \oc8051_golden_model_1.ACC [7]);
  and _74292_ (_23320_, _23227_, \oc8051_golden_model_1.ACC [7]);
  nor _74293_ (_23321_, _23320_, _23318_);
  nor _74294_ (_23322_, _23321_, _23274_);
  and _74295_ (_23323_, _23321_, _23274_);
  or _74296_ (_23324_, _23323_, _23322_);
  or _74297_ (_23325_, _23324_, _05966_);
  and _74298_ (_23326_, _23325_, _04081_);
  and _74299_ (_23327_, _23326_, _23317_);
  not _74300_ (_23328_, _16816_);
  not _74301_ (_23329_, _14988_);
  nor _74302_ (_23331_, _15232_, _23329_);
  and _74303_ (_23332_, _15232_, _23329_);
  nor _74304_ (_23333_, _23332_, _23331_);
  and _74305_ (_23334_, _23333_, _15497_);
  nor _74306_ (_23335_, _23333_, _15497_);
  nor _74307_ (_23336_, _23335_, _23334_);
  and _74308_ (_23337_, _23336_, _16497_);
  nor _74309_ (_23338_, _23336_, _16497_);
  or _74310_ (_23339_, _23338_, _23337_);
  nor _74311_ (_23340_, _16167_, _15855_);
  and _74312_ (_23342_, _16167_, _15855_);
  nor _74313_ (_23343_, _23342_, _23340_);
  and _74314_ (_23344_, _23343_, _23339_);
  nor _74315_ (_23345_, _23343_, _23339_);
  nor _74316_ (_23346_, _23345_, _23344_);
  nor _74317_ (_23347_, _23346_, _23328_);
  and _74318_ (_23348_, _23346_, _23328_);
  or _74319_ (_23349_, _23348_, _23347_);
  and _74320_ (_23350_, _23349_, _08091_);
  nor _74321_ (_23351_, _23349_, _08091_);
  or _74322_ (_23352_, _23351_, _23350_);
  and _74323_ (_23353_, _23352_, _03610_);
  or _74324_ (_23354_, _23353_, _08089_);
  or _74325_ (_23355_, _23354_, _23327_);
  and _74326_ (_23356_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor _74327_ (_23357_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or _74328_ (_23358_, _23357_, _23356_);
  and _74329_ (_23359_, _23358_, _15238_);
  nor _74330_ (_23360_, _23358_, _15238_);
  nor _74331_ (_23361_, _23360_, _23359_);
  nor _74332_ (_23363_, _15861_, _07484_);
  and _74333_ (_23364_, _15861_, _07484_);
  nor _74334_ (_23365_, _23364_, _23363_);
  and _74335_ (_23366_, _23365_, _23361_);
  nor _74336_ (_23367_, _23365_, _23361_);
  nor _74337_ (_23368_, _23367_, _23366_);
  nor _74338_ (_23369_, _23368_, _16504_);
  and _74339_ (_23370_, _23368_, _16504_);
  or _74340_ (_23371_, _23370_, _23369_);
  nor _74341_ (_23372_, _16835_, _08114_);
  and _74342_ (_23374_, _16835_, _08114_);
  nor _74343_ (_23375_, _23374_, _23372_);
  nor _74344_ (_23376_, _23375_, _23371_);
  and _74345_ (_23377_, _23375_, _23371_);
  or _74346_ (_23378_, _23377_, _09882_);
  or _74347_ (_23379_, _23378_, _23376_);
  and _74348_ (_23380_, _23379_, _23355_);
  or _74349_ (_23381_, _23380_, _09895_);
  or _74350_ (_23382_, _23211_, _09896_);
  and _74351_ (_23383_, _23382_, _04055_);
  and _74352_ (_23384_, _23383_, _23381_);
  and _74353_ (_23385_, _15245_, _14994_);
  nor _74354_ (_23386_, _15245_, _14994_);
  or _74355_ (_23387_, _23386_, _23385_);
  nor _74356_ (_23388_, _16841_, _16179_);
  and _74357_ (_23389_, _16841_, _16179_);
  nor _74358_ (_23390_, _23389_, _23388_);
  nor _74359_ (_23391_, _23390_, _23387_);
  and _74360_ (_23392_, _23390_, _23387_);
  or _74361_ (_23393_, _23392_, _23391_);
  not _74362_ (_23394_, _16508_);
  nor _74363_ (_23395_, _15867_, _15511_);
  and _74364_ (_23396_, _15867_, _15511_);
  nor _74365_ (_23397_, _23396_, _23395_);
  nor _74366_ (_23398_, _23397_, _23394_);
  and _74367_ (_23399_, _23397_, _23394_);
  nor _74368_ (_23400_, _23399_, _23398_);
  and _74369_ (_23401_, _23400_, _23393_);
  nor _74370_ (_23402_, _23400_, _23393_);
  nor _74371_ (_23403_, _23402_, _23401_);
  and _74372_ (_23404_, _23403_, _08120_);
  nor _74373_ (_23405_, _23403_, _08120_);
  or _74374_ (_23406_, _23405_, _23404_);
  and _74375_ (_23407_, _23406_, _03715_);
  or _74376_ (_23408_, _23407_, _23384_);
  and _74377_ (_23409_, _23408_, _03230_);
  and _74378_ (_23410_, _23211_, _04768_);
  or _74379_ (_23411_, _23410_, _23409_);
  or _74380_ (_23412_, _23411_, _03723_);
  and _74381_ (_23413_, _15213_, _14971_);
  nor _74382_ (_23414_, _15213_, _14971_);
  nor _74383_ (_23415_, _23414_, _23413_);
  and _74384_ (_23416_, _23415_, _15481_);
  nor _74385_ (_23417_, _23415_, _15481_);
  or _74386_ (_23418_, _23417_, _23416_);
  and _74387_ (_23419_, _23418_, _15818_);
  nor _74388_ (_23420_, _23418_, _15818_);
  or _74389_ (_23421_, _23420_, _23419_);
  and _74390_ (_23422_, _23421_, _16131_);
  nor _74391_ (_23423_, _23421_, _16131_);
  or _74392_ (_23424_, _23423_, _23422_);
  and _74393_ (_23425_, _23424_, _16461_);
  nor _74394_ (_23426_, _23424_, _16461_);
  or _74395_ (_23427_, _23426_, _23425_);
  and _74396_ (_23428_, _23427_, _16793_);
  nor _74397_ (_23429_, _23427_, _16793_);
  or _74398_ (_23430_, _23429_, _23428_);
  and _74399_ (_23431_, _23430_, _07910_);
  nor _74400_ (_23432_, _23430_, _07910_);
  or _74401_ (_23433_, _23432_, _23431_);
  or _74402_ (_23435_, _23433_, _03996_);
  and _74403_ (_23436_, _23435_, _08062_);
  and _74404_ (_23437_, _23436_, _23412_);
  not _74405_ (_23438_, _08062_);
  and _74406_ (_23439_, _23301_, _23438_);
  or _74407_ (_23440_, _23439_, _23437_);
  and _74408_ (_23441_, _23440_, _08061_);
  and _74409_ (_23442_, _23301_, _04759_);
  or _74410_ (_23443_, _23442_, _04443_);
  or _74411_ (_23444_, _23443_, _23441_);
  or _74412_ (_23446_, _23285_, _08128_);
  and _74413_ (_23447_, _23446_, _03737_);
  and _74414_ (_23448_, _23447_, _23444_);
  not _74415_ (_23449_, _08285_);
  nor _74416_ (_23450_, _08271_, _08260_);
  and _74417_ (_23451_, _08271_, _08260_);
  nor _74418_ (_23452_, _23451_, _23450_);
  nor _74419_ (_23453_, _23452_, _23449_);
  and _74420_ (_23454_, _23452_, _23449_);
  nor _74421_ (_23455_, _23454_, _23453_);
  and _74422_ (_23456_, _08235_, _08218_);
  nor _74423_ (_23457_, _23456_, _08517_);
  and _74424_ (_23458_, _08248_, _08203_);
  nor _74425_ (_23459_, _08248_, _08203_);
  or _74426_ (_23460_, _23459_, _23458_);
  and _74427_ (_23461_, _23460_, _23457_);
  nor _74428_ (_23462_, _23460_, _23457_);
  nor _74429_ (_23463_, _23462_, _23461_);
  nor _74430_ (_23464_, _23463_, _23455_);
  and _74431_ (_23465_, _23463_, _23455_);
  nor _74432_ (_23467_, _23465_, _23464_);
  or _74433_ (_23468_, _23467_, _06133_);
  nand _74434_ (_23469_, _23467_, _06133_);
  and _74435_ (_23470_, _23469_, _03729_);
  and _74436_ (_23471_, _23470_, _23468_);
  or _74437_ (_23472_, _23471_, _11668_);
  or _74438_ (_23473_, _23472_, _23448_);
  or _74439_ (_23474_, _23211_, _11666_);
  and _74440_ (_23475_, _23474_, _03736_);
  and _74441_ (_23476_, _23475_, _23473_);
  nand _74442_ (_23478_, _23193_, _03714_);
  nand _74443_ (_23479_, _23478_, _23268_);
  or _74444_ (_23480_, _23479_, _23476_);
  nand _74445_ (_23481_, _23480_, _23269_);
  not _74446_ (_23482_, _03606_);
  and _74447_ (_23483_, _03618_, _23482_);
  and _74448_ (_23484_, _23483_, _09856_);
  and _74449_ (_23485_, _11358_, _23484_);
  nand _74450_ (_23486_, _23485_, _23481_);
  or _74451_ (_23487_, _23485_, _23211_);
  and _74452_ (_23489_, _23487_, _06840_);
  and _74453_ (_23490_, _23489_, _23486_);
  nor _74454_ (_23491_, _15837_, _23329_);
  and _74455_ (_23492_, _15837_, _23329_);
  nor _74456_ (_23493_, _23492_, _23491_);
  and _74457_ (_23494_, _23493_, _16204_);
  nor _74458_ (_23495_, _23493_, _16204_);
  nor _74459_ (_23496_, _23495_, _23494_);
  nor _74460_ (_23497_, _16868_, _08145_);
  and _74461_ (_23498_, _16868_, _08145_);
  nor _74462_ (_23500_, _23498_, _23497_);
  not _74463_ (_23501_, _23500_);
  nor _74464_ (_23502_, _23501_, _23496_);
  and _74465_ (_23503_, _23501_, _23496_);
  nor _74466_ (_23504_, _23503_, _23502_);
  not _74467_ (_23505_, _15534_);
  and _74468_ (_23506_, _23505_, _15268_);
  nor _74469_ (_23507_, _23505_, _15268_);
  nor _74470_ (_23508_, _23507_, _23506_);
  and _74471_ (_23509_, _23508_, _16482_);
  nor _74472_ (_23510_, _23508_, _16482_);
  or _74473_ (_23511_, _23510_, _23509_);
  nand _74474_ (_23512_, _23511_, _23504_);
  or _74475_ (_23513_, _23511_, _23504_);
  and _74476_ (_23514_, _23513_, _03719_);
  nand _74477_ (_23515_, _23514_, _23512_);
  nand _74478_ (_23516_, _23515_, _23263_);
  or _74479_ (_23517_, _23516_, _23490_);
  nand _74480_ (_23518_, _23517_, _23265_);
  nor _74481_ (_23519_, _04463_, _04753_);
  and _74482_ (_23521_, _23519_, _11353_);
  nand _74483_ (_23522_, _23521_, _23518_);
  or _74484_ (_23523_, _23521_, _23211_);
  and _74485_ (_23524_, _23523_, _06875_);
  and _74486_ (_23525_, _23524_, _23522_);
  nor _74487_ (_23526_, _03753_, _11727_);
  and _74488_ (_23527_, _23526_, _08848_);
  nor _74489_ (_23528_, _15274_, _15020_);
  and _74490_ (_23529_, _15274_, _15020_);
  or _74491_ (_23530_, _23529_, _23528_);
  nor _74492_ (_23532_, _23530_, _15539_);
  and _74493_ (_23533_, _23530_, _15539_);
  nor _74494_ (_23534_, _23533_, _23532_);
  nor _74495_ (_23535_, _23534_, _15895_);
  and _74496_ (_23536_, _23534_, _15895_);
  nor _74497_ (_23537_, _23536_, _23535_);
  not _74498_ (_23538_, _23537_);
  nor _74499_ (_23539_, _23538_, _16210_);
  and _74500_ (_23540_, _23538_, _16210_);
  nor _74501_ (_23541_, _23540_, _23539_);
  nor _74502_ (_23543_, _23541_, _16537_);
  and _74503_ (_23544_, _23541_, _16537_);
  or _74504_ (_23545_, _23544_, _23543_);
  and _74505_ (_23546_, _23545_, _16873_);
  nor _74506_ (_23547_, _23545_, _16873_);
  nor _74507_ (_23548_, _23547_, _23546_);
  or _74508_ (_23549_, _23548_, _08150_);
  nand _74509_ (_23550_, _23548_, _08150_);
  and _74510_ (_23551_, _23550_, _06869_);
  nand _74511_ (_23552_, _23551_, _23549_);
  nand _74512_ (_23554_, _23552_, _23527_);
  or _74513_ (_23555_, _23554_, _23525_);
  or _74514_ (_23556_, _23527_, _23211_);
  and _74515_ (_23557_, _23556_, _09668_);
  and _74516_ (_23558_, _23557_, _23555_);
  nand _74517_ (_23559_, _23211_, _03752_);
  nand _74518_ (_23560_, _23559_, _08059_);
  or _74519_ (_23561_, _23560_, _23558_);
  not _74520_ (_23562_, _08180_);
  nor _74521_ (_23563_, _15285_, _08170_);
  and _74522_ (_23565_, _15285_, _08170_);
  nor _74523_ (_23566_, _23565_, _23563_);
  or _74524_ (_23567_, _23566_, _15911_);
  nand _74525_ (_23568_, _23566_, _15911_);
  and _74526_ (_23569_, _23568_, _23567_);
  or _74527_ (_23570_, _23569_, _15557_);
  nand _74528_ (_23571_, _23569_, _15557_);
  and _74529_ (_23572_, _23571_, _23570_);
  nor _74530_ (_23573_, _23572_, _16229_);
  and _74531_ (_23574_, _23572_, _16229_);
  nor _74532_ (_23575_, _23574_, _23573_);
  nor _74533_ (_23576_, _23575_, _16554_);
  and _74534_ (_23577_, _23575_, _16554_);
  or _74535_ (_23578_, _23577_, _23576_);
  nor _74536_ (_23579_, _23578_, _16890_);
  and _74537_ (_23580_, _23578_, _16890_);
  nor _74538_ (_23581_, _23580_, _23579_);
  nor _74539_ (_23582_, _23581_, _23562_);
  and _74540_ (_23583_, _23581_, _23562_);
  or _74541_ (_23584_, _23583_, _23582_);
  or _74542_ (_23586_, _23584_, _08059_);
  and _74543_ (_23587_, _23586_, _23561_);
  or _74544_ (_23588_, _23587_, _08051_);
  nor _74545_ (_23589_, _15293_, _15029_);
  and _74546_ (_23590_, _15293_, _15029_);
  or _74547_ (_23591_, _23590_, _23589_);
  and _74548_ (_23592_, _23591_, _15573_);
  nor _74549_ (_23593_, _23591_, _15573_);
  or _74550_ (_23594_, _23593_, _23592_);
  nor _74551_ (_23595_, _23594_, _15930_);
  and _74552_ (_23597_, _23594_, _15930_);
  nor _74553_ (_23598_, _23597_, _23595_);
  or _74554_ (_23599_, _23598_, _16152_);
  nand _74555_ (_23600_, _23598_, _16152_);
  and _74556_ (_23601_, _23600_, _23599_);
  nor _74557_ (_23602_, _23601_, _16576_);
  and _74558_ (_23603_, _23601_, _16576_);
  or _74559_ (_23604_, _23603_, _23602_);
  nor _74560_ (_23605_, _23604_, _16812_);
  and _74561_ (_23606_, _23604_, _16812_);
  nor _74562_ (_23608_, _23606_, _23605_);
  nor _74563_ (_23609_, _23608_, _08050_);
  and _74564_ (_23610_, _23608_, _08050_);
  or _74565_ (_23611_, _23610_, _10201_);
  or _74566_ (_23612_, _23611_, _23609_);
  and _74567_ (_23613_, _23612_, _03766_);
  and _74568_ (_23614_, _23613_, _23588_);
  not _74569_ (_23615_, _08330_);
  not _74570_ (_23616_, _16134_);
  and _74571_ (_23617_, _15301_, _15034_);
  nor _74572_ (_23619_, _15301_, _15034_);
  nor _74573_ (_23620_, _23619_, _23617_);
  nor _74574_ (_23621_, _23620_, _15583_);
  and _74575_ (_23622_, _23620_, _15583_);
  nor _74576_ (_23623_, _23622_, _23621_);
  nor _74577_ (_23624_, _23623_, _15940_);
  and _74578_ (_23625_, _23623_, _15940_);
  or _74579_ (_23626_, _23625_, _23624_);
  and _74580_ (_23627_, _23626_, _23616_);
  nor _74581_ (_23628_, _23626_, _23616_);
  nor _74582_ (_23630_, _23628_, _23627_);
  and _74583_ (_23631_, _23630_, _16582_);
  nor _74584_ (_23632_, _23630_, _16582_);
  or _74585_ (_23633_, _23632_, _23631_);
  nor _74586_ (_23634_, _23633_, _16796_);
  and _74587_ (_23635_, _23633_, _16796_);
  or _74588_ (_23636_, _23635_, _23634_);
  and _74589_ (_23637_, _23636_, _23615_);
  nor _74590_ (_23638_, _23636_, _23615_);
  or _74591_ (_23639_, _23638_, _23637_);
  and _74592_ (_23640_, _23639_, _03761_);
  or _74593_ (_23641_, _23640_, _07913_);
  or _74594_ (_23642_, _23641_, _23614_);
  not _74595_ (_23643_, _07974_);
  nand _74596_ (_23644_, _15309_, _23643_);
  nand _74597_ (_23645_, _23644_, _07975_);
  nor _74598_ (_23646_, _23645_, _15599_);
  and _74599_ (_23647_, _23645_, _15599_);
  nor _74600_ (_23648_, _23647_, _23646_);
  nand _74601_ (_23649_, _23648_, _15831_);
  or _74602_ (_23651_, _23648_, _15831_);
  and _74603_ (_23652_, _23651_, _23649_);
  or _74604_ (_23653_, _23652_, _16248_);
  nand _74605_ (_23654_, _23652_, _16248_);
  and _74606_ (_23655_, _23654_, _23653_);
  nor _74607_ (_23656_, _23655_, _16476_);
  and _74608_ (_23657_, _23655_, _16476_);
  or _74609_ (_23658_, _23657_, _23656_);
  nor _74610_ (_23659_, _23658_, _16907_);
  and _74611_ (_23660_, _23658_, _16907_);
  nor _74612_ (_23662_, _23660_, _23659_);
  not _74613_ (_23663_, _23662_);
  nor _74614_ (_23664_, _23663_, _07984_);
  and _74615_ (_23665_, _23663_, _07984_);
  or _74616_ (_23666_, _23665_, _23664_);
  or _74617_ (_23667_, _23666_, _07914_);
  and _74618_ (_23668_, _23667_, _23642_);
  or _74619_ (_23669_, _23668_, _07912_);
  or _74620_ (_23670_, _05223_, _05210_);
  nor _74621_ (_23671_, _05206_, _03550_);
  and _74622_ (_23673_, _23671_, _23670_);
  nor _74623_ (_23674_, _23671_, _23670_);
  or _74624_ (_23675_, _23674_, _23673_);
  nor _74625_ (_23676_, _05261_, _05233_);
  not _74626_ (_23677_, _23676_);
  nor _74627_ (_23678_, _05227_, _05219_);
  and _74628_ (_23679_, _23678_, _23677_);
  nor _74629_ (_23680_, _23678_, _23677_);
  nor _74630_ (_23681_, _23680_, _23679_);
  nor _74631_ (_23682_, _23681_, _23675_);
  and _74632_ (_23684_, _23681_, _23675_);
  or _74633_ (_23685_, _23684_, _23682_);
  or _74634_ (_23686_, _23685_, _03248_);
  and _74635_ (_23687_, _23686_, _03710_);
  and _74636_ (_23688_, _23687_, _23669_);
  nor _74637_ (_23689_, _03625_, _03224_);
  not _74638_ (_23690_, _23689_);
  not _74639_ (_23691_, _08341_);
  and _74640_ (_23692_, _15317_, _15044_);
  nor _74641_ (_23693_, _15317_, _15044_);
  or _74642_ (_23695_, _23693_, _23692_);
  nor _74643_ (_23696_, _15951_, _15607_);
  and _74644_ (_23697_, _15951_, _15607_);
  nor _74645_ (_23698_, _23697_, _23696_);
  nor _74646_ (_23699_, _23698_, _23695_);
  and _74647_ (_23700_, _23698_, _23695_);
  nor _74648_ (_23701_, _23700_, _23699_);
  not _74649_ (_23702_, _16916_);
  nor _74650_ (_23703_, _16593_, _16257_);
  and _74651_ (_23704_, _16593_, _16257_);
  nor _74652_ (_23705_, _23704_, _23703_);
  nor _74653_ (_23706_, _23705_, _23702_);
  and _74654_ (_23707_, _23705_, _23702_);
  nor _74655_ (_23708_, _23707_, _23706_);
  nor _74656_ (_23709_, _23708_, _23701_);
  and _74657_ (_23710_, _23708_, _23701_);
  or _74658_ (_23711_, _23710_, _23709_);
  nand _74659_ (_23712_, _23711_, _23691_);
  and _74660_ (_23713_, _23711_, _03505_);
  or _74661_ (_23714_, _23713_, _08342_);
  and _74662_ (_23716_, _23714_, _23712_);
  or _74663_ (_23717_, _23716_, _23690_);
  or _74664_ (_23718_, _23717_, _23688_);
  or _74665_ (_23719_, _23689_, _23211_);
  and _74666_ (_23720_, _23719_, _23718_);
  or _74667_ (_23721_, _23720_, _10658_);
  and _74668_ (_23722_, _23433_, _06834_);
  or _74669_ (_23723_, _23722_, _06838_);
  and _74670_ (_23724_, _23723_, _23721_);
  and _74671_ (_23725_, _23433_, _06833_);
  or _74672_ (_23727_, _23725_, _04481_);
  or _74673_ (_23728_, _23727_, _23724_);
  and _74674_ (_23729_, _15324_, _15051_);
  nor _74675_ (_23730_, _15324_, _15051_);
  nor _74676_ (_23731_, _23730_, _23729_);
  not _74677_ (_23732_, _15959_);
  and _74678_ (_23733_, _23732_, _15614_);
  nor _74679_ (_23734_, _23732_, _15614_);
  nor _74680_ (_23735_, _23734_, _23733_);
  nor _74681_ (_23736_, _23735_, _23731_);
  and _74682_ (_23738_, _23735_, _23731_);
  or _74683_ (_23739_, _23738_, _23736_);
  not _74684_ (_23740_, _16600_);
  and _74685_ (_23741_, _23740_, _16265_);
  nor _74686_ (_23742_, _23740_, _16265_);
  nor _74687_ (_23743_, _23742_, _23741_);
  nand _74688_ (_23744_, _23743_, _16924_);
  or _74689_ (_23745_, _23743_, _16924_);
  and _74690_ (_23746_, _23745_, _23744_);
  or _74691_ (_23747_, _23746_, _23739_);
  nand _74692_ (_23749_, _23746_, _23739_);
  and _74693_ (_23750_, _23749_, _23747_);
  nor _74694_ (_23751_, _23750_, _08348_);
  and _74695_ (_23752_, _23750_, _08348_);
  or _74696_ (_23753_, _23752_, _07400_);
  or _74697_ (_23754_, _23753_, _23751_);
  and _74698_ (_23755_, _23754_, _03589_);
  and _74699_ (_23756_, _23755_, _23728_);
  and _74700_ (_23757_, _15329_, _15056_);
  nor _74701_ (_23758_, _15329_, _15056_);
  nor _74702_ (_23760_, _23758_, _23757_);
  and _74703_ (_23761_, _23760_, _15619_);
  nor _74704_ (_23762_, _23760_, _15619_);
  or _74705_ (_23763_, _23762_, _23761_);
  and _74706_ (_23764_, _23763_, _15965_);
  nor _74707_ (_23765_, _23763_, _15965_);
  or _74708_ (_23766_, _23765_, _23764_);
  not _74709_ (_23767_, _16606_);
  and _74710_ (_23768_, _23767_, _16270_);
  nor _74711_ (_23769_, _23767_, _16270_);
  nor _74712_ (_23770_, _23769_, _23768_);
  not _74713_ (_23771_, _16929_);
  and _74714_ (_23772_, _23771_, _08353_);
  nor _74715_ (_23773_, _23771_, _08353_);
  nor _74716_ (_23774_, _23773_, _23772_);
  or _74717_ (_23775_, _23774_, _23770_);
  nand _74718_ (_23776_, _23774_, _23770_);
  and _74719_ (_23777_, _23776_, _23775_);
  or _74720_ (_23778_, _23777_, _23766_);
  nand _74721_ (_23779_, _23777_, _23766_);
  and _74722_ (_23781_, _23779_, _03222_);
  and _74723_ (_23782_, _23781_, _23778_);
  or _74724_ (_23783_, _23782_, _07405_);
  or _74725_ (_23784_, _23783_, _23756_);
  and _74726_ (_23785_, _07463_, _16935_);
  nor _74727_ (_23786_, _07463_, _16935_);
  nor _74728_ (_23787_, _23786_, _23785_);
  nor _74729_ (_23788_, _07604_, _07547_);
  and _74730_ (_23789_, _07604_, _07547_);
  nor _74731_ (_23790_, _23789_, _23788_);
  nor _74732_ (_23792_, _23790_, _07493_);
  and _74733_ (_23793_, _23790_, _07493_);
  nor _74734_ (_23794_, _23793_, _23792_);
  nor _74735_ (_23795_, _23794_, _23787_);
  and _74736_ (_23796_, _23794_, _23787_);
  nor _74737_ (_23797_, _23796_, _23795_);
  not _74738_ (_23798_, _23797_);
  nor _74739_ (_23799_, _07674_, _07424_);
  and _74740_ (_23800_, _07674_, _07424_);
  nor _74741_ (_23801_, _23800_, _23799_);
  nor _74742_ (_23803_, _23801_, _23798_);
  and _74743_ (_23804_, _23801_, _23798_);
  nor _74744_ (_23805_, _23804_, _23803_);
  and _74745_ (_23806_, _23805_, _07760_);
  nor _74746_ (_23807_, _23805_, _07760_);
  or _74747_ (_23808_, _23807_, _07411_);
  or _74748_ (_23809_, _23808_, _23806_);
  and _74749_ (_23810_, _23809_, _03217_);
  and _74750_ (_23811_, _23810_, _23784_);
  nand _74751_ (_23812_, _23685_, _03216_);
  nor _74752_ (_23814_, _11764_, _04754_);
  and _74753_ (_23815_, _23814_, _11760_);
  and _74754_ (_23816_, _23815_, _04734_);
  and _74755_ (_23817_, _05889_, _04733_);
  and _74756_ (_23818_, _23817_, _23816_);
  nand _74757_ (_23819_, _23818_, _23812_);
  or _74758_ (_23820_, _23819_, _23811_);
  or _74759_ (_23821_, _23818_, _23211_);
  and _74760_ (_23822_, _23821_, _05886_);
  and _74761_ (_23823_, _23822_, _23820_);
  nor _74762_ (_23825_, _15339_, _14959_);
  and _74763_ (_23826_, _15339_, _14959_);
  or _74764_ (_23827_, _23826_, _23825_);
  nor _74765_ (_23828_, _15976_, _15630_);
  and _74766_ (_23829_, _15976_, _15630_);
  nor _74767_ (_23830_, _23829_, _23828_);
  nor _74768_ (_23831_, _23830_, _23827_);
  and _74769_ (_23832_, _23830_, _23827_);
  or _74770_ (_23833_, _23832_, _23831_);
  nor _74771_ (_23834_, _16445_, _16281_);
  and _74772_ (_23835_, _16445_, _16281_);
  nor _74773_ (_23836_, _23835_, _23834_);
  and _74774_ (_23837_, _23836_, _16780_);
  nor _74775_ (_23838_, _23836_, _16780_);
  nor _74776_ (_23839_, _23838_, _23837_);
  nor _74777_ (_23840_, _23839_, _23833_);
  and _74778_ (_23841_, _23839_, _23833_);
  nor _74779_ (_23842_, _23841_, _23840_);
  and _74780_ (_23843_, _23842_, _08366_);
  nor _74781_ (_23844_, _23842_, _08366_);
  or _74782_ (_23846_, _23844_, _23843_);
  and _74783_ (_23847_, _23846_, _03601_);
  or _74784_ (_23848_, _23847_, _23823_);
  and _74785_ (_23849_, _23848_, _08364_);
  nand _74786_ (_23850_, _23685_, _08363_);
  and _74787_ (_23851_, _11815_, _11348_);
  and _74788_ (_23852_, _23851_, _11820_);
  nand _74789_ (_23853_, _23852_, _23850_);
  or _74790_ (_23854_, _23853_, _23849_);
  or _74791_ (_23855_, _23852_, _23211_);
  and _74792_ (_23857_, _23855_, _11343_);
  and _74793_ (_23858_, _23857_, _23854_);
  nor _74794_ (_23859_, _15799_, _08676_);
  and _74795_ (_23860_, _15799_, _08676_);
  nor _74796_ (_23861_, _23860_, _23859_);
  and _74797_ (_23862_, _15072_, _08680_);
  nor _74798_ (_23863_, _23862_, _15550_);
  nor _74799_ (_23864_, _23863_, _23861_);
  and _74800_ (_23865_, _23863_, _23861_);
  nor _74801_ (_23866_, _23865_, _23864_);
  nor _74802_ (_23868_, _16453_, _08669_);
  and _74803_ (_23869_, _16453_, _08669_);
  nor _74804_ (_23870_, _23869_, _23868_);
  nor _74805_ (_23871_, _23870_, _23866_);
  and _74806_ (_23872_, _23870_, _23866_);
  nor _74807_ (_23873_, _23872_, _23871_);
  not _74808_ (_23874_, _23873_);
  and _74809_ (_23875_, _08664_, _08376_);
  nor _74810_ (_23876_, _08664_, _08376_);
  nor _74811_ (_23877_, _23876_, _23875_);
  nor _74812_ (_23879_, _23877_, _23874_);
  and _74813_ (_23880_, _23877_, _23874_);
  or _74814_ (_23881_, _23880_, _23879_);
  and _74815_ (_23882_, _23881_, _11344_);
  or _74816_ (_23883_, _23882_, _08392_);
  or _74817_ (_23884_, _23883_, _23858_);
  nor _74818_ (_23885_, _15921_, _08640_);
  and _74819_ (_23886_, _15921_, _08640_);
  nor _74820_ (_23887_, _23886_, _23885_);
  and _74821_ (_23888_, _15083_, _08644_);
  nor _74822_ (_23890_, _23888_, _15568_);
  nor _74823_ (_23891_, _23890_, _23887_);
  and _74824_ (_23892_, _23890_, _23887_);
  nor _74825_ (_23893_, _23892_, _23891_);
  nor _74826_ (_23894_, _08630_, _08634_);
  and _74827_ (_23895_, _08630_, _08634_);
  nor _74828_ (_23896_, _23895_, _23894_);
  nor _74829_ (_23897_, _23896_, _23893_);
  and _74830_ (_23898_, _23896_, _23893_);
  nor _74831_ (_23899_, _23898_, _23897_);
  nor _74832_ (_23900_, _23899_, _08627_);
  and _74833_ (_23901_, _23899_, _08627_);
  or _74834_ (_23902_, _23901_, _23900_);
  and _74835_ (_23903_, _23902_, _08400_);
  nor _74836_ (_23904_, _23902_, _08400_);
  or _74837_ (_23905_, _23904_, _23903_);
  or _74838_ (_23906_, _23905_, _08393_);
  and _74839_ (_23907_, _23906_, _03779_);
  and _74840_ (_23908_, _23907_, _23884_);
  nor _74841_ (_23909_, _12739_, _12539_);
  and _74842_ (_23911_, _12739_, _12539_);
  nor _74843_ (_23912_, _23911_, _23909_);
  nor _74844_ (_23913_, _12333_, _12128_);
  and _74845_ (_23914_, _12333_, _12128_);
  nor _74846_ (_23915_, _23914_, _23913_);
  not _74847_ (_23916_, _23915_);
  and _74848_ (_23917_, _23916_, _23912_);
  nor _74849_ (_23918_, _23916_, _23912_);
  nor _74850_ (_23919_, _23918_, _23917_);
  or _74851_ (_23920_, _23919_, _12817_);
  nand _74852_ (_23922_, _23919_, _12817_);
  and _74853_ (_23923_, _23922_, _23920_);
  or _74854_ (_23924_, _23923_, _13147_);
  nand _74855_ (_23925_, _23923_, _13147_);
  and _74856_ (_23926_, _23925_, _23924_);
  or _74857_ (_23927_, _23926_, _13353_);
  nand _74858_ (_23928_, _23926_, _13353_);
  and _74859_ (_23929_, _23928_, _23927_);
  nor _74860_ (_23930_, _23929_, _06378_);
  and _74861_ (_23931_, _23929_, _06378_);
  or _74862_ (_23933_, _23931_, _23930_);
  and _74863_ (_23934_, _23933_, _03778_);
  or _74864_ (_23935_, _23934_, _07904_);
  or _74865_ (_23936_, _23935_, _23908_);
  and _74866_ (_23937_, _16734_, _08737_);
  and _74867_ (_23938_, _10026_, _08738_);
  nor _74868_ (_23939_, _23938_, _23937_);
  not _74869_ (_23940_, _10058_);
  nor _74870_ (_23941_, _08753_, _23940_);
  and _74871_ (_23942_, _08753_, _23940_);
  nor _74872_ (_23944_, _23942_, _23941_);
  and _74873_ (_23945_, _10030_, _08748_);
  nor _74874_ (_23946_, _23945_, _10031_);
  and _74875_ (_23947_, _23946_, _23944_);
  nor _74876_ (_23948_, _23946_, _23944_);
  nor _74877_ (_23949_, _23948_, _23947_);
  nor _74878_ (_23950_, _23949_, _08743_);
  and _74879_ (_23951_, _23949_, _08743_);
  or _74880_ (_23952_, _23951_, _23950_);
  nor _74881_ (_23953_, _23952_, _23939_);
  and _74882_ (_23955_, _23952_, _23939_);
  nor _74883_ (_23956_, _23955_, _23953_);
  nand _74884_ (_23957_, _23956_, _08407_);
  or _74885_ (_23958_, _23956_, _08407_);
  and _74886_ (_23959_, _23958_, _23957_);
  or _74887_ (_23960_, _23959_, _07905_);
  and _74888_ (_23961_, _23960_, _07766_);
  and _74889_ (_23962_, _23961_, _23936_);
  and _74890_ (_23963_, _15209_, _14965_);
  nor _74891_ (_23964_, _15209_, _14965_);
  nor _74892_ (_23966_, _23964_, _23963_);
  and _74893_ (_23967_, _23966_, _15474_);
  nor _74894_ (_23968_, _23966_, _15474_);
  or _74895_ (_23969_, _23968_, _23967_);
  nand _74896_ (_23970_, _23969_, _15813_);
  or _74897_ (_23971_, _23969_, _15813_);
  and _74898_ (_23972_, _23971_, _23970_);
  nor _74899_ (_23973_, _16784_, _16450_);
  and _74900_ (_23974_, _16784_, _16450_);
  nor _74901_ (_23975_, _23974_, _23973_);
  not _74902_ (_23977_, _16124_);
  and _74903_ (_23978_, _23977_, _07902_);
  nor _74904_ (_23979_, _23977_, _07902_);
  nor _74905_ (_23980_, _23979_, _23978_);
  nor _74906_ (_23981_, _23980_, _23975_);
  and _74907_ (_23982_, _23980_, _23975_);
  nor _74908_ (_23983_, _23982_, _23981_);
  nand _74909_ (_23984_, _23983_, _23972_);
  or _74910_ (_23985_, _23983_, _23972_);
  and _74911_ (_23986_, _23985_, _03600_);
  and _74912_ (_23988_, _23986_, _23984_);
  or _74913_ (_23989_, _23988_, _23962_);
  and _74914_ (_23990_, _23989_, _07778_);
  nor _74915_ (_23991_, _11841_, _03182_);
  nand _74916_ (_23992_, _23211_, _03780_);
  or _74917_ (_23993_, _23992_, _05254_);
  nand _74918_ (_23994_, _23993_, _23991_);
  or _74919_ (_23995_, _23994_, _23990_);
  or _74920_ (_23996_, _23991_, _23211_);
  and _74921_ (_23997_, _23996_, _08414_);
  and _74922_ (_23999_, _23997_, _08416_);
  and _74923_ (_24000_, _23999_, _23995_);
  or _74924_ (_24001_, _08681_, _08678_);
  nand _74925_ (_24002_, _08681_, _08678_);
  and _74926_ (_24003_, _24002_, _24001_);
  nor _74927_ (_24004_, _08672_, _08674_);
  and _74928_ (_24005_, _08672_, _08674_);
  nor _74929_ (_24006_, _24005_, _24004_);
  and _74930_ (_24007_, _24006_, _24003_);
  nor _74931_ (_24008_, _24006_, _24003_);
  nor _74932_ (_24010_, _24008_, _24007_);
  and _74933_ (_24011_, _08662_, _08375_);
  or _74934_ (_24012_, _24011_, _10329_);
  nor _74935_ (_24013_, _08665_, _08667_);
  and _74936_ (_24014_, _08665_, _08667_);
  nor _74937_ (_24015_, _24014_, _24013_);
  not _74938_ (_24016_, _24015_);
  and _74939_ (_24017_, _24016_, _24012_);
  nor _74940_ (_24018_, _24016_, _24012_);
  nor _74941_ (_24019_, _24018_, _24017_);
  nor _74942_ (_24021_, _24019_, _24010_);
  and _74943_ (_24022_, _24019_, _24010_);
  or _74944_ (_24023_, _24022_, _24021_);
  and _74945_ (_24024_, _24023_, _08421_);
  or _74946_ (_24025_, _24024_, _08420_);
  or _74947_ (_24026_, _24025_, _24000_);
  not _74948_ (_24027_, _08638_);
  or _74949_ (_24028_, _08645_, _08642_);
  nand _74950_ (_24029_, _08645_, _08642_);
  and _74951_ (_24030_, _24029_, _24028_);
  nand _74952_ (_24032_, _24030_, _24027_);
  or _74953_ (_24033_, _24030_, _24027_);
  and _74954_ (_24034_, _24033_, _24032_);
  nor _74955_ (_24035_, _24034_, _08635_);
  and _74956_ (_24036_, _24034_, _08635_);
  or _74957_ (_24037_, _24036_, _24035_);
  not _74958_ (_24038_, _08628_);
  nor _74959_ (_24039_, _08632_, _08625_);
  and _74960_ (_24040_, _08632_, _08625_);
  nor _74961_ (_24041_, _24040_, _24039_);
  nor _74962_ (_24043_, _24041_, _24038_);
  and _74963_ (_24044_, _24041_, _24038_);
  nor _74964_ (_24045_, _24044_, _24043_);
  nor _74965_ (_24046_, _24045_, _24037_);
  and _74966_ (_24047_, _24045_, _24037_);
  nor _74967_ (_24048_, _24047_, _24046_);
  and _74968_ (_24049_, _24048_, _08399_);
  nor _74969_ (_24050_, _24048_, _08399_);
  or _74970_ (_24051_, _24050_, _24049_);
  or _74971_ (_24052_, _24051_, _08425_);
  and _74972_ (_24054_, _24052_, _03789_);
  and _74973_ (_24055_, _24054_, _24026_);
  nor _74974_ (_24056_, _12331_, _12005_);
  and _74975_ (_24057_, _12331_, _12005_);
  nor _74976_ (_24058_, _24057_, _24056_);
  not _74977_ (_24059_, _24058_);
  not _74978_ (_24060_, _12737_);
  and _74979_ (_24061_, _24060_, _12537_);
  nor _74980_ (_24062_, _24060_, _12537_);
  nor _74981_ (_24063_, _24062_, _24061_);
  nor _74982_ (_24065_, _24063_, _24059_);
  and _74983_ (_24066_, _24063_, _24059_);
  nor _74984_ (_24067_, _24066_, _24065_);
  not _74985_ (_24068_, _13351_);
  nor _74986_ (_24069_, _13145_, _12815_);
  and _74987_ (_24070_, _13145_, _12815_);
  nor _74988_ (_24071_, _24070_, _24069_);
  nor _74989_ (_24072_, _24071_, _24068_);
  and _74990_ (_24073_, _24071_, _24068_);
  nor _74991_ (_24074_, _24073_, _24072_);
  not _74992_ (_24076_, _24074_);
  nor _74993_ (_24077_, _24076_, _24067_);
  and _74994_ (_24078_, _24076_, _24067_);
  nor _74995_ (_24079_, _24078_, _24077_);
  or _74996_ (_24080_, _24079_, _06376_);
  nand _74997_ (_24081_, _24079_, _06376_);
  and _74998_ (_24082_, _24081_, _03788_);
  and _74999_ (_24083_, _24082_, _24080_);
  or _75000_ (_24084_, _24083_, _08429_);
  or _75001_ (_24085_, _24084_, _24055_);
  not _75002_ (_24087_, _08741_);
  or _75003_ (_24088_, _08750_, _08751_);
  nand _75004_ (_24089_, _08750_, _08751_);
  and _75005_ (_24090_, _24089_, _24088_);
  not _75006_ (_24091_, _08744_);
  and _75007_ (_24092_, _24091_, _08746_);
  nor _75008_ (_24093_, _24091_, _08746_);
  nor _75009_ (_24094_, _24093_, _24092_);
  not _75010_ (_24095_, _24094_);
  and _75011_ (_24096_, _24095_, _24090_);
  nor _75012_ (_24098_, _24095_, _24090_);
  nor _75013_ (_24099_, _24098_, _24096_);
  nand _75014_ (_24100_, _24099_, _24087_);
  or _75015_ (_24101_, _24099_, _24087_);
  and _75016_ (_24102_, _24101_, _24100_);
  or _75017_ (_24103_, _24102_, _08739_);
  nand _75018_ (_24104_, _24102_, _08739_);
  and _75019_ (_24105_, _24104_, _24103_);
  or _75020_ (_24106_, _24105_, _08735_);
  nand _75021_ (_24107_, _24105_, _08735_);
  and _75022_ (_24109_, _24107_, _24106_);
  nor _75023_ (_24110_, _24109_, _08405_);
  and _75024_ (_24111_, _24109_, _08405_);
  or _75025_ (_24112_, _24111_, _24110_);
  or _75026_ (_24113_, _24112_, _08435_);
  and _75027_ (_24114_, _24113_, _07777_);
  and _75028_ (_24115_, _24114_, _24085_);
  and _75029_ (_24116_, _11338_, _10753_);
  nor _75030_ (_24117_, _15687_, _14960_);
  and _75031_ (_24118_, _15687_, _14960_);
  nor _75032_ (_24120_, _24118_, _24117_);
  nor _75033_ (_24121_, _16781_, _16333_);
  and _75034_ (_24122_, _16781_, _16333_);
  nor _75035_ (_24123_, _24122_, _24121_);
  and _75036_ (_24124_, _24123_, _24120_);
  nor _75037_ (_24125_, _24123_, _24120_);
  nor _75038_ (_24126_, _24125_, _24124_);
  nor _75039_ (_24127_, _16447_, _16017_);
  and _75040_ (_24128_, _16447_, _16017_);
  nor _75041_ (_24129_, _24128_, _24127_);
  nor _75042_ (_24131_, _15206_, _08439_);
  and _75043_ (_24132_, _15206_, _08439_);
  nor _75044_ (_24133_, _24132_, _24131_);
  and _75045_ (_24134_, _24133_, _24129_);
  nor _75046_ (_24135_, _24133_, _24129_);
  nor _75047_ (_24136_, _24135_, _24134_);
  not _75048_ (_24137_, _24136_);
  nand _75049_ (_24138_, _24137_, _24126_);
  or _75050_ (_24139_, _24137_, _24126_);
  and _75051_ (_24140_, _24139_, _03622_);
  nand _75052_ (_24142_, _24140_, _24138_);
  nand _75053_ (_24143_, _24142_, _24116_);
  or _75054_ (_24144_, _24143_, _24115_);
  or _75055_ (_24145_, _23211_, _24116_);
  and _75056_ (_24146_, _24145_, _08447_);
  and _75057_ (_24147_, _24146_, _24144_);
  nor _75058_ (_24148_, _15071_, _08679_);
  and _75059_ (_24149_, _15071_, _08679_);
  nor _75060_ (_24150_, _24149_, _24148_);
  and _75061_ (_24151_, _24150_, _08675_);
  nor _75062_ (_24153_, _24150_, _08675_);
  or _75063_ (_24154_, _24153_, _24151_);
  nand _75064_ (_24155_, _24154_, _08673_);
  or _75065_ (_24156_, _24154_, _08673_);
  and _75066_ (_24157_, _24156_, _24155_);
  not _75067_ (_24158_, _08666_);
  nor _75068_ (_24159_, _08668_, _08663_);
  and _75069_ (_24160_, _08668_, _08663_);
  nor _75070_ (_24161_, _24160_, _24159_);
  nor _75071_ (_24162_, _24161_, _24158_);
  and _75072_ (_24164_, _24161_, _24158_);
  nor _75073_ (_24165_, _24164_, _24162_);
  and _75074_ (_24166_, _24165_, _24157_);
  nor _75075_ (_24167_, _24165_, _24157_);
  or _75076_ (_24168_, _24167_, _24166_);
  and _75077_ (_24169_, _24168_, _08374_);
  nor _75078_ (_24170_, _24168_, _08374_);
  or _75079_ (_24171_, _24170_, _24169_);
  and _75080_ (_24172_, _24171_, _08446_);
  or _75081_ (_24173_, _24172_, _08450_);
  or _75082_ (_24175_, _24173_, _24147_);
  not _75083_ (_24176_, _08398_);
  nor _75084_ (_24177_, _15082_, _08643_);
  and _75085_ (_24178_, _15082_, _08643_);
  nor _75086_ (_24179_, _24178_, _24177_);
  and _75087_ (_24180_, _24179_, _08639_);
  nor _75088_ (_24181_, _24179_, _08639_);
  or _75089_ (_24182_, _24181_, _24180_);
  nand _75090_ (_24183_, _24182_, _08637_);
  or _75091_ (_24184_, _24182_, _08637_);
  and _75092_ (_24187_, _24184_, _24183_);
  nor _75093_ (_24188_, _08633_, _08626_);
  and _75094_ (_24189_, _08633_, _08626_);
  nor _75095_ (_24190_, _24189_, _24188_);
  and _75096_ (_24191_, _24190_, _08629_);
  nor _75097_ (_24192_, _24190_, _08629_);
  nor _75098_ (_24193_, _24192_, _24191_);
  and _75099_ (_24194_, _24193_, _24187_);
  nor _75100_ (_24195_, _24193_, _24187_);
  or _75101_ (_24196_, _24195_, _24194_);
  nor _75102_ (_24199_, _24196_, _24176_);
  and _75103_ (_24200_, _24196_, _24176_);
  nor _75104_ (_24201_, _24200_, _24199_);
  nand _75105_ (_24202_, _24201_, _08450_);
  and _75106_ (_24203_, _24202_, _03784_);
  and _75107_ (_24204_, _24203_, _24175_);
  or _75108_ (_24205_, _24204_, _23261_);
  and _75109_ (_24206_, _24205_, _08461_);
  nor _75110_ (_24207_, _08752_, _10057_);
  and _75111_ (_24208_, _08752_, _10057_);
  nor _75112_ (_24211_, _24208_, _24207_);
  not _75113_ (_24212_, _24211_);
  not _75114_ (_24213_, _08745_);
  and _75115_ (_24214_, _24213_, _08747_);
  nor _75116_ (_24215_, _24213_, _08747_);
  nor _75117_ (_24216_, _24215_, _24214_);
  nor _75118_ (_24217_, _24216_, _24212_);
  and _75119_ (_24218_, _24216_, _24212_);
  nor _75120_ (_24219_, _24218_, _24217_);
  and _75121_ (_24220_, _24219_, _08742_);
  nor _75122_ (_24223_, _24219_, _08742_);
  or _75123_ (_24224_, _24223_, _24220_);
  and _75124_ (_24225_, _24224_, _08740_);
  nor _75125_ (_24226_, _24224_, _08740_);
  or _75126_ (_24227_, _24226_, _24225_);
  and _75127_ (_24228_, _24227_, _08736_);
  nor _75128_ (_24229_, _24227_, _08736_);
  or _75129_ (_24230_, _24229_, _24228_);
  and _75130_ (_24231_, _24230_, _08406_);
  nor _75131_ (_24232_, _24230_, _08406_);
  or _75132_ (_24235_, _24232_, _24231_);
  and _75133_ (_24236_, _24235_, _08458_);
  or _75134_ (_24237_, _24236_, _24206_);
  and _75135_ (_24238_, _24237_, _07795_);
  and _75136_ (_24239_, _11881_, _11877_);
  nor _75137_ (_24240_, _15401_, _15144_);
  and _75138_ (_24241_, _15401_, _15144_);
  or _75139_ (_24242_, _24241_, _24240_);
  nor _75140_ (_24243_, _16037_, _15710_);
  and _75141_ (_24244_, _16037_, _15710_);
  nor _75142_ (_24247_, _24244_, _24243_);
  nor _75143_ (_24248_, _24247_, _24242_);
  and _75144_ (_24249_, _24247_, _24242_);
  nor _75145_ (_24250_, _24249_, _24248_);
  not _75146_ (_24251_, _24250_);
  nor _75147_ (_24252_, _17004_, _16442_);
  and _75148_ (_24253_, _17004_, _16442_);
  nor _75149_ (_24254_, _24253_, _24252_);
  not _75150_ (_24255_, _16352_);
  and _75151_ (_24256_, _24255_, _08470_);
  nor _75152_ (_24259_, _24255_, _08470_);
  nor _75153_ (_24260_, _24259_, _24256_);
  nor _75154_ (_24261_, _24260_, _24254_);
  and _75155_ (_24262_, _24260_, _24254_);
  nor _75156_ (_24263_, _24262_, _24261_);
  nand _75157_ (_24264_, _24263_, _24251_);
  or _75158_ (_24265_, _24263_, _24251_);
  and _75159_ (_24266_, _24265_, _03624_);
  nand _75160_ (_24267_, _24266_, _24264_);
  nand _75161_ (_24268_, _24267_, _24239_);
  or _75162_ (_24270_, _24268_, _24238_);
  or _75163_ (_24271_, _23211_, _24239_);
  and _75164_ (_24272_, _24271_, _07898_);
  and _75165_ (_24273_, _24272_, _24270_);
  not _75166_ (_24274_, _15805_);
  nor _75167_ (_24275_, _15406_, _08170_);
  and _75168_ (_24276_, _15406_, _08170_);
  or _75169_ (_24277_, _24276_, _24275_);
  nor _75170_ (_24278_, _24277_, _15716_);
  and _75171_ (_24279_, _24277_, _15716_);
  nor _75172_ (_24281_, _24279_, _24278_);
  and _75173_ (_24282_, _24281_, _24274_);
  nor _75174_ (_24283_, _24281_, _24274_);
  nor _75175_ (_24284_, _24283_, _24282_);
  nor _75176_ (_24285_, _24284_, _16357_);
  and _75177_ (_24286_, _24284_, _16357_);
  or _75178_ (_24287_, _24286_, _24285_);
  and _75179_ (_24288_, _24287_, _16684_);
  nor _75180_ (_24289_, _24287_, _16684_);
  nor _75181_ (_24290_, _24289_, _24288_);
  nor _75182_ (_24292_, _24290_, _17010_);
  and _75183_ (_24293_, _24290_, _17010_);
  or _75184_ (_24294_, _24293_, _24292_);
  nor _75185_ (_24295_, _24294_, _07890_);
  and _75186_ (_24296_, _24294_, _07890_);
  or _75187_ (_24297_, _24296_, _24295_);
  and _75188_ (_24298_, _24297_, _08468_);
  or _75189_ (_24299_, _24298_, _08475_);
  or _75190_ (_24300_, _24299_, _24273_);
  not _75191_ (_24301_, _16690_);
  not _75192_ (_24303_, _16045_);
  nor _75193_ (_24304_, _15411_, _15029_);
  and _75194_ (_24305_, _15411_, _15029_);
  or _75195_ (_24306_, _24305_, _24304_);
  nor _75196_ (_24307_, _24306_, _15721_);
  and _75197_ (_24308_, _24306_, _15721_);
  nor _75198_ (_24309_, _24308_, _24307_);
  and _75199_ (_24310_, _24309_, _24303_);
  nor _75200_ (_24311_, _24309_, _24303_);
  nor _75201_ (_24312_, _24311_, _24310_);
  nor _75202_ (_24314_, _24312_, _16363_);
  and _75203_ (_24315_, _24312_, _16363_);
  or _75204_ (_24316_, _24315_, _24314_);
  nor _75205_ (_24317_, _24316_, _24301_);
  and _75206_ (_24318_, _24316_, _24301_);
  nor _75207_ (_24319_, _24318_, _24317_);
  and _75208_ (_24320_, _24319_, _17015_);
  nor _75209_ (_24321_, _24319_, _17015_);
  or _75210_ (_24322_, _24321_, _24320_);
  not _75211_ (_24323_, _24322_);
  nor _75212_ (_24325_, _24323_, _08502_);
  and _75213_ (_24326_, _24323_, _08502_);
  or _75214_ (_24327_, _24326_, _24325_);
  or _75215_ (_24328_, _24327_, _08477_);
  and _75216_ (_24329_, _24328_, _03777_);
  and _75217_ (_24330_, _24329_, _24300_);
  nor _75218_ (_24331_, _15416_, _15034_);
  and _75219_ (_24332_, _15416_, _15034_);
  or _75220_ (_24333_, _24332_, _24331_);
  nor _75221_ (_24334_, _24333_, _15727_);
  and _75222_ (_24336_, _24333_, _15727_);
  nor _75223_ (_24337_, _24336_, _24334_);
  nor _75224_ (_24338_, _24337_, _16050_);
  and _75225_ (_24339_, _24337_, _16050_);
  or _75226_ (_24340_, _24339_, _24338_);
  nor _75227_ (_24341_, _24340_, _16368_);
  and _75228_ (_24342_, _24340_, _16368_);
  or _75229_ (_24343_, _24342_, _24341_);
  nor _75230_ (_24344_, _24343_, _16695_);
  and _75231_ (_24345_, _24343_, _16695_);
  or _75232_ (_24347_, _24345_, _24344_);
  and _75233_ (_24348_, _24347_, _17021_);
  nor _75234_ (_24349_, _24347_, _17021_);
  or _75235_ (_24350_, _24349_, _24348_);
  or _75236_ (_24351_, _24350_, _08583_);
  nand _75237_ (_24352_, _24350_, _08583_);
  and _75238_ (_24353_, _24352_, _03776_);
  and _75239_ (_24354_, _24353_, _24351_);
  or _75240_ (_24355_, _24354_, _08506_);
  or _75241_ (_24356_, _24355_, _24330_);
  not _75242_ (_24358_, _08613_);
  and _75243_ (_24359_, _15421_, _07974_);
  and _75244_ (_24360_, _23643_, _07972_);
  nor _75245_ (_24361_, _24360_, _24359_);
  nor _75246_ (_24362_, _24361_, _15732_);
  and _75247_ (_24363_, _24361_, _15732_);
  nor _75248_ (_24364_, _24363_, _24362_);
  or _75249_ (_24365_, _24364_, _16056_);
  nand _75250_ (_24366_, _24364_, _16056_);
  and _75251_ (_24367_, _24366_, _24365_);
  nor _75252_ (_24369_, _24367_, _16374_);
  and _75253_ (_24370_, _24367_, _16374_);
  nor _75254_ (_24371_, _24370_, _24369_);
  nor _75255_ (_24372_, _24371_, _16701_);
  and _75256_ (_24373_, _24371_, _16701_);
  or _75257_ (_24374_, _24373_, _24372_);
  and _75258_ (_24375_, _24374_, _17026_);
  nor _75259_ (_24376_, _24374_, _17026_);
  nor _75260_ (_24377_, _24376_, _24375_);
  nor _75261_ (_24378_, _24377_, _24358_);
  and _75262_ (_24380_, _24377_, _24358_);
  or _75263_ (_24381_, _24380_, _24378_);
  or _75264_ (_24382_, _24381_, _08589_);
  and _75265_ (_24383_, _24382_, _08588_);
  and _75266_ (_24384_, _24383_, _24356_);
  or _75267_ (_24385_, _24384_, _23235_);
  and _75268_ (_24386_, _10774_, _11903_);
  and _75269_ (_24387_, _24386_, _24385_);
  not _75270_ (_24388_, _24386_);
  nand _75271_ (_24389_, _24388_, _23211_);
  nand _75272_ (_24391_, _24389_, _16706_);
  or _75273_ (_24392_, _24391_, _24387_);
  not _75274_ (_24393_, _15071_);
  and _75275_ (_24394_, _24393_, _08680_);
  nor _75276_ (_24395_, _24393_, _08680_);
  nor _75277_ (_24396_, _24395_, _24394_);
  and _75278_ (_24397_, _24396_, _15741_);
  nor _75279_ (_24398_, _24396_, _15741_);
  nor _75280_ (_24399_, _24398_, _24397_);
  and _75281_ (_24400_, _24399_, _15802_);
  nor _75282_ (_24402_, _24399_, _15802_);
  or _75283_ (_24403_, _24402_, _24400_);
  and _75284_ (_24404_, _24403_, _16383_);
  nor _75285_ (_24405_, _24403_, _16383_);
  nor _75286_ (_24406_, _24405_, _24404_);
  nor _75287_ (_24407_, _24406_, _16715_);
  and _75288_ (_24408_, _24406_, _16715_);
  nor _75289_ (_24409_, _24408_, _24407_);
  and _75290_ (_24410_, _24409_, _17035_);
  nor _75291_ (_24411_, _24409_, _17035_);
  or _75292_ (_24413_, _24411_, _24410_);
  nor _75293_ (_24414_, _24413_, _08696_);
  and _75294_ (_24415_, _24413_, _08696_);
  or _75295_ (_24416_, _24415_, _24414_);
  or _75296_ (_24417_, _24416_, _16706_);
  and _75297_ (_24418_, _24417_, _16712_);
  and _75298_ (_24419_, _24418_, _24392_);
  and _75299_ (_24420_, _24416_, _16710_);
  or _75300_ (_24421_, _24420_, _08620_);
  or _75301_ (_24422_, _24421_, _24419_);
  not _75302_ (_24424_, _08660_);
  and _75303_ (_24425_, _15082_, _08644_);
  nor _75304_ (_24426_, _15082_, _08644_);
  or _75305_ (_24427_, _24426_, _24425_);
  and _75306_ (_24428_, _24427_, _15747_);
  nor _75307_ (_24429_, _24427_, _15747_);
  nor _75308_ (_24430_, _24429_, _24428_);
  nor _75309_ (_24431_, _24430_, _16068_);
  and _75310_ (_24432_, _24430_, _16068_);
  or _75311_ (_24433_, _24432_, _24431_);
  nor _75312_ (_24435_, _24433_, _16388_);
  and _75313_ (_24436_, _24433_, _16388_);
  or _75314_ (_24437_, _24436_, _24435_);
  and _75315_ (_24438_, _24437_, _16724_);
  nor _75316_ (_24439_, _24437_, _16724_);
  nor _75317_ (_24440_, _24439_, _24438_);
  nor _75318_ (_24441_, _24440_, _17041_);
  and _75319_ (_24442_, _24440_, _17041_);
  or _75320_ (_24443_, _24442_, _24441_);
  nor _75321_ (_24444_, _24443_, _24424_);
  and _75322_ (_24446_, _24443_, _24424_);
  or _75323_ (_24447_, _24446_, _24444_);
  or _75324_ (_24448_, _24447_, _08624_);
  and _75325_ (_24449_, _24448_, _03518_);
  and _75326_ (_24450_, _24449_, _24422_);
  nor _75327_ (_24451_, _15436_, _08318_);
  and _75328_ (_24452_, _15436_, _08318_);
  or _75329_ (_24453_, _24452_, _24451_);
  nor _75330_ (_24454_, _24453_, _15752_);
  and _75331_ (_24455_, _24453_, _15752_);
  nor _75332_ (_24457_, _24455_, _24454_);
  and _75333_ (_24458_, _24457_, _16075_);
  nor _75334_ (_24459_, _24457_, _16075_);
  nor _75335_ (_24460_, _24459_, _24458_);
  and _75336_ (_24461_, _24460_, _16394_);
  nor _75337_ (_24462_, _24460_, _16394_);
  nor _75338_ (_24463_, _24462_, _24461_);
  nor _75339_ (_24464_, _24463_, _16729_);
  and _75340_ (_24465_, _24463_, _16729_);
  or _75341_ (_24466_, _24465_, _24464_);
  nor _75342_ (_24468_, _24466_, _17046_);
  and _75343_ (_24469_, _24466_, _17046_);
  or _75344_ (_24470_, _24469_, _24468_);
  or _75345_ (_24471_, _24470_, _08728_);
  nand _75346_ (_24472_, _24470_, _08728_);
  and _75347_ (_24473_, _24472_, _03517_);
  and _75348_ (_24474_, _24473_, _24471_);
  or _75349_ (_24475_, _24474_, _24450_);
  and _75350_ (_24476_, _24475_, _08734_);
  and _75351_ (_24477_, _15441_, _23940_);
  nor _75352_ (_24479_, _24477_, _23941_);
  and _75353_ (_24480_, _24479_, _15758_);
  nor _75354_ (_24481_, _24479_, _15758_);
  nor _75355_ (_24482_, _24481_, _24480_);
  nor _75356_ (_24483_, _24482_, _16081_);
  and _75357_ (_24484_, _24482_, _16081_);
  nor _75358_ (_24485_, _24484_, _24483_);
  nor _75359_ (_24486_, _24485_, _16399_);
  and _75360_ (_24487_, _24485_, _16399_);
  or _75361_ (_24488_, _24487_, _24486_);
  nor _75362_ (_24490_, _24488_, _16737_);
  and _75363_ (_24491_, _24488_, _16737_);
  or _75364_ (_24492_, _24491_, _24490_);
  nor _75365_ (_24493_, _24492_, _17052_);
  and _75366_ (_24494_, _24492_, _17052_);
  or _75367_ (_24495_, _24494_, _24493_);
  nor _75368_ (_24496_, _24495_, _08768_);
  and _75369_ (_24497_, _24495_, _08768_);
  or _75370_ (_24498_, _24497_, _24496_);
  nand _75371_ (_24499_, _24498_, _08701_);
  nand _75372_ (_24501_, _24499_, _23218_);
  or _75373_ (_24502_, _24501_, _24476_);
  and _75374_ (_24503_, _24502_, _23219_);
  or _75375_ (_24504_, _24503_, _03815_);
  or _75376_ (_24505_, _23352_, _04246_);
  and _75377_ (_24506_, _24505_, _08776_);
  and _75378_ (_24507_, _24506_, _24504_);
  not _75379_ (_24508_, _08781_);
  and _75380_ (_24509_, _15503_, _24508_);
  and _75381_ (_24510_, _24509_, \oc8051_golden_model_1.ACC [3]);
  nor _75382_ (_24512_, _24509_, \oc8051_golden_model_1.ACC [3]);
  nor _75383_ (_24513_, _24512_, _24510_);
  and _75384_ (_24514_, _24513_, _16412_);
  nor _75385_ (_24515_, _24513_, _16412_);
  nor _75386_ (_24516_, _24515_, _24514_);
  and _75387_ (_24517_, _16748_, _07433_);
  nor _75388_ (_24518_, _16748_, _07433_);
  nor _75389_ (_24519_, _24518_, _24517_);
  nor _75390_ (_24520_, _24519_, _24516_);
  and _75391_ (_24521_, _24519_, _24516_);
  or _75392_ (_24523_, _24521_, _24520_);
  or _75393_ (_24524_, _24523_, _08788_);
  nand _75394_ (_24525_, _24523_, _08788_);
  and _75395_ (_24526_, _24525_, _24524_);
  and _75396_ (_24527_, _24526_, _08775_);
  or _75397_ (_24528_, _24527_, _24507_);
  and _75398_ (_24529_, _24528_, _10359_);
  and _75399_ (_24530_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor _75400_ (_24531_, _24530_, _08110_);
  nand _75401_ (_24532_, _24531_, _23230_);
  or _75402_ (_24534_, _24531_, _23230_);
  and _75403_ (_24535_, _24534_, _24532_);
  nand _75404_ (_24536_, _24535_, _08780_);
  nand _75405_ (_24537_, _24536_, _04540_);
  or _75406_ (_24538_, _24537_, _24529_);
  or _75407_ (_24539_, _23211_, _04540_);
  and _75408_ (_24540_, _24539_, _03823_);
  and _75409_ (_24541_, _24540_, _24538_);
  or _75410_ (_24542_, _24541_, _23194_);
  and _75411_ (_24543_, _24542_, _11955_);
  and _75412_ (_24545_, _23211_, _11956_);
  or _75413_ (_24546_, _24545_, _04552_);
  or _75414_ (_24547_, _24546_, _24543_);
  or _75415_ (_24548_, _23211_, _06785_);
  and _75416_ (_24549_, _24548_, _03514_);
  and _75417_ (_24550_, _24549_, _24547_);
  or _75418_ (_24551_, _24550_, _23170_);
  and _75419_ (_24552_, _24551_, _08799_);
  nor _75420_ (_24553_, _11975_, _03196_);
  nor _75421_ (_24554_, _08805_, _03631_);
  and _75422_ (_24556_, _24554_, _24553_);
  not _75423_ (_24557_, _08806_);
  and _75424_ (_24558_, _15503_, _24557_);
  and _75425_ (_24559_, _24558_, _07578_);
  nor _75426_ (_24560_, _24558_, _07578_);
  nor _75427_ (_24561_, _24560_, _24559_);
  nor _75428_ (_24562_, _17080_, _16430_);
  and _75429_ (_24563_, _17080_, _16430_);
  or _75430_ (_24564_, _24563_, _24562_);
  or _75431_ (_24565_, _24564_, _24561_);
  nand _75432_ (_24567_, _24564_, _24561_);
  and _75433_ (_24568_, _24567_, _24565_);
  nor _75434_ (_24569_, _16767_, _08813_);
  and _75435_ (_24570_, _16767_, _08813_);
  nor _75436_ (_24571_, _24570_, _24569_);
  not _75437_ (_24572_, _24571_);
  nand _75438_ (_24573_, _24572_, _24568_);
  or _75439_ (_24574_, _24572_, _24568_);
  and _75440_ (_24575_, _24574_, _08798_);
  nand _75441_ (_24576_, _24575_, _24573_);
  nand _75442_ (_24578_, _24576_, _24556_);
  or _75443_ (_24579_, _24578_, _24552_);
  or _75444_ (_24580_, _24556_, _23211_);
  and _75445_ (_24581_, _24580_, _43000_);
  and _75446_ (_24582_, _24581_, _24579_);
  or _75447_ (_24583_, _24582_, _23144_);
  and _75448_ (_43570_, _24583_, _41806_);
  or _75449_ (_24584_, _05245_, \oc8051_golden_model_1.PSW [1]);
  and _75450_ (_24585_, _12213_, _05245_);
  not _75451_ (_24586_, _24585_);
  and _75452_ (_24588_, _24586_, _24584_);
  or _75453_ (_24589_, _24588_, _04081_);
  nand _75454_ (_24590_, _05245_, _03274_);
  and _75455_ (_24591_, _24590_, _24584_);
  and _75456_ (_24592_, _24591_, _04409_);
  not _75457_ (_24593_, \oc8051_golden_model_1.PSW [1]);
  nor _75458_ (_24594_, _04409_, _24593_);
  or _75459_ (_24595_, _24594_, _03610_);
  or _75460_ (_24596_, _24595_, _24592_);
  and _75461_ (_24597_, _24596_, _04055_);
  and _75462_ (_24599_, _24597_, _24589_);
  and _75463_ (_24600_, _12224_, _05901_);
  nor _75464_ (_24601_, _05901_, _24593_);
  or _75465_ (_24602_, _24601_, _03723_);
  or _75466_ (_24603_, _24602_, _24600_);
  and _75467_ (_24604_, _24603_, _14265_);
  or _75468_ (_24605_, _24604_, _24599_);
  nor _75469_ (_24606_, _05245_, _24593_);
  and _75470_ (_24607_, _05245_, _06764_);
  or _75471_ (_24608_, _24607_, _24606_);
  or _75472_ (_24610_, _24608_, _03996_);
  and _75473_ (_24611_, _24610_, _24605_);
  or _75474_ (_24612_, _24611_, _03729_);
  or _75475_ (_24613_, _24591_, _03737_);
  and _75476_ (_24614_, _24613_, _03736_);
  and _75477_ (_24615_, _24614_, _24612_);
  and _75478_ (_24616_, _12211_, _05901_);
  or _75479_ (_24617_, _24616_, _24601_);
  and _75480_ (_24618_, _24617_, _03714_);
  or _75481_ (_24619_, _24618_, _03719_);
  or _75482_ (_24622_, _24619_, _24615_);
  and _75483_ (_24623_, _24600_, _12239_);
  or _75484_ (_24624_, _24601_, _06840_);
  or _75485_ (_24625_, _24624_, _24623_);
  and _75486_ (_24626_, _24625_, _24622_);
  and _75487_ (_24627_, _24626_, _03710_);
  not _75488_ (_24628_, _05901_);
  nor _75489_ (_24629_, _12256_, _24628_);
  or _75490_ (_24630_, _24601_, _24629_);
  and _75491_ (_24631_, _24630_, _03505_);
  or _75492_ (_24633_, _24631_, _07390_);
  or _75493_ (_24634_, _24633_, _24627_);
  or _75494_ (_24635_, _24608_, _06838_);
  and _75495_ (_24636_, _24635_, _24634_);
  or _75496_ (_24637_, _24636_, _04481_);
  and _75497_ (_24638_, _06501_, _05245_);
  or _75498_ (_24639_, _24606_, _07400_);
  or _75499_ (_24640_, _24639_, _24638_);
  and _75500_ (_24641_, _24640_, _03589_);
  and _75501_ (_24642_, _24641_, _24637_);
  nor _75502_ (_24644_, _12313_, _09661_);
  or _75503_ (_24645_, _24644_, _24606_);
  and _75504_ (_24646_, _24645_, _03222_);
  or _75505_ (_24647_, _24646_, _24642_);
  and _75506_ (_24648_, _24647_, _03602_);
  or _75507_ (_24649_, _12327_, _09661_);
  and _75508_ (_24650_, _24649_, _03600_);
  nand _75509_ (_24651_, _05245_, _04303_);
  and _75510_ (_24652_, _24651_, _03601_);
  or _75511_ (_24653_, _24652_, _24650_);
  and _75512_ (_24655_, _24653_, _24584_);
  or _75513_ (_24656_, _24655_, _24648_);
  and _75514_ (_24657_, _24656_, _07778_);
  or _75515_ (_24658_, _12333_, _09661_);
  and _75516_ (_24659_, _24584_, _03780_);
  and _75517_ (_24660_, _24659_, _24658_);
  or _75518_ (_24661_, _24660_, _24657_);
  and _75519_ (_24662_, _24661_, _07777_);
  or _75520_ (_24663_, _12207_, _09661_);
  and _75521_ (_24664_, _24584_, _03622_);
  and _75522_ (_24666_, _24664_, _24663_);
  or _75523_ (_24667_, _24666_, _24662_);
  and _75524_ (_24668_, _24667_, _06828_);
  or _75525_ (_24669_, _24606_, _05618_);
  and _75526_ (_24670_, _24591_, _03790_);
  and _75527_ (_24671_, _24670_, _24669_);
  or _75528_ (_24672_, _24671_, _24668_);
  and _75529_ (_24673_, _24672_, _03786_);
  or _75530_ (_24674_, _24651_, _05618_);
  and _75531_ (_24675_, _24584_, _03624_);
  and _75532_ (_24677_, _24675_, _24674_);
  or _75533_ (_24678_, _24590_, _05618_);
  and _75534_ (_24679_, _24584_, _03785_);
  and _75535_ (_24680_, _24679_, _24678_);
  or _75536_ (_24681_, _24680_, _03815_);
  or _75537_ (_24682_, _24681_, _24677_);
  or _75538_ (_24683_, _24682_, _24673_);
  or _75539_ (_24684_, _24588_, _04246_);
  and _75540_ (_24685_, _24684_, _03823_);
  and _75541_ (_24686_, _24685_, _24683_);
  and _75542_ (_24688_, _24617_, _03453_);
  or _75543_ (_24689_, _24688_, _03447_);
  or _75544_ (_24690_, _24689_, _24686_);
  or _75545_ (_24691_, _24606_, _03514_);
  or _75546_ (_24692_, _24691_, _24585_);
  and _75547_ (_24693_, _24692_, _24690_);
  or _75548_ (_24694_, _24693_, _43004_);
  or _75549_ (_24695_, _43000_, \oc8051_golden_model_1.PSW [1]);
  and _75550_ (_24696_, _24695_, _41806_);
  and _75551_ (_43571_, _24696_, _24694_);
  and _75552_ (_24698_, _07821_, \oc8051_golden_model_1.ACC [7]);
  nor _75553_ (_24699_, _07821_, \oc8051_golden_model_1.ACC [7]);
  nor _75554_ (_24700_, _24699_, _10295_);
  nor _75555_ (_24701_, _24700_, _24698_);
  nand _75556_ (_24702_, _24701_, _07890_);
  and _75557_ (_24703_, _24698_, _07887_);
  nor _75558_ (_24704_, _24703_, _07898_);
  and _75559_ (_24705_, _24704_, _24702_);
  not _75560_ (_24706_, \oc8051_golden_model_1.PSW [2]);
  nor _75561_ (_24707_, _05245_, _24706_);
  not _75562_ (_24709_, _24707_);
  or _75563_ (_24710_, _12519_, _09661_);
  and _75564_ (_24711_, _24710_, _24709_);
  or _75565_ (_24712_, _24711_, _03589_);
  or _75566_ (_24713_, _09661_, _04875_);
  and _75567_ (_24714_, _24713_, _24709_);
  and _75568_ (_24715_, _24714_, _07390_);
  not _75569_ (_24716_, _08050_);
  nor _75570_ (_24717_, _07987_, \oc8051_golden_model_1.ACC [7]);
  and _75571_ (_24718_, _07987_, \oc8051_golden_model_1.ACC [7]);
  nor _75572_ (_24720_, _24718_, _24717_);
  and _75573_ (_24721_, _24720_, _10197_);
  nor _75574_ (_24722_, _24720_, _10197_);
  or _75575_ (_24723_, _24722_, _24721_);
  or _75576_ (_24724_, _24723_, _24716_);
  nand _75577_ (_24725_, _24723_, _24716_);
  and _75578_ (_24726_, _24725_, _24724_);
  and _75579_ (_24727_, _24726_, _08051_);
  not _75580_ (_24728_, _07822_);
  and _75581_ (_24729_, _10183_, _24728_);
  nor _75582_ (_24731_, _10183_, _24728_);
  nor _75583_ (_24732_, _24731_, _24729_);
  nor _75584_ (_24733_, _24732_, _08177_);
  and _75585_ (_24734_, _24732_, _08177_);
  or _75586_ (_24735_, _24734_, _24733_);
  or _75587_ (_24736_, _24735_, _08059_);
  nor _75588_ (_24737_, _05901_, _24706_);
  and _75589_ (_24738_, _12409_, _05901_);
  nor _75590_ (_24739_, _24738_, _24737_);
  or _75591_ (_24740_, _24739_, _03736_);
  and _75592_ (_24742_, _24714_, _03723_);
  nor _75593_ (_24743_, _12416_, _09661_);
  nor _75594_ (_24744_, _24743_, _24707_);
  and _75595_ (_24745_, _24744_, _03610_);
  and _75596_ (_24746_, _05245_, \oc8051_golden_model_1.ACC [2]);
  nor _75597_ (_24747_, _24746_, _24707_);
  or _75598_ (_24748_, _24747_, _09029_);
  or _75599_ (_24749_, _04409_, _24706_);
  and _75600_ (_24750_, _24749_, _04081_);
  and _75601_ (_24751_, _24750_, _24748_);
  or _75602_ (_24753_, _24751_, _03715_);
  or _75603_ (_24754_, _24753_, _24745_);
  not _75604_ (_24755_, _24737_);
  nand _75605_ (_24756_, _12411_, _05901_);
  and _75606_ (_24757_, _24756_, _24755_);
  or _75607_ (_24758_, _24757_, _04055_);
  and _75608_ (_24759_, _24758_, _03996_);
  and _75609_ (_24760_, _24759_, _24754_);
  or _75610_ (_24761_, _24760_, _24742_);
  and _75611_ (_24762_, _24761_, _03737_);
  and _75612_ (_24764_, _24747_, _03729_);
  or _75613_ (_24765_, _24764_, _03714_);
  or _75614_ (_24766_, _24765_, _24762_);
  and _75615_ (_24767_, _24766_, _24740_);
  or _75616_ (_24768_, _24767_, _03719_);
  and _75617_ (_24769_, _24755_, _10084_);
  or _75618_ (_24770_, _24769_, _06840_);
  or _75619_ (_24771_, _24770_, _24757_);
  and _75620_ (_24772_, _24771_, _06875_);
  and _75621_ (_24773_, _24772_, _24768_);
  or _75622_ (_24775_, _14294_, _14181_);
  or _75623_ (_24776_, _24775_, _14408_);
  or _75624_ (_24777_, _24776_, _14527_);
  or _75625_ (_24778_, _24777_, _14643_);
  or _75626_ (_24779_, _24778_, _14758_);
  or _75627_ (_24780_, _24779_, _07386_);
  nor _75628_ (_24781_, _24780_, _14875_);
  or _75629_ (_24782_, _24781_, _08060_);
  or _75630_ (_24783_, _24782_, _24773_);
  and _75631_ (_24784_, _24783_, _10201_);
  and _75632_ (_24786_, _24784_, _24736_);
  or _75633_ (_24787_, _24786_, _03761_);
  or _75634_ (_24788_, _24787_, _24727_);
  nor _75635_ (_24789_, _08520_, \oc8051_golden_model_1.ACC [7]);
  and _75636_ (_24790_, _08520_, \oc8051_golden_model_1.ACC [7]);
  nor _75637_ (_24791_, _24790_, _24789_);
  not _75638_ (_24792_, _24791_);
  or _75639_ (_24793_, _24792_, _10227_);
  nand _75640_ (_24794_, _24792_, _10227_);
  and _75641_ (_24795_, _24794_, _24793_);
  nand _75642_ (_24797_, _24795_, _23615_);
  or _75643_ (_24798_, _24795_, _23615_);
  and _75644_ (_24799_, _24798_, _24797_);
  or _75645_ (_24800_, _24799_, _03766_);
  and _75646_ (_24801_, _24800_, _07914_);
  and _75647_ (_24802_, _24801_, _24788_);
  nor _75648_ (_24803_, _07919_, \oc8051_golden_model_1.ACC [7]);
  and _75649_ (_24804_, _07919_, \oc8051_golden_model_1.ACC [7]);
  nor _75650_ (_24805_, _24804_, _24803_);
  nor _75651_ (_24806_, _24805_, _10239_);
  and _75652_ (_24808_, _24805_, _10239_);
  or _75653_ (_24809_, _24808_, _24806_);
  or _75654_ (_24810_, _24809_, _07984_);
  nand _75655_ (_24811_, _24809_, _07984_);
  and _75656_ (_24812_, _24811_, _24810_);
  and _75657_ (_24813_, _24812_, _07913_);
  or _75658_ (_24814_, _24813_, _03505_);
  or _75659_ (_24815_, _24814_, _24802_);
  or _75660_ (_24816_, _12461_, _24628_);
  and _75661_ (_24817_, _24816_, _24755_);
  or _75662_ (_24819_, _24817_, _03710_);
  and _75663_ (_24820_, _24819_, _06838_);
  and _75664_ (_24821_, _24820_, _24815_);
  or _75665_ (_24822_, _24821_, _24715_);
  and _75666_ (_24823_, _24822_, _07400_);
  nand _75667_ (_24824_, _06637_, _05245_);
  nor _75668_ (_24825_, _24707_, _07400_);
  and _75669_ (_24826_, _24825_, _24824_);
  or _75670_ (_24827_, _24826_, _03222_);
  or _75671_ (_24828_, _24827_, _24823_);
  and _75672_ (_24830_, _24828_, _24712_);
  or _75673_ (_24831_, _24830_, _07405_);
  nor _75674_ (_24832_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and _75675_ (_24833_, _24832_, _07431_);
  nand _75676_ (_24834_, _24833_, _07405_);
  and _75677_ (_24835_, _24834_, _03602_);
  and _75678_ (_24836_, _24835_, _24831_);
  nand _75679_ (_24837_, _12533_, _05245_);
  nor _75680_ (_24838_, _24707_, _07766_);
  and _75681_ (_24839_, _24838_, _24837_);
  and _75682_ (_24841_, _05245_, _06332_);
  nor _75683_ (_24842_, _24841_, _24707_);
  and _75684_ (_24843_, _24842_, _03601_);
  or _75685_ (_24844_, _24843_, _03780_);
  or _75686_ (_24845_, _24844_, _24839_);
  or _75687_ (_24846_, _24845_, _24836_);
  nand _75688_ (_24847_, _12539_, _05245_);
  and _75689_ (_24848_, _24847_, _24709_);
  or _75690_ (_24849_, _24848_, _07778_);
  and _75691_ (_24850_, _24849_, _24846_);
  or _75692_ (_24852_, _24850_, _03622_);
  and _75693_ (_24853_, _24709_, _05717_);
  or _75694_ (_24854_, _24842_, _07777_);
  or _75695_ (_24855_, _24854_, _24853_);
  and _75696_ (_24856_, _24855_, _24852_);
  or _75697_ (_24857_, _24856_, _03790_);
  or _75698_ (_24858_, _24747_, _06828_);
  or _75699_ (_24859_, _24858_, _24853_);
  and _75700_ (_24860_, _24859_, _07795_);
  and _75701_ (_24861_, _24860_, _24857_);
  or _75702_ (_24863_, _12532_, _09661_);
  nor _75703_ (_24864_, _24707_, _07795_);
  and _75704_ (_24865_, _24864_, _24863_);
  or _75705_ (_24866_, _24865_, _03785_);
  or _75706_ (_24867_, _24866_, _24861_);
  or _75707_ (_24868_, _12538_, _09661_);
  and _75708_ (_24869_, _24868_, _24709_);
  or _75709_ (_24870_, _24869_, _07793_);
  and _75710_ (_24871_, _24870_, _07898_);
  and _75711_ (_24872_, _24871_, _24867_);
  or _75712_ (_24874_, _24872_, _24705_);
  and _75713_ (_24875_, _24874_, _08477_);
  nand _75714_ (_24876_, _24718_, _08499_);
  nor _75715_ (_24877_, _24717_, _10301_);
  nor _75716_ (_24878_, _24877_, _24718_);
  nand _75717_ (_24879_, _24878_, _08502_);
  and _75718_ (_24880_, _24879_, _24876_);
  and _75719_ (_24881_, _24880_, _08475_);
  or _75720_ (_24882_, _24881_, _03776_);
  or _75721_ (_24883_, _24882_, _24875_);
  nand _75722_ (_24885_, _24790_, _08580_);
  nor _75723_ (_24886_, _24792_, _10307_);
  nor _75724_ (_24887_, _24886_, _24790_);
  nand _75725_ (_24888_, _24887_, _08583_);
  and _75726_ (_24889_, _24888_, _24885_);
  or _75727_ (_24890_, _24889_, _03777_);
  and _75728_ (_24891_, _24890_, _08589_);
  and _75729_ (_24892_, _24891_, _24883_);
  nand _75730_ (_24893_, _24804_, _08610_);
  nor _75731_ (_24894_, _24803_, _10313_);
  or _75732_ (_24896_, _24804_, _24358_);
  or _75733_ (_24897_, _24896_, _24894_);
  and _75734_ (_24898_, _24897_, _24893_);
  and _75735_ (_24899_, _24898_, _08506_);
  or _75736_ (_24900_, _24899_, _08618_);
  or _75737_ (_24901_, _24900_, _24892_);
  nor _75738_ (_24902_, _08693_, _08374_);
  nand _75739_ (_24903_, _10331_, _08618_);
  or _75740_ (_24904_, _24903_, _24902_);
  and _75741_ (_24905_, _24904_, _08624_);
  nand _75742_ (_24907_, _24905_, _24901_);
  nor _75743_ (_24908_, _08657_, _24176_);
  and _75744_ (_24909_, _08657_, _08399_);
  or _75745_ (_24910_, _24909_, _08624_);
  or _75746_ (_24911_, _24910_, _24908_);
  and _75747_ (_24912_, _24911_, _08702_);
  and _75748_ (_24913_, _24912_, _24907_);
  or _75749_ (_24914_, _08725_, _08188_);
  and _75750_ (_24915_, _24914_, _10354_);
  or _75751_ (_24916_, _08765_, _08406_);
  and _75752_ (_24918_, _10349_, _24916_);
  or _75753_ (_24919_, _24918_, _03815_);
  or _75754_ (_24920_, _24919_, _24915_);
  or _75755_ (_24921_, _24920_, _24913_);
  nand _75756_ (_24922_, _24744_, _03815_);
  and _75757_ (_24923_, _24922_, _03823_);
  and _75758_ (_24924_, _24923_, _24921_);
  nor _75759_ (_24925_, _24739_, _03823_);
  or _75760_ (_24926_, _24925_, _03447_);
  or _75761_ (_24927_, _24926_, _24924_);
  and _75762_ (_24929_, _12592_, _05245_);
  or _75763_ (_24930_, _24707_, _03514_);
  or _75764_ (_24931_, _24930_, _24929_);
  and _75765_ (_24932_, _24931_, _24927_);
  or _75766_ (_24933_, _24932_, _43004_);
  or _75767_ (_24934_, _43000_, \oc8051_golden_model_1.PSW [2]);
  and _75768_ (_24935_, _24934_, _41806_);
  and _75769_ (_43572_, _24935_, _24933_);
  nor _75770_ (_24936_, _05245_, _05018_);
  and _75771_ (_24937_, _05245_, _06276_);
  nor _75772_ (_24939_, _24937_, _24936_);
  and _75773_ (_24940_, _24939_, _03601_);
  nor _75774_ (_24941_, _09661_, _05005_);
  nor _75775_ (_24942_, _24941_, _24936_);
  and _75776_ (_24943_, _24942_, _07390_);
  and _75777_ (_24944_, _05245_, \oc8051_golden_model_1.ACC [3]);
  nor _75778_ (_24945_, _24944_, _24936_);
  nor _75779_ (_24946_, _24945_, _09029_);
  nor _75780_ (_24947_, _04409_, _05018_);
  or _75781_ (_24948_, _24947_, _24946_);
  and _75782_ (_24950_, _24948_, _04081_);
  nor _75783_ (_24951_, _12627_, _09661_);
  nor _75784_ (_24952_, _24951_, _24936_);
  nor _75785_ (_24953_, _24952_, _04081_);
  or _75786_ (_24954_, _24953_, _24950_);
  and _75787_ (_24955_, _24954_, _04055_);
  nor _75788_ (_24956_, _05901_, _05018_);
  and _75789_ (_24957_, _12631_, _05901_);
  nor _75790_ (_24958_, _24957_, _24956_);
  nor _75791_ (_24959_, _24958_, _04055_);
  or _75792_ (_24961_, _24959_, _03723_);
  or _75793_ (_24962_, _24961_, _24955_);
  nand _75794_ (_24963_, _24942_, _03723_);
  and _75795_ (_24964_, _24963_, _24962_);
  and _75796_ (_24965_, _24964_, _03737_);
  nor _75797_ (_24966_, _24945_, _03737_);
  or _75798_ (_24967_, _24966_, _24965_);
  and _75799_ (_24968_, _24967_, _03736_);
  and _75800_ (_24969_, _12641_, _05901_);
  nor _75801_ (_24970_, _24969_, _24956_);
  nor _75802_ (_24972_, _24970_, _03736_);
  or _75803_ (_24973_, _24972_, _03719_);
  or _75804_ (_24974_, _24973_, _24968_);
  nor _75805_ (_24975_, _24956_, _12648_);
  nor _75806_ (_24976_, _24975_, _24958_);
  or _75807_ (_24977_, _24976_, _06840_);
  and _75808_ (_24978_, _24977_, _03710_);
  and _75809_ (_24979_, _24978_, _24974_);
  nor _75810_ (_24980_, _12612_, _24628_);
  nor _75811_ (_24981_, _24980_, _24956_);
  nor _75812_ (_24983_, _24981_, _03710_);
  nor _75813_ (_24984_, _24983_, _07390_);
  not _75814_ (_24985_, _24984_);
  nor _75815_ (_24986_, _24985_, _24979_);
  nor _75816_ (_24987_, _24986_, _24943_);
  nor _75817_ (_24988_, _24987_, _04481_);
  and _75818_ (_24989_, _06592_, _05245_);
  nor _75819_ (_24990_, _24936_, _07400_);
  not _75820_ (_24991_, _24990_);
  nor _75821_ (_24992_, _24991_, _24989_);
  or _75822_ (_24994_, _24992_, _03222_);
  nor _75823_ (_24995_, _24994_, _24988_);
  nor _75824_ (_24996_, _12718_, _09661_);
  nor _75825_ (_24997_, _24936_, _24996_);
  nor _75826_ (_24998_, _24997_, _03589_);
  or _75827_ (_24999_, _24998_, _03601_);
  nor _75828_ (_25000_, _24999_, _24995_);
  nor _75829_ (_25001_, _25000_, _24940_);
  or _75830_ (_25002_, _25001_, _03600_);
  and _75831_ (_25003_, _12733_, _05245_);
  or _75832_ (_25005_, _25003_, _24936_);
  or _75833_ (_25006_, _25005_, _07766_);
  and _75834_ (_25007_, _25006_, _07778_);
  and _75835_ (_25008_, _25007_, _25002_);
  and _75836_ (_25009_, _12739_, _05245_);
  nor _75837_ (_25010_, _25009_, _24936_);
  nor _75838_ (_25011_, _25010_, _07778_);
  nor _75839_ (_25012_, _25011_, _25008_);
  nor _75840_ (_25013_, _25012_, _03622_);
  nor _75841_ (_25014_, _24936_, _05567_);
  not _75842_ (_25016_, _25014_);
  nor _75843_ (_25017_, _24939_, _07777_);
  and _75844_ (_25018_, _25017_, _25016_);
  nor _75845_ (_25019_, _25018_, _25013_);
  nor _75846_ (_25020_, _25019_, _03790_);
  nor _75847_ (_25021_, _24945_, _06828_);
  and _75848_ (_25022_, _25021_, _25016_);
  nor _75849_ (_25023_, _25022_, _03624_);
  not _75850_ (_25024_, _25023_);
  nor _75851_ (_25025_, _25024_, _25020_);
  nor _75852_ (_25027_, _12732_, _09661_);
  or _75853_ (_25028_, _24936_, _07795_);
  nor _75854_ (_25029_, _25028_, _25027_);
  or _75855_ (_25030_, _25029_, _03785_);
  nor _75856_ (_25031_, _25030_, _25025_);
  nor _75857_ (_25032_, _12738_, _09661_);
  nor _75858_ (_25033_, _25032_, _24936_);
  nor _75859_ (_25034_, _25033_, _07793_);
  or _75860_ (_25035_, _25034_, _25031_);
  and _75861_ (_25036_, _25035_, _04246_);
  nor _75862_ (_25038_, _24952_, _04246_);
  or _75863_ (_25039_, _25038_, _25036_);
  and _75864_ (_25040_, _25039_, _03823_);
  nor _75865_ (_25041_, _24970_, _03823_);
  or _75866_ (_25042_, _25041_, _25040_);
  and _75867_ (_25043_, _25042_, _03514_);
  and _75868_ (_25044_, _12794_, _05245_);
  nor _75869_ (_25045_, _25044_, _24936_);
  nor _75870_ (_25046_, _25045_, _03514_);
  or _75871_ (_25047_, _25046_, _25043_);
  or _75872_ (_25049_, _25047_, _43004_);
  or _75873_ (_25050_, _43000_, \oc8051_golden_model_1.PSW [3]);
  and _75874_ (_25051_, _25050_, _41806_);
  and _75875_ (_43573_, _25051_, _25049_);
  not _75876_ (_25052_, \oc8051_golden_model_1.PSW [4]);
  nor _75877_ (_25053_, _05245_, _25052_);
  nor _75878_ (_25054_, _05777_, _09661_);
  nor _75879_ (_25055_, _25054_, _25053_);
  and _75880_ (_25056_, _25055_, _07390_);
  nor _75881_ (_25057_, _05901_, _25052_);
  and _75882_ (_25059_, _12827_, _05901_);
  nor _75883_ (_25060_, _25059_, _25057_);
  nor _75884_ (_25061_, _25060_, _03736_);
  and _75885_ (_25062_, _05245_, \oc8051_golden_model_1.ACC [4]);
  nor _75886_ (_25063_, _25062_, _25053_);
  nor _75887_ (_25064_, _25063_, _09029_);
  nor _75888_ (_25065_, _04409_, _25052_);
  or _75889_ (_25066_, _25065_, _25064_);
  and _75890_ (_25067_, _25066_, _04081_);
  nor _75891_ (_25068_, _12841_, _09661_);
  nor _75892_ (_25070_, _25068_, _25053_);
  nor _75893_ (_25071_, _25070_, _04081_);
  or _75894_ (_25072_, _25071_, _25067_);
  and _75895_ (_25073_, _25072_, _04055_);
  and _75896_ (_25074_, _12845_, _05901_);
  nor _75897_ (_25075_, _25074_, _25057_);
  nor _75898_ (_25076_, _25075_, _04055_);
  or _75899_ (_25077_, _25076_, _03723_);
  or _75900_ (_25078_, _25077_, _25073_);
  nand _75901_ (_25079_, _25055_, _03723_);
  and _75902_ (_25081_, _25079_, _25078_);
  and _75903_ (_25082_, _25081_, _03737_);
  nor _75904_ (_25083_, _25063_, _03737_);
  or _75905_ (_25084_, _25083_, _25082_);
  and _75906_ (_25085_, _25084_, _03736_);
  nor _75907_ (_25086_, _25085_, _25061_);
  nor _75908_ (_25087_, _25086_, _03719_);
  nor _75909_ (_25088_, _25057_, _12860_);
  or _75910_ (_25089_, _25075_, _06840_);
  nor _75911_ (_25090_, _25089_, _25088_);
  nor _75912_ (_25092_, _25090_, _25087_);
  nor _75913_ (_25093_, _25092_, _03505_);
  nor _75914_ (_25094_, _12825_, _24628_);
  nor _75915_ (_25095_, _25094_, _25057_);
  nor _75916_ (_25096_, _25095_, _03710_);
  nor _75917_ (_25097_, _25096_, _07390_);
  not _75918_ (_25098_, _25097_);
  nor _75919_ (_25099_, _25098_, _25093_);
  nor _75920_ (_25100_, _25099_, _25056_);
  nor _75921_ (_25101_, _25100_, _04481_);
  and _75922_ (_25102_, _06730_, _05245_);
  nor _75923_ (_25103_, _25053_, _07400_);
  not _75924_ (_25104_, _25103_);
  nor _75925_ (_25105_, _25104_, _25102_);
  nor _75926_ (_25106_, _25105_, _03222_);
  not _75927_ (_25107_, _25106_);
  nor _75928_ (_25108_, _25107_, _25101_);
  nor _75929_ (_25109_, _12933_, _09661_);
  nor _75930_ (_25110_, _25109_, _25053_);
  nor _75931_ (_25111_, _25110_, _03589_);
  or _75932_ (_25114_, _25111_, _08828_);
  or _75933_ (_25115_, _25114_, _25108_);
  and _75934_ (_25116_, _12821_, _05245_);
  or _75935_ (_25117_, _25053_, _07766_);
  or _75936_ (_25118_, _25117_, _25116_);
  and _75937_ (_25119_, _06298_, _05245_);
  nor _75938_ (_25120_, _25119_, _25053_);
  and _75939_ (_25121_, _25120_, _03601_);
  nor _75940_ (_25122_, _25121_, _03780_);
  and _75941_ (_25123_, _25122_, _25118_);
  and _75942_ (_25125_, _25123_, _25115_);
  and _75943_ (_25126_, _12817_, _05245_);
  nor _75944_ (_25127_, _25126_, _25053_);
  nor _75945_ (_25128_, _25127_, _07778_);
  nor _75946_ (_25129_, _25128_, _25125_);
  nor _75947_ (_25130_, _25129_, _03622_);
  nor _75948_ (_25131_, _25053_, _05825_);
  not _75949_ (_25132_, _25131_);
  nor _75950_ (_25133_, _25120_, _07777_);
  and _75951_ (_25134_, _25133_, _25132_);
  nor _75952_ (_25136_, _25134_, _25130_);
  nor _75953_ (_25137_, _25136_, _03790_);
  nor _75954_ (_25138_, _25063_, _06828_);
  and _75955_ (_25139_, _25138_, _25132_);
  nor _75956_ (_25140_, _25139_, _03624_);
  not _75957_ (_25141_, _25140_);
  nor _75958_ (_25142_, _25141_, _25137_);
  nor _75959_ (_25143_, _12819_, _09661_);
  or _75960_ (_25144_, _25053_, _07795_);
  nor _75961_ (_25145_, _25144_, _25143_);
  or _75962_ (_25146_, _25145_, _03785_);
  nor _75963_ (_25147_, _25146_, _25142_);
  nor _75964_ (_25148_, _12816_, _09661_);
  nor _75965_ (_25149_, _25148_, _25053_);
  nor _75966_ (_25150_, _25149_, _07793_);
  or _75967_ (_25151_, _25150_, _25147_);
  and _75968_ (_25152_, _25151_, _04246_);
  nor _75969_ (_25153_, _25070_, _04246_);
  or _75970_ (_25154_, _25153_, _25152_);
  and _75971_ (_25155_, _25154_, _03823_);
  nor _75972_ (_25158_, _25060_, _03823_);
  or _75973_ (_25159_, _25158_, _25155_);
  and _75974_ (_25160_, _25159_, _03514_);
  and _75975_ (_25161_, _13003_, _05245_);
  nor _75976_ (_25162_, _25161_, _25053_);
  nor _75977_ (_25163_, _25162_, _03514_);
  or _75978_ (_25164_, _25163_, _25160_);
  or _75979_ (_25165_, _25164_, _43004_);
  or _75980_ (_25166_, _43000_, \oc8051_golden_model_1.PSW [4]);
  and _75981_ (_25167_, _25166_, _41806_);
  and _75982_ (_43574_, _25167_, _25165_);
  not _75983_ (_25169_, \oc8051_golden_model_1.PSW [5]);
  nor _75984_ (_25170_, _05245_, _25169_);
  and _75985_ (_25171_, _06684_, _05245_);
  or _75986_ (_25172_, _25171_, _25170_);
  and _75987_ (_25173_, _25172_, _04481_);
  and _75988_ (_25174_, _05245_, \oc8051_golden_model_1.ACC [5]);
  nor _75989_ (_25175_, _25174_, _25170_);
  nor _75990_ (_25176_, _25175_, _09029_);
  nor _75991_ (_25177_, _04409_, _25169_);
  or _75992_ (_25178_, _25177_, _25176_);
  and _75993_ (_25179_, _25178_, _04081_);
  nor _75994_ (_25180_, _13014_, _09661_);
  nor _75995_ (_25181_, _25180_, _25170_);
  nor _75996_ (_25182_, _25181_, _04081_);
  or _75997_ (_25183_, _25182_, _25179_);
  and _75998_ (_25184_, _25183_, _04055_);
  nor _75999_ (_25185_, _05901_, _25169_);
  and _76000_ (_25186_, _13037_, _05901_);
  nor _76001_ (_25187_, _25186_, _25185_);
  nor _76002_ (_25190_, _25187_, _04055_);
  or _76003_ (_25191_, _25190_, _03723_);
  or _76004_ (_25192_, _25191_, _25184_);
  nor _76005_ (_25193_, _05469_, _09661_);
  nor _76006_ (_25194_, _25193_, _25170_);
  nand _76007_ (_25195_, _25194_, _03723_);
  and _76008_ (_25196_, _25195_, _25192_);
  and _76009_ (_25197_, _25196_, _03737_);
  nor _76010_ (_25198_, _25175_, _03737_);
  or _76011_ (_25199_, _25198_, _25197_);
  and _76012_ (_25201_, _25199_, _03736_);
  and _76013_ (_25202_, _13047_, _05901_);
  nor _76014_ (_25203_, _25202_, _25185_);
  nor _76015_ (_25204_, _25203_, _03736_);
  or _76016_ (_25205_, _25204_, _25201_);
  and _76017_ (_25206_, _25205_, _06840_);
  nor _76018_ (_25207_, _25185_, _13054_);
  nor _76019_ (_25208_, _25207_, _25187_);
  and _76020_ (_25209_, _25208_, _03719_);
  or _76021_ (_25210_, _25209_, _25206_);
  and _76022_ (_25212_, _25210_, _03710_);
  nor _76023_ (_25213_, _13020_, _24628_);
  nor _76024_ (_25214_, _25213_, _25185_);
  nor _76025_ (_25215_, _25214_, _03710_);
  nor _76026_ (_25216_, _25215_, _07390_);
  not _76027_ (_25217_, _25216_);
  nor _76028_ (_25218_, _25217_, _25212_);
  and _76029_ (_25219_, _25194_, _07390_);
  or _76030_ (_25220_, _25219_, _04481_);
  nor _76031_ (_25221_, _25220_, _25218_);
  or _76032_ (_25223_, _25221_, _25173_);
  and _76033_ (_25224_, _25223_, _03589_);
  nor _76034_ (_25225_, _13127_, _09661_);
  nor _76035_ (_25226_, _25225_, _25170_);
  nor _76036_ (_25227_, _25226_, _03589_);
  or _76037_ (_25228_, _25227_, _08828_);
  or _76038_ (_25229_, _25228_, _25224_);
  and _76039_ (_25230_, _13141_, _05245_);
  or _76040_ (_25231_, _25170_, _07766_);
  or _76041_ (_25232_, _25231_, _25230_);
  and _76042_ (_25233_, _06306_, _05245_);
  nor _76043_ (_25234_, _25233_, _25170_);
  and _76044_ (_25235_, _25234_, _03601_);
  nor _76045_ (_25236_, _25235_, _03780_);
  and _76046_ (_25237_, _25236_, _25232_);
  and _76047_ (_25238_, _25237_, _25229_);
  and _76048_ (_25239_, _13147_, _05245_);
  nor _76049_ (_25240_, _25239_, _25170_);
  nor _76050_ (_25241_, _25240_, _07778_);
  nor _76051_ (_25242_, _25241_, _25238_);
  nor _76052_ (_25245_, _25242_, _03622_);
  nor _76053_ (_25246_, _25170_, _05518_);
  not _76054_ (_25247_, _25246_);
  nor _76055_ (_25248_, _25234_, _07777_);
  and _76056_ (_25249_, _25248_, _25247_);
  nor _76057_ (_25250_, _25249_, _25245_);
  nor _76058_ (_25251_, _25250_, _03790_);
  nor _76059_ (_25252_, _25175_, _06828_);
  and _76060_ (_25253_, _25252_, _25247_);
  nor _76061_ (_25254_, _25253_, _03624_);
  not _76062_ (_25256_, _25254_);
  nor _76063_ (_25257_, _25256_, _25251_);
  nor _76064_ (_25258_, _13140_, _09661_);
  or _76065_ (_25259_, _25170_, _07795_);
  nor _76066_ (_25260_, _25259_, _25258_);
  or _76067_ (_25261_, _25260_, _03785_);
  nor _76068_ (_25262_, _25261_, _25257_);
  nor _76069_ (_25263_, _13146_, _09661_);
  nor _76070_ (_25264_, _25263_, _25170_);
  nor _76071_ (_25265_, _25264_, _07793_);
  or _76072_ (_25267_, _25265_, _25262_);
  and _76073_ (_25268_, _25267_, _04246_);
  nor _76074_ (_25269_, _25181_, _04246_);
  or _76075_ (_25270_, _25269_, _25268_);
  and _76076_ (_25271_, _25270_, _03823_);
  nor _76077_ (_25272_, _25203_, _03823_);
  or _76078_ (_25273_, _25272_, _25271_);
  and _76079_ (_25274_, _25273_, _03514_);
  and _76080_ (_25275_, _13199_, _05245_);
  nor _76081_ (_25276_, _25275_, _25170_);
  nor _76082_ (_25278_, _25276_, _03514_);
  or _76083_ (_25279_, _25278_, _25274_);
  or _76084_ (_25280_, _25279_, _43004_);
  or _76085_ (_25281_, _43000_, \oc8051_golden_model_1.PSW [5]);
  and _76086_ (_25282_, _25281_, _41806_);
  and _76087_ (_43575_, _25282_, _25280_);
  not _76088_ (_25283_, _08574_);
  nor _76089_ (_25284_, _25283_, _08516_);
  nor _76090_ (_25285_, _25284_, _03777_);
  nor _76091_ (_25286_, _05245_, _15859_);
  nor _76092_ (_25288_, _05363_, _09661_);
  nor _76093_ (_25289_, _25288_, _25286_);
  and _76094_ (_25290_, _25289_, _07390_);
  nor _76095_ (_25291_, _08516_, _03766_);
  not _76096_ (_25292_, _25291_);
  nor _76097_ (_25293_, _25292_, _10223_);
  nor _76098_ (_25294_, _08042_, _08006_);
  or _76099_ (_25295_, _25294_, _10201_);
  or _76100_ (_25296_, _08059_, _07834_);
  nor _76101_ (_25297_, _25296_, _08173_);
  nor _76102_ (_25299_, _05901_, _15859_);
  and _76103_ (_25300_, _13253_, _05901_);
  nor _76104_ (_25301_, _25300_, _25299_);
  nor _76105_ (_25302_, _25301_, _03736_);
  and _76106_ (_25303_, _05245_, \oc8051_golden_model_1.ACC [6]);
  nor _76107_ (_25304_, _25303_, _25286_);
  nor _76108_ (_25305_, _25304_, _09029_);
  nor _76109_ (_25306_, _04409_, _15859_);
  or _76110_ (_25307_, _25306_, _25305_);
  and _76111_ (_25308_, _25307_, _04081_);
  nor _76112_ (_25310_, _13242_, _09661_);
  nor _76113_ (_25311_, _25310_, _25286_);
  nor _76114_ (_25312_, _25311_, _04081_);
  or _76115_ (_25313_, _25312_, _25308_);
  and _76116_ (_25314_, _25313_, _04055_);
  and _76117_ (_25315_, _13229_, _05901_);
  nor _76118_ (_25316_, _25315_, _25299_);
  nor _76119_ (_25317_, _25316_, _04055_);
  or _76120_ (_25318_, _25317_, _03723_);
  or _76121_ (_25319_, _25318_, _25314_);
  nand _76122_ (_25321_, _25289_, _03723_);
  and _76123_ (_25322_, _25321_, _25319_);
  and _76124_ (_25323_, _25322_, _03737_);
  nor _76125_ (_25324_, _25304_, _03737_);
  or _76126_ (_25325_, _25324_, _25323_);
  and _76127_ (_25326_, _25325_, _03736_);
  nor _76128_ (_25327_, _25326_, _25302_);
  nor _76129_ (_25328_, _25327_, _03719_);
  nor _76130_ (_25329_, _25299_, _13260_);
  or _76131_ (_25330_, _25329_, _06840_);
  nor _76132_ (_25332_, _25330_, _25316_);
  or _76133_ (_25333_, _25332_, _08060_);
  nor _76134_ (_25334_, _25333_, _25328_);
  or _76135_ (_25335_, _25334_, _25297_);
  or _76136_ (_25336_, _25335_, _08051_);
  and _76137_ (_25337_, _25336_, _03766_);
  and _76138_ (_25338_, _25337_, _25295_);
  nor _76139_ (_25339_, _25338_, _25293_);
  nor _76140_ (_25340_, _25339_, _07913_);
  or _76141_ (_25341_, _07916_, _07914_);
  nor _76142_ (_25343_, _25341_, _07977_);
  or _76143_ (_25344_, _25343_, _03505_);
  nor _76144_ (_25345_, _25344_, _25340_);
  nor _76145_ (_25346_, _13226_, _24628_);
  nor _76146_ (_25347_, _25346_, _25299_);
  nor _76147_ (_25348_, _25347_, _03710_);
  nor _76148_ (_25349_, _25348_, _07390_);
  not _76149_ (_25350_, _25349_);
  nor _76150_ (_25351_, _25350_, _25345_);
  nor _76151_ (_25352_, _25351_, _25290_);
  nor _76152_ (_25354_, _25352_, _04481_);
  and _76153_ (_25355_, _06455_, _05245_);
  nor _76154_ (_25356_, _25286_, _07400_);
  not _76155_ (_25357_, _25356_);
  nor _76156_ (_25358_, _25357_, _25355_);
  nor _76157_ (_25359_, _25358_, _03222_);
  not _76158_ (_25360_, _25359_);
  nor _76159_ (_25361_, _25360_, _25354_);
  nor _76160_ (_25362_, _13332_, _09661_);
  nor _76161_ (_25363_, _25362_, _25286_);
  nor _76162_ (_25364_, _25363_, _03589_);
  or _76163_ (_25365_, _25364_, _08828_);
  or _76164_ (_25366_, _25365_, _25361_);
  and _76165_ (_25367_, _13347_, _05245_);
  or _76166_ (_25368_, _25286_, _07766_);
  or _76167_ (_25369_, _25368_, _25367_);
  and _76168_ (_25370_, _13339_, _05245_);
  nor _76169_ (_25371_, _25370_, _25286_);
  and _76170_ (_25372_, _25371_, _03601_);
  nor _76171_ (_25373_, _25372_, _03780_);
  and _76172_ (_25376_, _25373_, _25369_);
  and _76173_ (_25377_, _25376_, _25366_);
  and _76174_ (_25378_, _13353_, _05245_);
  nor _76175_ (_25379_, _25378_, _25286_);
  nor _76176_ (_25380_, _25379_, _07778_);
  nor _76177_ (_25381_, _25380_, _25377_);
  nor _76178_ (_25382_, _25381_, _03622_);
  nor _76179_ (_25383_, _25286_, _05412_);
  not _76180_ (_25384_, _25383_);
  nor _76181_ (_25385_, _25371_, _07777_);
  and _76182_ (_25387_, _25385_, _25384_);
  nor _76183_ (_25388_, _25387_, _25382_);
  nor _76184_ (_25389_, _25388_, _03790_);
  nor _76185_ (_25390_, _25304_, _06828_);
  and _76186_ (_25391_, _25390_, _25384_);
  or _76187_ (_25392_, _25391_, _25389_);
  and _76188_ (_25393_, _25392_, _07795_);
  nor _76189_ (_25394_, _13346_, _09661_);
  nor _76190_ (_25395_, _25394_, _25286_);
  nor _76191_ (_25396_, _25395_, _07795_);
  or _76192_ (_25398_, _25396_, _25393_);
  and _76193_ (_25399_, _25398_, _07793_);
  not _76194_ (_25400_, _07897_);
  nor _76195_ (_25401_, _13352_, _09661_);
  nor _76196_ (_25402_, _25401_, _25286_);
  nor _76197_ (_25403_, _25402_, _07793_);
  nor _76198_ (_25404_, _25403_, _25400_);
  not _76199_ (_25405_, _25404_);
  nor _76200_ (_25406_, _25405_, _25399_);
  not _76201_ (_25407_, _07834_);
  and _76202_ (_25409_, _07881_, _25407_);
  nor _76203_ (_25410_, _25409_, _07891_);
  nor _76204_ (_25411_, _25410_, _07898_);
  nor _76205_ (_25412_, _25411_, _25406_);
  nor _76206_ (_25413_, _25409_, _07892_);
  nor _76207_ (_25414_, _25413_, _08475_);
  not _76208_ (_25415_, _25414_);
  nor _76209_ (_25416_, _25415_, _25412_);
  nor _76210_ (_25417_, _08477_, _08006_);
  and _76211_ (_25418_, _25417_, _08493_);
  nor _76212_ (_25420_, _25418_, _03776_);
  not _76213_ (_25421_, _25420_);
  nor _76214_ (_25422_, _25421_, _25416_);
  nor _76215_ (_25423_, _25422_, _25285_);
  nor _76216_ (_25424_, _25423_, _08506_);
  not _76217_ (_25425_, _07916_);
  and _76218_ (_25426_, _08604_, _25425_);
  nor _76219_ (_25427_, _25426_, _08589_);
  nor _76220_ (_25428_, _25427_, _11907_);
  not _76221_ (_25429_, _25428_);
  nor _76222_ (_25431_, _25429_, _25424_);
  and _76223_ (_25432_, _08687_, _08618_);
  nor _76224_ (_25433_, _08651_, _08624_);
  or _76225_ (_25434_, _25433_, _03517_);
  nor _76226_ (_25435_, _25434_, _25432_);
  not _76227_ (_25436_, _25435_);
  nor _76228_ (_25437_, _25436_, _25431_);
  and _76229_ (_25438_, _08719_, _03517_);
  or _76230_ (_25439_, _25438_, _08701_);
  nor _76231_ (_25440_, _25439_, _25437_);
  nor _76232_ (_25442_, _08759_, _08734_);
  nor _76233_ (_25443_, _25442_, _25440_);
  and _76234_ (_25444_, _25443_, _04246_);
  nor _76235_ (_25445_, _25311_, _04246_);
  or _76236_ (_25446_, _25445_, _25444_);
  and _76237_ (_25447_, _25446_, _03823_);
  nor _76238_ (_25448_, _25301_, _03823_);
  or _76239_ (_25449_, _25448_, _25447_);
  and _76240_ (_25450_, _25449_, _03514_);
  and _76241_ (_25451_, _13402_, _05245_);
  nor _76242_ (_25453_, _25286_, _25451_);
  nor _76243_ (_25454_, _25453_, _03514_);
  or _76244_ (_25455_, _25454_, _25450_);
  or _76245_ (_25456_, _25455_, _43004_);
  or _76246_ (_25457_, _43000_, \oc8051_golden_model_1.PSW [6]);
  and _76247_ (_25458_, _25457_, _41806_);
  and _76248_ (_43576_, _25458_, _25456_);
  not _76249_ (_25459_, \oc8051_golden_model_1.PCON [0]);
  nor _76250_ (_25460_, _05212_, _25459_);
  nor _76251_ (_25461_, _05666_, _10377_);
  nor _76252_ (_25463_, _25461_, _25460_);
  and _76253_ (_25464_, _25463_, _17166_);
  and _76254_ (_25465_, _05212_, \oc8051_golden_model_1.ACC [0]);
  nor _76255_ (_25466_, _25465_, _25460_);
  nor _76256_ (_25467_, _25466_, _03737_);
  nor _76257_ (_25468_, _25467_, _07390_);
  nor _76258_ (_25469_, _25463_, _04081_);
  nor _76259_ (_25470_, _04409_, _25459_);
  nor _76260_ (_25471_, _25466_, _09029_);
  nor _76261_ (_25472_, _25471_, _25470_);
  nor _76262_ (_25474_, _25472_, _03610_);
  or _76263_ (_25475_, _25474_, _03723_);
  nor _76264_ (_25476_, _25475_, _25469_);
  or _76265_ (_25477_, _25476_, _03729_);
  and _76266_ (_25478_, _25477_, _25468_);
  and _76267_ (_25479_, _05212_, _04620_);
  and _76268_ (_25480_, _06838_, _03996_);
  or _76269_ (_25481_, _25480_, _25460_);
  nor _76270_ (_25482_, _25481_, _25479_);
  nor _76271_ (_25483_, _25482_, _25478_);
  nor _76272_ (_25485_, _25483_, _04481_);
  and _76273_ (_25486_, _06546_, _05212_);
  nor _76274_ (_25487_, _25460_, _07400_);
  not _76275_ (_25488_, _25487_);
  nor _76276_ (_25489_, _25488_, _25486_);
  nor _76277_ (_25490_, _25489_, _25485_);
  nor _76278_ (_25491_, _25490_, _03222_);
  nor _76279_ (_25492_, _12109_, _10377_);
  or _76280_ (_25493_, _25460_, _03589_);
  nor _76281_ (_25494_, _25493_, _25492_);
  or _76282_ (_25496_, _25494_, _03601_);
  nor _76283_ (_25497_, _25496_, _25491_);
  and _76284_ (_25498_, _05212_, _06274_);
  nor _76285_ (_25499_, _25498_, _25460_);
  nand _76286_ (_25500_, _25499_, _07766_);
  and _76287_ (_25501_, _25500_, _08828_);
  nor _76288_ (_25502_, _25501_, _25497_);
  and _76289_ (_25503_, _12124_, _05212_);
  nor _76290_ (_25504_, _25503_, _25460_);
  and _76291_ (_25505_, _25504_, _03600_);
  nor _76292_ (_25507_, _25505_, _25502_);
  nor _76293_ (_25508_, _25507_, _03780_);
  and _76294_ (_25509_, _12128_, _05212_);
  or _76295_ (_25510_, _25460_, _07778_);
  nor _76296_ (_25511_, _25510_, _25509_);
  or _76297_ (_25512_, _25511_, _03622_);
  nor _76298_ (_25513_, _25512_, _25508_);
  or _76299_ (_25514_, _25499_, _07777_);
  nor _76300_ (_25515_, _25514_, _25461_);
  nor _76301_ (_25516_, _25515_, _25513_);
  nor _76302_ (_25518_, _25516_, _03790_);
  and _76303_ (_25519_, _12005_, _05212_);
  or _76304_ (_25520_, _25519_, _25460_);
  and _76305_ (_25521_, _25520_, _03790_);
  or _76306_ (_25522_, _25521_, _25518_);
  and _76307_ (_25523_, _25522_, _07795_);
  nor _76308_ (_25524_, _12122_, _10377_);
  nor _76309_ (_25525_, _25524_, _25460_);
  nor _76310_ (_25526_, _25525_, _07795_);
  or _76311_ (_25527_, _25526_, _25523_);
  and _76312_ (_25529_, _25527_, _07793_);
  nor _76313_ (_25530_, _12003_, _10377_);
  nor _76314_ (_25531_, _25530_, _25460_);
  nor _76315_ (_25532_, _25531_, _07793_);
  nor _76316_ (_25533_, _25532_, _17166_);
  not _76317_ (_25534_, _25533_);
  nor _76318_ (_25535_, _25534_, _25529_);
  nor _76319_ (_25536_, _25535_, _25464_);
  or _76320_ (_25537_, _25536_, _43004_);
  or _76321_ (_25538_, _43000_, \oc8051_golden_model_1.PCON [0]);
  and _76322_ (_25539_, _25538_, _41806_);
  and _76323_ (_43579_, _25539_, _25537_);
  and _76324_ (_25540_, _06501_, _05212_);
  not _76325_ (_25541_, \oc8051_golden_model_1.PCON [1]);
  nor _76326_ (_25542_, _05212_, _25541_);
  nor _76327_ (_25543_, _25542_, _07400_);
  not _76328_ (_25544_, _25543_);
  nor _76329_ (_25545_, _25544_, _25540_);
  not _76330_ (_25546_, _25545_);
  nor _76331_ (_25547_, _05212_, \oc8051_golden_model_1.PCON [1]);
  and _76332_ (_25550_, _05212_, _03274_);
  nor _76333_ (_25551_, _25550_, _25547_);
  and _76334_ (_25552_, _25551_, _03729_);
  and _76335_ (_25553_, _25551_, _04409_);
  nor _76336_ (_25554_, _04409_, _25541_);
  or _76337_ (_25555_, _25554_, _25553_);
  and _76338_ (_25556_, _25555_, _04081_);
  and _76339_ (_25557_, _12213_, _05212_);
  nor _76340_ (_25558_, _25557_, _25547_);
  and _76341_ (_25559_, _25558_, _03610_);
  or _76342_ (_25561_, _25559_, _25556_);
  and _76343_ (_25562_, _25561_, _03996_);
  and _76344_ (_25563_, _05212_, _06764_);
  nor _76345_ (_25564_, _25563_, _25542_);
  nor _76346_ (_25565_, _25564_, _03996_);
  nor _76347_ (_25566_, _25565_, _25562_);
  nor _76348_ (_25567_, _25566_, _03729_);
  or _76349_ (_25568_, _25567_, _07390_);
  nor _76350_ (_25569_, _25568_, _25552_);
  and _76351_ (_25570_, _25564_, _07390_);
  nor _76352_ (_25572_, _25570_, _25569_);
  nor _76353_ (_25573_, _25572_, _04481_);
  nor _76354_ (_25574_, _25573_, _03222_);
  and _76355_ (_25575_, _25574_, _25546_);
  not _76356_ (_25576_, _25547_);
  and _76357_ (_25577_, _12313_, _05212_);
  nor _76358_ (_25578_, _25577_, _03589_);
  and _76359_ (_25579_, _25578_, _25576_);
  nor _76360_ (_25580_, _25579_, _25575_);
  nor _76361_ (_25581_, _25580_, _08828_);
  nor _76362_ (_25583_, _12327_, _10377_);
  nor _76363_ (_25584_, _25583_, _07766_);
  and _76364_ (_25585_, _05212_, _04303_);
  nor _76365_ (_25586_, _25585_, _05886_);
  nor _76366_ (_25587_, _25586_, _25584_);
  nor _76367_ (_25588_, _25587_, _25547_);
  nor _76368_ (_25589_, _25588_, _25581_);
  nor _76369_ (_25590_, _25589_, _03780_);
  nor _76370_ (_25591_, _12333_, _10377_);
  nor _76371_ (_25592_, _25591_, _07778_);
  and _76372_ (_25594_, _25592_, _25576_);
  nor _76373_ (_25595_, _25594_, _25590_);
  nor _76374_ (_25596_, _25595_, _03622_);
  nor _76375_ (_25597_, _12207_, _10377_);
  nor _76376_ (_25598_, _25597_, _07777_);
  and _76377_ (_25599_, _25598_, _25576_);
  nor _76378_ (_25600_, _25599_, _25596_);
  nor _76379_ (_25601_, _25600_, _03790_);
  nor _76380_ (_25602_, _25542_, _05618_);
  nor _76381_ (_25603_, _25602_, _06828_);
  and _76382_ (_25605_, _25603_, _25551_);
  nor _76383_ (_25606_, _25605_, _25601_);
  or _76384_ (_25607_, _25606_, _18499_);
  and _76385_ (_25608_, _25585_, _05617_);
  or _76386_ (_25609_, _25547_, _07795_);
  or _76387_ (_25610_, _25609_, _25608_);
  and _76388_ (_25611_, _25550_, _05617_);
  or _76389_ (_25612_, _25547_, _07793_);
  or _76390_ (_25613_, _25612_, _25611_);
  and _76391_ (_25614_, _25613_, _04246_);
  and _76392_ (_25616_, _25614_, _25610_);
  and _76393_ (_25617_, _25616_, _25607_);
  nor _76394_ (_25618_, _25558_, _04246_);
  nor _76395_ (_25619_, _25618_, _25617_);
  and _76396_ (_25620_, _25619_, _03514_);
  nor _76397_ (_25621_, _25557_, _25542_);
  nor _76398_ (_25622_, _25621_, _03514_);
  or _76399_ (_25623_, _25622_, _25620_);
  or _76400_ (_25624_, _25623_, _43004_);
  or _76401_ (_25625_, _43000_, \oc8051_golden_model_1.PCON [1]);
  and _76402_ (_25627_, _25625_, _41806_);
  and _76403_ (_43580_, _25627_, _25624_);
  not _76404_ (_25628_, \oc8051_golden_model_1.PCON [2]);
  nor _76405_ (_25629_, _05212_, _25628_);
  nor _76406_ (_25630_, _12538_, _10377_);
  nor _76407_ (_25631_, _25630_, _25629_);
  nor _76408_ (_25632_, _25631_, _07793_);
  and _76409_ (_25633_, _12539_, _05212_);
  nor _76410_ (_25634_, _25633_, _25629_);
  nor _76411_ (_25635_, _25634_, _07778_);
  nor _76412_ (_25637_, _10377_, _04875_);
  nor _76413_ (_25638_, _25637_, _25629_);
  and _76414_ (_25639_, _25638_, _07390_);
  and _76415_ (_25640_, _05212_, \oc8051_golden_model_1.ACC [2]);
  nor _76416_ (_25641_, _25640_, _25629_);
  nor _76417_ (_25642_, _25641_, _03737_);
  nor _76418_ (_25643_, _25641_, _09029_);
  nor _76419_ (_25644_, _04409_, _25628_);
  or _76420_ (_25645_, _25644_, _25643_);
  and _76421_ (_25646_, _25645_, _04081_);
  nor _76422_ (_25648_, _12416_, _10377_);
  nor _76423_ (_25649_, _25648_, _25629_);
  nor _76424_ (_25650_, _25649_, _04081_);
  or _76425_ (_25651_, _25650_, _25646_);
  and _76426_ (_25652_, _25651_, _03996_);
  nor _76427_ (_25653_, _25638_, _03996_);
  nor _76428_ (_25654_, _25653_, _25652_);
  nor _76429_ (_25655_, _25654_, _03729_);
  or _76430_ (_25656_, _25655_, _07390_);
  nor _76431_ (_25657_, _25656_, _25642_);
  nor _76432_ (_25659_, _25657_, _25639_);
  nor _76433_ (_25660_, _25659_, _04481_);
  and _76434_ (_25661_, _06637_, _05212_);
  nor _76435_ (_25662_, _25629_, _07400_);
  not _76436_ (_25663_, _25662_);
  nor _76437_ (_25664_, _25663_, _25661_);
  nor _76438_ (_25665_, _25664_, _03222_);
  not _76439_ (_25666_, _25665_);
  nor _76440_ (_25667_, _25666_, _25660_);
  nor _76441_ (_25668_, _12519_, _10377_);
  nor _76442_ (_25670_, _25668_, _25629_);
  nor _76443_ (_25671_, _25670_, _03589_);
  or _76444_ (_25672_, _25671_, _08828_);
  or _76445_ (_25673_, _25672_, _25667_);
  and _76446_ (_25674_, _12533_, _05212_);
  or _76447_ (_25675_, _25629_, _07766_);
  or _76448_ (_25676_, _25675_, _25674_);
  and _76449_ (_25677_, _05212_, _06332_);
  nor _76450_ (_25678_, _25677_, _25629_);
  and _76451_ (_25679_, _25678_, _03601_);
  nor _76452_ (_25681_, _25679_, _03780_);
  and _76453_ (_25682_, _25681_, _25676_);
  and _76454_ (_25683_, _25682_, _25673_);
  nor _76455_ (_25684_, _25683_, _25635_);
  nor _76456_ (_25685_, _25684_, _03622_);
  nor _76457_ (_25686_, _25629_, _05718_);
  not _76458_ (_25687_, _25686_);
  nor _76459_ (_25688_, _25678_, _07777_);
  and _76460_ (_25689_, _25688_, _25687_);
  nor _76461_ (_25690_, _25689_, _25685_);
  nor _76462_ (_25692_, _25690_, _03790_);
  nor _76463_ (_25693_, _25641_, _06828_);
  and _76464_ (_25694_, _25693_, _25687_);
  nor _76465_ (_25695_, _25694_, _03624_);
  not _76466_ (_25696_, _25695_);
  nor _76467_ (_25697_, _25696_, _25692_);
  nor _76468_ (_25698_, _12532_, _10377_);
  or _76469_ (_25699_, _25629_, _07795_);
  nor _76470_ (_25700_, _25699_, _25698_);
  or _76471_ (_25701_, _25700_, _03785_);
  nor _76472_ (_25703_, _25701_, _25697_);
  nor _76473_ (_25704_, _25703_, _25632_);
  nor _76474_ (_25705_, _25704_, _03815_);
  nor _76475_ (_25706_, _25649_, _04246_);
  or _76476_ (_25707_, _25706_, _03447_);
  nor _76477_ (_25708_, _25707_, _25705_);
  and _76478_ (_25709_, _12592_, _05212_);
  or _76479_ (_25710_, _25629_, _03514_);
  nor _76480_ (_25711_, _25710_, _25709_);
  nor _76481_ (_25712_, _25711_, _25708_);
  or _76482_ (_25714_, _25712_, _43004_);
  or _76483_ (_25715_, _43000_, \oc8051_golden_model_1.PCON [2]);
  and _76484_ (_25716_, _25715_, _41806_);
  and _76485_ (_43581_, _25716_, _25714_);
  not _76486_ (_25717_, \oc8051_golden_model_1.PCON [3]);
  nor _76487_ (_25718_, _05212_, _25717_);
  nor _76488_ (_25719_, _12738_, _10377_);
  nor _76489_ (_25720_, _25719_, _25718_);
  nor _76490_ (_25721_, _25720_, _07793_);
  and _76491_ (_25722_, _12739_, _05212_);
  nor _76492_ (_25724_, _25722_, _25718_);
  nor _76493_ (_25725_, _25724_, _07778_);
  and _76494_ (_25726_, _06592_, _05212_);
  or _76495_ (_25727_, _25726_, _25718_);
  and _76496_ (_25728_, _25727_, _04481_);
  and _76497_ (_25729_, _05212_, \oc8051_golden_model_1.ACC [3]);
  nor _76498_ (_25730_, _25729_, _25718_);
  nor _76499_ (_25731_, _25730_, _03737_);
  nor _76500_ (_25732_, _25730_, _09029_);
  nor _76501_ (_25733_, _04409_, _25717_);
  or _76502_ (_25734_, _25733_, _25732_);
  and _76503_ (_25735_, _25734_, _04081_);
  nor _76504_ (_25736_, _12627_, _10377_);
  nor _76505_ (_25737_, _25736_, _25718_);
  nor _76506_ (_25738_, _25737_, _04081_);
  or _76507_ (_25739_, _25738_, _25735_);
  and _76508_ (_25740_, _25739_, _03996_);
  nor _76509_ (_25741_, _10377_, _05005_);
  nor _76510_ (_25742_, _25741_, _25718_);
  nor _76511_ (_25743_, _25742_, _03996_);
  nor _76512_ (_25746_, _25743_, _25740_);
  nor _76513_ (_25747_, _25746_, _03729_);
  or _76514_ (_25748_, _25747_, _07390_);
  nor _76515_ (_25749_, _25748_, _25731_);
  and _76516_ (_25750_, _25742_, _07390_);
  or _76517_ (_25751_, _25750_, _04481_);
  nor _76518_ (_25752_, _25751_, _25749_);
  or _76519_ (_25753_, _25752_, _25728_);
  and _76520_ (_25754_, _25753_, _03589_);
  nor _76521_ (_25755_, _12718_, _10377_);
  nor _76522_ (_25757_, _25755_, _25718_);
  nor _76523_ (_25758_, _25757_, _03589_);
  or _76524_ (_25759_, _25758_, _08828_);
  or _76525_ (_25760_, _25759_, _25754_);
  and _76526_ (_25761_, _12733_, _05212_);
  or _76527_ (_25762_, _25718_, _07766_);
  or _76528_ (_25763_, _25762_, _25761_);
  and _76529_ (_25764_, _05212_, _06276_);
  nor _76530_ (_25765_, _25764_, _25718_);
  and _76531_ (_25766_, _25765_, _03601_);
  nor _76532_ (_25768_, _25766_, _03780_);
  and _76533_ (_25769_, _25768_, _25763_);
  and _76534_ (_25770_, _25769_, _25760_);
  nor _76535_ (_25771_, _25770_, _25725_);
  nor _76536_ (_25772_, _25771_, _03622_);
  nor _76537_ (_25773_, _25718_, _05567_);
  not _76538_ (_25774_, _25773_);
  nor _76539_ (_25775_, _25765_, _07777_);
  and _76540_ (_25776_, _25775_, _25774_);
  nor _76541_ (_25777_, _25776_, _25772_);
  nor _76542_ (_25779_, _25777_, _03790_);
  nor _76543_ (_25780_, _25730_, _06828_);
  and _76544_ (_25781_, _25780_, _25774_);
  or _76545_ (_25782_, _25781_, _25779_);
  and _76546_ (_25783_, _25782_, _07795_);
  nor _76547_ (_25784_, _12732_, _10377_);
  nor _76548_ (_25785_, _25784_, _25718_);
  nor _76549_ (_25786_, _25785_, _07795_);
  or _76550_ (_25787_, _25786_, _25783_);
  and _76551_ (_25788_, _25787_, _07793_);
  nor _76552_ (_25790_, _25788_, _25721_);
  nor _76553_ (_25791_, _25790_, _03815_);
  nor _76554_ (_25792_, _25737_, _04246_);
  or _76555_ (_25793_, _25792_, _03447_);
  nor _76556_ (_25794_, _25793_, _25791_);
  and _76557_ (_25795_, _12794_, _05212_);
  nor _76558_ (_25796_, _25795_, _25718_);
  and _76559_ (_25797_, _25796_, _03447_);
  nor _76560_ (_25798_, _25797_, _25794_);
  or _76561_ (_25799_, _25798_, _43004_);
  or _76562_ (_25801_, _43000_, \oc8051_golden_model_1.PCON [3]);
  and _76563_ (_25802_, _25801_, _41806_);
  and _76564_ (_43582_, _25802_, _25799_);
  not _76565_ (_25803_, \oc8051_golden_model_1.PCON [4]);
  nor _76566_ (_25804_, _05212_, _25803_);
  nor _76567_ (_25805_, _12816_, _10377_);
  nor _76568_ (_25806_, _25805_, _25804_);
  nor _76569_ (_25807_, _25806_, _07793_);
  and _76570_ (_25808_, _12817_, _05212_);
  nor _76571_ (_25809_, _25808_, _25804_);
  nor _76572_ (_25811_, _25809_, _07778_);
  and _76573_ (_25812_, _06298_, _05212_);
  nor _76574_ (_25813_, _25812_, _25804_);
  and _76575_ (_25814_, _25813_, _03601_);
  and _76576_ (_25815_, _05212_, \oc8051_golden_model_1.ACC [4]);
  nor _76577_ (_25816_, _25815_, _25804_);
  nor _76578_ (_25817_, _25816_, _03737_);
  nor _76579_ (_25818_, _25816_, _09029_);
  nor _76580_ (_25819_, _04409_, _25803_);
  or _76581_ (_25820_, _25819_, _25818_);
  and _76582_ (_25822_, _25820_, _04081_);
  nor _76583_ (_25823_, _12841_, _10377_);
  nor _76584_ (_25824_, _25823_, _25804_);
  nor _76585_ (_25825_, _25824_, _04081_);
  or _76586_ (_25826_, _25825_, _25822_);
  and _76587_ (_25827_, _25826_, _03996_);
  nor _76588_ (_25828_, _05777_, _10377_);
  nor _76589_ (_25829_, _25828_, _25804_);
  nor _76590_ (_25830_, _25829_, _03996_);
  nor _76591_ (_25831_, _25830_, _25827_);
  nor _76592_ (_25833_, _25831_, _03729_);
  or _76593_ (_25834_, _25833_, _07390_);
  nor _76594_ (_25835_, _25834_, _25817_);
  and _76595_ (_25836_, _25829_, _07390_);
  nor _76596_ (_25837_, _25836_, _25835_);
  nor _76597_ (_25838_, _25837_, _04481_);
  and _76598_ (_25839_, _06730_, _05212_);
  nor _76599_ (_25840_, _25804_, _07400_);
  not _76600_ (_25841_, _25840_);
  nor _76601_ (_25842_, _25841_, _25839_);
  or _76602_ (_25844_, _25842_, _03222_);
  nor _76603_ (_25845_, _25844_, _25838_);
  nor _76604_ (_25846_, _12933_, _10377_);
  nor _76605_ (_25847_, _25846_, _25804_);
  nor _76606_ (_25848_, _25847_, _03589_);
  or _76607_ (_25849_, _25848_, _03601_);
  nor _76608_ (_25850_, _25849_, _25845_);
  nor _76609_ (_25851_, _25850_, _25814_);
  or _76610_ (_25852_, _25851_, _03600_);
  and _76611_ (_25853_, _12821_, _05212_);
  or _76612_ (_25855_, _25853_, _25804_);
  or _76613_ (_25856_, _25855_, _07766_);
  and _76614_ (_25857_, _25856_, _07778_);
  and _76615_ (_25858_, _25857_, _25852_);
  nor _76616_ (_25859_, _25858_, _25811_);
  nor _76617_ (_25860_, _25859_, _03622_);
  nor _76618_ (_25861_, _25804_, _05825_);
  not _76619_ (_25862_, _25861_);
  nor _76620_ (_25863_, _25813_, _07777_);
  and _76621_ (_25864_, _25863_, _25862_);
  nor _76622_ (_25866_, _25864_, _25860_);
  nor _76623_ (_25867_, _25866_, _03790_);
  nor _76624_ (_25868_, _25816_, _06828_);
  and _76625_ (_25869_, _25868_, _25862_);
  or _76626_ (_25870_, _25869_, _25867_);
  and _76627_ (_25871_, _25870_, _07795_);
  nor _76628_ (_25872_, _12819_, _10377_);
  nor _76629_ (_25873_, _25872_, _25804_);
  nor _76630_ (_25874_, _25873_, _07795_);
  or _76631_ (_25875_, _25874_, _25871_);
  and _76632_ (_25877_, _25875_, _07793_);
  nor _76633_ (_25878_, _25877_, _25807_);
  nor _76634_ (_25879_, _25878_, _03815_);
  nor _76635_ (_25880_, _25824_, _04246_);
  or _76636_ (_25881_, _25880_, _03447_);
  nor _76637_ (_25882_, _25881_, _25879_);
  and _76638_ (_25883_, _13003_, _05212_);
  or _76639_ (_25884_, _25804_, _03514_);
  nor _76640_ (_25885_, _25884_, _25883_);
  nor _76641_ (_25886_, _25885_, _25882_);
  or _76642_ (_25888_, _25886_, _43004_);
  or _76643_ (_25889_, _43000_, \oc8051_golden_model_1.PCON [4]);
  and _76644_ (_25890_, _25889_, _41806_);
  and _76645_ (_43583_, _25890_, _25888_);
  not _76646_ (_25891_, \oc8051_golden_model_1.PCON [5]);
  nor _76647_ (_25892_, _05212_, _25891_);
  nor _76648_ (_25893_, _13146_, _10377_);
  nor _76649_ (_25894_, _25893_, _25892_);
  nor _76650_ (_25895_, _25894_, _07793_);
  and _76651_ (_25896_, _13147_, _05212_);
  nor _76652_ (_25898_, _25896_, _25892_);
  nor _76653_ (_25899_, _25898_, _07778_);
  and _76654_ (_25900_, _06684_, _05212_);
  or _76655_ (_25901_, _25900_, _25892_);
  and _76656_ (_25902_, _25901_, _04481_);
  and _76657_ (_25903_, _05212_, \oc8051_golden_model_1.ACC [5]);
  nor _76658_ (_25904_, _25903_, _25892_);
  nor _76659_ (_25905_, _25904_, _03737_);
  nor _76660_ (_25906_, _25904_, _09029_);
  nor _76661_ (_25907_, _04409_, _25891_);
  or _76662_ (_25909_, _25907_, _25906_);
  and _76663_ (_25910_, _25909_, _04081_);
  nor _76664_ (_25911_, _13014_, _10377_);
  nor _76665_ (_25912_, _25911_, _25892_);
  nor _76666_ (_25913_, _25912_, _04081_);
  or _76667_ (_25914_, _25913_, _25910_);
  and _76668_ (_25915_, _25914_, _03996_);
  nor _76669_ (_25916_, _05469_, _10377_);
  nor _76670_ (_25917_, _25916_, _25892_);
  nor _76671_ (_25918_, _25917_, _03996_);
  nor _76672_ (_25920_, _25918_, _25915_);
  nor _76673_ (_25921_, _25920_, _03729_);
  or _76674_ (_25922_, _25921_, _07390_);
  nor _76675_ (_25923_, _25922_, _25905_);
  and _76676_ (_25924_, _25917_, _07390_);
  or _76677_ (_25925_, _25924_, _04481_);
  nor _76678_ (_25926_, _25925_, _25923_);
  or _76679_ (_25927_, _25926_, _25902_);
  and _76680_ (_25928_, _25927_, _03589_);
  nor _76681_ (_25929_, _13127_, _10377_);
  nor _76682_ (_25931_, _25929_, _25892_);
  nor _76683_ (_25932_, _25931_, _03589_);
  or _76684_ (_25933_, _25932_, _08828_);
  or _76685_ (_25934_, _25933_, _25928_);
  and _76686_ (_25935_, _13141_, _05212_);
  or _76687_ (_25936_, _25892_, _07766_);
  or _76688_ (_25937_, _25936_, _25935_);
  and _76689_ (_25938_, _06306_, _05212_);
  nor _76690_ (_25939_, _25938_, _25892_);
  and _76691_ (_25940_, _25939_, _03601_);
  nor _76692_ (_25942_, _25940_, _03780_);
  and _76693_ (_25943_, _25942_, _25937_);
  and _76694_ (_25944_, _25943_, _25934_);
  nor _76695_ (_25945_, _25944_, _25899_);
  nor _76696_ (_25946_, _25945_, _03622_);
  nor _76697_ (_25947_, _25892_, _05518_);
  not _76698_ (_25948_, _25947_);
  nor _76699_ (_25949_, _25939_, _07777_);
  and _76700_ (_25950_, _25949_, _25948_);
  nor _76701_ (_25951_, _25950_, _25946_);
  nor _76702_ (_25953_, _25951_, _03790_);
  nor _76703_ (_25954_, _25904_, _06828_);
  and _76704_ (_25955_, _25954_, _25948_);
  nor _76705_ (_25956_, _25955_, _03624_);
  not _76706_ (_25957_, _25956_);
  nor _76707_ (_25958_, _25957_, _25953_);
  nor _76708_ (_25959_, _13140_, _10377_);
  or _76709_ (_25960_, _25892_, _07795_);
  nor _76710_ (_25961_, _25960_, _25959_);
  or _76711_ (_25962_, _25961_, _03785_);
  nor _76712_ (_25964_, _25962_, _25958_);
  nor _76713_ (_25965_, _25964_, _25895_);
  nor _76714_ (_25966_, _25965_, _03815_);
  nor _76715_ (_25967_, _25912_, _04246_);
  or _76716_ (_25968_, _25967_, _03447_);
  nor _76717_ (_25969_, _25968_, _25966_);
  and _76718_ (_25970_, _13199_, _05212_);
  or _76719_ (_25971_, _25892_, _03514_);
  nor _76720_ (_25972_, _25971_, _25970_);
  nor _76721_ (_25973_, _25972_, _25969_);
  or _76722_ (_25975_, _25973_, _43004_);
  or _76723_ (_25976_, _43000_, \oc8051_golden_model_1.PCON [5]);
  and _76724_ (_25977_, _25976_, _41806_);
  and _76725_ (_43584_, _25977_, _25975_);
  not _76726_ (_25978_, \oc8051_golden_model_1.PCON [6]);
  nor _76727_ (_25979_, _05212_, _25978_);
  nor _76728_ (_25980_, _13352_, _10377_);
  nor _76729_ (_25981_, _25980_, _25979_);
  nor _76730_ (_25982_, _25981_, _07793_);
  and _76731_ (_25983_, _13353_, _05212_);
  nor _76732_ (_25985_, _25983_, _25979_);
  nor _76733_ (_25986_, _25985_, _07778_);
  and _76734_ (_25987_, _06455_, _05212_);
  or _76735_ (_25988_, _25987_, _25979_);
  and _76736_ (_25989_, _25988_, _04481_);
  and _76737_ (_25990_, _05212_, \oc8051_golden_model_1.ACC [6]);
  nor _76738_ (_25991_, _25990_, _25979_);
  nor _76739_ (_25992_, _25991_, _03737_);
  nor _76740_ (_25993_, _25991_, _09029_);
  nor _76741_ (_25994_, _04409_, _25978_);
  or _76742_ (_25996_, _25994_, _25993_);
  and _76743_ (_25997_, _25996_, _04081_);
  nor _76744_ (_25998_, _13242_, _10377_);
  nor _76745_ (_25999_, _25998_, _25979_);
  nor _76746_ (_26000_, _25999_, _04081_);
  or _76747_ (_26001_, _26000_, _25997_);
  and _76748_ (_26002_, _26001_, _03996_);
  nor _76749_ (_26003_, _05363_, _10377_);
  nor _76750_ (_26004_, _26003_, _25979_);
  nor _76751_ (_26005_, _26004_, _03996_);
  nor _76752_ (_26007_, _26005_, _26002_);
  nor _76753_ (_26008_, _26007_, _03729_);
  or _76754_ (_26009_, _26008_, _07390_);
  nor _76755_ (_26010_, _26009_, _25992_);
  and _76756_ (_26011_, _26004_, _07390_);
  or _76757_ (_26012_, _26011_, _04481_);
  nor _76758_ (_26013_, _26012_, _26010_);
  or _76759_ (_26014_, _26013_, _25989_);
  and _76760_ (_26015_, _26014_, _03589_);
  nor _76761_ (_26016_, _13332_, _10377_);
  nor _76762_ (_26018_, _26016_, _25979_);
  nor _76763_ (_26019_, _26018_, _03589_);
  or _76764_ (_26020_, _26019_, _08828_);
  or _76765_ (_26021_, _26020_, _26015_);
  and _76766_ (_26022_, _13347_, _05212_);
  or _76767_ (_26023_, _25979_, _07766_);
  or _76768_ (_26024_, _26023_, _26022_);
  and _76769_ (_26025_, _13339_, _05212_);
  nor _76770_ (_26026_, _26025_, _25979_);
  and _76771_ (_26027_, _26026_, _03601_);
  nor _76772_ (_26029_, _26027_, _03780_);
  and _76773_ (_26030_, _26029_, _26024_);
  and _76774_ (_26031_, _26030_, _26021_);
  nor _76775_ (_26032_, _26031_, _25986_);
  nor _76776_ (_26033_, _26032_, _03622_);
  nor _76777_ (_26034_, _25979_, _05412_);
  not _76778_ (_26035_, _26034_);
  nor _76779_ (_26036_, _26026_, _07777_);
  and _76780_ (_26037_, _26036_, _26035_);
  nor _76781_ (_26038_, _26037_, _26033_);
  nor _76782_ (_26040_, _26038_, _03790_);
  nor _76783_ (_26041_, _25991_, _06828_);
  and _76784_ (_26042_, _26041_, _26035_);
  or _76785_ (_26043_, _26042_, _26040_);
  and _76786_ (_26044_, _26043_, _07795_);
  nor _76787_ (_26045_, _13346_, _10377_);
  nor _76788_ (_26046_, _26045_, _25979_);
  nor _76789_ (_26047_, _26046_, _07795_);
  or _76790_ (_26048_, _26047_, _26044_);
  and _76791_ (_26049_, _26048_, _07793_);
  nor _76792_ (_26051_, _26049_, _25982_);
  nor _76793_ (_26052_, _26051_, _03815_);
  nor _76794_ (_26053_, _25999_, _04246_);
  or _76795_ (_26054_, _26053_, _03447_);
  nor _76796_ (_26055_, _26054_, _26052_);
  and _76797_ (_26056_, _13402_, _05212_);
  or _76798_ (_26057_, _25979_, _03514_);
  nor _76799_ (_26058_, _26057_, _26056_);
  nor _76800_ (_26059_, _26058_, _26055_);
  or _76801_ (_26060_, _26059_, _43004_);
  or _76802_ (_26062_, _43000_, \oc8051_golden_model_1.PCON [6]);
  and _76803_ (_26063_, _26062_, _41806_);
  and _76804_ (_43585_, _26063_, _26060_);
  not _76805_ (_26064_, \oc8051_golden_model_1.SBUF [0]);
  nor _76806_ (_26065_, _05221_, _26064_);
  nor _76807_ (_26066_, _05666_, _10458_);
  nor _76808_ (_26067_, _26066_, _26065_);
  and _76809_ (_26068_, _26067_, _17166_);
  and _76810_ (_26069_, _05221_, \oc8051_golden_model_1.ACC [0]);
  nor _76811_ (_26070_, _26069_, _26065_);
  nor _76812_ (_26072_, _26070_, _03737_);
  nor _76813_ (_26073_, _26072_, _07390_);
  nor _76814_ (_26074_, _26067_, _04081_);
  nor _76815_ (_26075_, _04409_, _26064_);
  nor _76816_ (_26076_, _26070_, _09029_);
  nor _76817_ (_26077_, _26076_, _26075_);
  nor _76818_ (_26078_, _26077_, _03610_);
  or _76819_ (_26079_, _26078_, _03723_);
  nor _76820_ (_26080_, _26079_, _26074_);
  or _76821_ (_26081_, _26080_, _03729_);
  and _76822_ (_26082_, _26081_, _26073_);
  and _76823_ (_26083_, _05221_, _04620_);
  or _76824_ (_26084_, _26065_, _25480_);
  nor _76825_ (_26085_, _26084_, _26083_);
  nor _76826_ (_26086_, _26085_, _26082_);
  nor _76827_ (_26087_, _26086_, _04481_);
  and _76828_ (_26088_, _06546_, _05221_);
  nor _76829_ (_26089_, _26065_, _07400_);
  not _76830_ (_26090_, _26089_);
  nor _76831_ (_26091_, _26090_, _26088_);
  nor _76832_ (_26094_, _26091_, _26087_);
  nor _76833_ (_26095_, _26094_, _03222_);
  nor _76834_ (_26096_, _12109_, _10458_);
  or _76835_ (_26097_, _26065_, _03589_);
  nor _76836_ (_26098_, _26097_, _26096_);
  or _76837_ (_26099_, _26098_, _03601_);
  nor _76838_ (_26100_, _26099_, _26095_);
  and _76839_ (_26101_, _05221_, _06274_);
  nor _76840_ (_26102_, _26101_, _26065_);
  nand _76841_ (_26103_, _26102_, _07766_);
  and _76842_ (_26105_, _26103_, _08828_);
  nor _76843_ (_26106_, _26105_, _26100_);
  and _76844_ (_26107_, _12124_, _05221_);
  nor _76845_ (_26108_, _26107_, _26065_);
  and _76846_ (_26109_, _26108_, _03600_);
  nor _76847_ (_26110_, _26109_, _26106_);
  nor _76848_ (_26111_, _26110_, _03780_);
  and _76849_ (_26112_, _12128_, _05221_);
  or _76850_ (_26113_, _26065_, _07778_);
  nor _76851_ (_26114_, _26113_, _26112_);
  or _76852_ (_26116_, _26114_, _03622_);
  nor _76853_ (_26117_, _26116_, _26111_);
  or _76854_ (_26118_, _26102_, _07777_);
  nor _76855_ (_26119_, _26118_, _26066_);
  nor _76856_ (_26120_, _26119_, _26117_);
  nor _76857_ (_26121_, _26120_, _03790_);
  nor _76858_ (_26122_, _26065_, _05666_);
  or _76859_ (_26123_, _26122_, _06828_);
  nor _76860_ (_26124_, _26123_, _26070_);
  or _76861_ (_26125_, _26124_, _26121_);
  and _76862_ (_26127_, _26125_, _07795_);
  nor _76863_ (_26128_, _12122_, _10458_);
  nor _76864_ (_26129_, _26128_, _26065_);
  nor _76865_ (_26130_, _26129_, _07795_);
  or _76866_ (_26131_, _26130_, _26127_);
  and _76867_ (_26132_, _26131_, _07793_);
  nor _76868_ (_26133_, _12003_, _10458_);
  nor _76869_ (_26134_, _26133_, _26065_);
  nor _76870_ (_26135_, _26134_, _07793_);
  nor _76871_ (_26136_, _26135_, _17166_);
  not _76872_ (_26138_, _26136_);
  nor _76873_ (_26139_, _26138_, _26132_);
  nor _76874_ (_26140_, _26139_, _26068_);
  or _76875_ (_26141_, _26140_, _43004_);
  or _76876_ (_26142_, _43000_, \oc8051_golden_model_1.SBUF [0]);
  and _76877_ (_26143_, _26142_, _41806_);
  and _76878_ (_43588_, _26143_, _26141_);
  and _76879_ (_26144_, _06501_, _05221_);
  not _76880_ (_26145_, \oc8051_golden_model_1.SBUF [1]);
  nor _76881_ (_26146_, _05221_, _26145_);
  nor _76882_ (_26148_, _26146_, _07400_);
  not _76883_ (_26149_, _26148_);
  nor _76884_ (_26150_, _26149_, _26144_);
  not _76885_ (_26151_, _26150_);
  and _76886_ (_26152_, _05221_, _06764_);
  nor _76887_ (_26153_, _26152_, _26146_);
  and _76888_ (_26154_, _26153_, _07390_);
  nor _76889_ (_26155_, _05221_, \oc8051_golden_model_1.SBUF [1]);
  and _76890_ (_26156_, _05221_, _03274_);
  nor _76891_ (_26157_, _26156_, _26155_);
  and _76892_ (_26159_, _26157_, _03729_);
  and _76893_ (_26160_, _26157_, _04409_);
  nor _76894_ (_26161_, _04409_, _26145_);
  or _76895_ (_26162_, _26161_, _26160_);
  and _76896_ (_26163_, _26162_, _04081_);
  and _76897_ (_26164_, _12213_, _05221_);
  nor _76898_ (_26165_, _26164_, _26155_);
  and _76899_ (_26166_, _26165_, _03610_);
  or _76900_ (_26167_, _26166_, _26163_);
  and _76901_ (_26168_, _26167_, _03996_);
  nor _76902_ (_26170_, _26153_, _03996_);
  nor _76903_ (_26171_, _26170_, _26168_);
  nor _76904_ (_26172_, _26171_, _03729_);
  or _76905_ (_26173_, _26172_, _07390_);
  nor _76906_ (_26174_, _26173_, _26159_);
  nor _76907_ (_26175_, _26174_, _26154_);
  nor _76908_ (_26176_, _26175_, _04481_);
  nor _76909_ (_26177_, _26176_, _03222_);
  and _76910_ (_26178_, _26177_, _26151_);
  not _76911_ (_26179_, _26155_);
  and _76912_ (_26181_, _12313_, _05221_);
  nor _76913_ (_26182_, _26181_, _03589_);
  and _76914_ (_26183_, _26182_, _26179_);
  nor _76915_ (_26184_, _26183_, _26178_);
  nor _76916_ (_26185_, _26184_, _08828_);
  nor _76917_ (_26186_, _12327_, _10458_);
  nor _76918_ (_26187_, _26186_, _07766_);
  and _76919_ (_26188_, _05221_, _04303_);
  nor _76920_ (_26189_, _26188_, _05886_);
  nor _76921_ (_26190_, _26189_, _26187_);
  nor _76922_ (_26191_, _26190_, _26155_);
  nor _76923_ (_26192_, _26191_, _26185_);
  nor _76924_ (_26193_, _26192_, _03780_);
  nor _76925_ (_26194_, _12333_, _10458_);
  nor _76926_ (_26195_, _26194_, _07778_);
  and _76927_ (_26196_, _26195_, _26179_);
  nor _76928_ (_26197_, _26196_, _26193_);
  nor _76929_ (_26198_, _26197_, _03622_);
  nor _76930_ (_26199_, _12207_, _10458_);
  nor _76931_ (_26200_, _26199_, _07777_);
  and _76932_ (_26203_, _26200_, _26179_);
  nor _76933_ (_26204_, _26203_, _26198_);
  nor _76934_ (_26205_, _26204_, _03790_);
  nor _76935_ (_26206_, _26146_, _05618_);
  nor _76936_ (_26207_, _26206_, _06828_);
  and _76937_ (_26208_, _26207_, _26157_);
  nor _76938_ (_26209_, _26208_, _26205_);
  or _76939_ (_26210_, _26209_, _18499_);
  and _76940_ (_26211_, _26188_, _05617_);
  nor _76941_ (_26212_, _26211_, _07795_);
  and _76942_ (_26214_, _26212_, _26179_);
  nand _76943_ (_26215_, _26156_, _05617_);
  nor _76944_ (_26216_, _26155_, _07793_);
  and _76945_ (_26217_, _26216_, _26215_);
  or _76946_ (_26218_, _26217_, _03815_);
  nor _76947_ (_26219_, _26218_, _26214_);
  and _76948_ (_26220_, _26219_, _26210_);
  nor _76949_ (_26221_, _26165_, _04246_);
  nor _76950_ (_26222_, _26221_, _26220_);
  and _76951_ (_26223_, _26222_, _03514_);
  nor _76952_ (_26225_, _26164_, _26146_);
  nor _76953_ (_26226_, _26225_, _03514_);
  or _76954_ (_26227_, _26226_, _26223_);
  or _76955_ (_26228_, _26227_, _43004_);
  or _76956_ (_26229_, _43000_, \oc8051_golden_model_1.SBUF [1]);
  and _76957_ (_26230_, _26229_, _41806_);
  and _76958_ (_43589_, _26230_, _26228_);
  not _76959_ (_26231_, \oc8051_golden_model_1.SBUF [2]);
  nor _76960_ (_26232_, _05221_, _26231_);
  nor _76961_ (_26233_, _12538_, _10458_);
  nor _76962_ (_26235_, _26233_, _26232_);
  nor _76963_ (_26236_, _26235_, _07793_);
  and _76964_ (_26237_, _12539_, _05221_);
  nor _76965_ (_26238_, _26237_, _26232_);
  nor _76966_ (_26239_, _26238_, _07778_);
  nor _76967_ (_26240_, _10458_, _04875_);
  nor _76968_ (_26241_, _26240_, _26232_);
  and _76969_ (_26242_, _26241_, _07390_);
  and _76970_ (_26243_, _05221_, \oc8051_golden_model_1.ACC [2]);
  nor _76971_ (_26244_, _26243_, _26232_);
  nor _76972_ (_26246_, _26244_, _03737_);
  nor _76973_ (_26247_, _26244_, _09029_);
  nor _76974_ (_26248_, _04409_, _26231_);
  or _76975_ (_26249_, _26248_, _26247_);
  and _76976_ (_26250_, _26249_, _04081_);
  nor _76977_ (_26251_, _12416_, _10458_);
  nor _76978_ (_26252_, _26251_, _26232_);
  nor _76979_ (_26253_, _26252_, _04081_);
  or _76980_ (_26254_, _26253_, _26250_);
  and _76981_ (_26255_, _26254_, _03996_);
  nor _76982_ (_26257_, _26241_, _03996_);
  nor _76983_ (_26258_, _26257_, _26255_);
  nor _76984_ (_26259_, _26258_, _03729_);
  or _76985_ (_26260_, _26259_, _07390_);
  nor _76986_ (_26261_, _26260_, _26246_);
  nor _76987_ (_26262_, _26261_, _26242_);
  nor _76988_ (_26263_, _26262_, _04481_);
  and _76989_ (_26264_, _06637_, _05221_);
  nor _76990_ (_26265_, _26232_, _07400_);
  not _76991_ (_26266_, _26265_);
  nor _76992_ (_26268_, _26266_, _26264_);
  nor _76993_ (_26269_, _26268_, _03222_);
  not _76994_ (_26270_, _26269_);
  nor _76995_ (_26271_, _26270_, _26263_);
  nor _76996_ (_26272_, _12519_, _10458_);
  nor _76997_ (_26273_, _26272_, _26232_);
  nor _76998_ (_26274_, _26273_, _03589_);
  or _76999_ (_26275_, _26274_, _08828_);
  or _77000_ (_26276_, _26275_, _26271_);
  and _77001_ (_26277_, _12533_, _05221_);
  or _77002_ (_26279_, _26232_, _07766_);
  or _77003_ (_26280_, _26279_, _26277_);
  and _77004_ (_26281_, _05221_, _06332_);
  nor _77005_ (_26282_, _26281_, _26232_);
  and _77006_ (_26283_, _26282_, _03601_);
  nor _77007_ (_26284_, _26283_, _03780_);
  and _77008_ (_26285_, _26284_, _26280_);
  and _77009_ (_26286_, _26285_, _26276_);
  nor _77010_ (_26287_, _26286_, _26239_);
  nor _77011_ (_26288_, _26287_, _03622_);
  nor _77012_ (_26290_, _26232_, _05718_);
  not _77013_ (_26291_, _26290_);
  nor _77014_ (_26292_, _26282_, _07777_);
  and _77015_ (_26293_, _26292_, _26291_);
  nor _77016_ (_26294_, _26293_, _26288_);
  nor _77017_ (_26295_, _26294_, _03790_);
  nor _77018_ (_26296_, _26244_, _06828_);
  and _77019_ (_26297_, _26296_, _26291_);
  nor _77020_ (_26298_, _26297_, _03624_);
  not _77021_ (_26299_, _26298_);
  nor _77022_ (_26301_, _26299_, _26295_);
  nor _77023_ (_26302_, _12532_, _10458_);
  or _77024_ (_26303_, _26232_, _07795_);
  nor _77025_ (_26304_, _26303_, _26302_);
  or _77026_ (_26305_, _26304_, _03785_);
  nor _77027_ (_26306_, _26305_, _26301_);
  nor _77028_ (_26307_, _26306_, _26236_);
  nor _77029_ (_26308_, _26307_, _03815_);
  nor _77030_ (_26309_, _26252_, _04246_);
  or _77031_ (_26310_, _26309_, _03447_);
  nor _77032_ (_26312_, _26310_, _26308_);
  and _77033_ (_26313_, _12592_, _05221_);
  or _77034_ (_26314_, _26232_, _03514_);
  nor _77035_ (_26315_, _26314_, _26313_);
  nor _77036_ (_26316_, _26315_, _26312_);
  or _77037_ (_26317_, _26316_, _43004_);
  or _77038_ (_26318_, _43000_, \oc8051_golden_model_1.SBUF [2]);
  and _77039_ (_26319_, _26318_, _41806_);
  and _77040_ (_43590_, _26319_, _26317_);
  not _77041_ (_26320_, \oc8051_golden_model_1.SBUF [3]);
  nor _77042_ (_26322_, _05221_, _26320_);
  nor _77043_ (_26323_, _12738_, _10458_);
  nor _77044_ (_26324_, _26323_, _26322_);
  nor _77045_ (_26325_, _26324_, _07793_);
  and _77046_ (_26326_, _12739_, _05221_);
  nor _77047_ (_26327_, _26326_, _26322_);
  nor _77048_ (_26328_, _26327_, _07778_);
  and _77049_ (_26329_, _06592_, _05221_);
  or _77050_ (_26330_, _26329_, _26322_);
  and _77051_ (_26331_, _26330_, _04481_);
  and _77052_ (_26333_, _05221_, \oc8051_golden_model_1.ACC [3]);
  nor _77053_ (_26334_, _26333_, _26322_);
  nor _77054_ (_26335_, _26334_, _03737_);
  nor _77055_ (_26336_, _26334_, _09029_);
  nor _77056_ (_26337_, _04409_, _26320_);
  or _77057_ (_26338_, _26337_, _26336_);
  and _77058_ (_26339_, _26338_, _04081_);
  nor _77059_ (_26340_, _12627_, _10458_);
  nor _77060_ (_26341_, _26340_, _26322_);
  nor _77061_ (_26342_, _26341_, _04081_);
  or _77062_ (_26344_, _26342_, _26339_);
  and _77063_ (_26345_, _26344_, _03996_);
  nor _77064_ (_26346_, _10458_, _05005_);
  nor _77065_ (_26347_, _26346_, _26322_);
  nor _77066_ (_26348_, _26347_, _03996_);
  nor _77067_ (_26349_, _26348_, _26345_);
  nor _77068_ (_26350_, _26349_, _03729_);
  or _77069_ (_26351_, _26350_, _07390_);
  nor _77070_ (_26352_, _26351_, _26335_);
  and _77071_ (_26353_, _26347_, _07390_);
  or _77072_ (_26355_, _26353_, _04481_);
  nor _77073_ (_26356_, _26355_, _26352_);
  or _77074_ (_26357_, _26356_, _26331_);
  and _77075_ (_26358_, _26357_, _03589_);
  nor _77076_ (_26359_, _12718_, _10458_);
  nor _77077_ (_26360_, _26359_, _26322_);
  nor _77078_ (_26361_, _26360_, _03589_);
  or _77079_ (_26362_, _26361_, _08828_);
  or _77080_ (_26363_, _26362_, _26358_);
  and _77081_ (_26364_, _12733_, _05221_);
  or _77082_ (_26366_, _26322_, _07766_);
  or _77083_ (_26367_, _26366_, _26364_);
  and _77084_ (_26368_, _05221_, _06276_);
  nor _77085_ (_26369_, _26368_, _26322_);
  and _77086_ (_26370_, _26369_, _03601_);
  nor _77087_ (_26371_, _26370_, _03780_);
  and _77088_ (_26372_, _26371_, _26367_);
  and _77089_ (_26373_, _26372_, _26363_);
  nor _77090_ (_26374_, _26373_, _26328_);
  nor _77091_ (_26375_, _26374_, _03622_);
  nor _77092_ (_26377_, _26322_, _05567_);
  not _77093_ (_26378_, _26377_);
  nor _77094_ (_26379_, _26369_, _07777_);
  and _77095_ (_26380_, _26379_, _26378_);
  nor _77096_ (_26381_, _26380_, _26375_);
  nor _77097_ (_26382_, _26381_, _03790_);
  nor _77098_ (_26383_, _26334_, _06828_);
  and _77099_ (_26384_, _26383_, _26378_);
  nor _77100_ (_26385_, _26384_, _03624_);
  not _77101_ (_26386_, _26385_);
  nor _77102_ (_26388_, _26386_, _26382_);
  nor _77103_ (_26389_, _12732_, _10458_);
  or _77104_ (_26390_, _26322_, _07795_);
  nor _77105_ (_26391_, _26390_, _26389_);
  or _77106_ (_26392_, _26391_, _03785_);
  nor _77107_ (_26393_, _26392_, _26388_);
  nor _77108_ (_26394_, _26393_, _26325_);
  nor _77109_ (_26395_, _26394_, _03815_);
  nor _77110_ (_26396_, _26341_, _04246_);
  or _77111_ (_26397_, _26396_, _03447_);
  nor _77112_ (_26399_, _26397_, _26395_);
  and _77113_ (_26400_, _12794_, _05221_);
  or _77114_ (_26401_, _26322_, _03514_);
  nor _77115_ (_26402_, _26401_, _26400_);
  nor _77116_ (_26403_, _26402_, _26399_);
  or _77117_ (_26404_, _26403_, _43004_);
  or _77118_ (_26405_, _43000_, \oc8051_golden_model_1.SBUF [3]);
  and _77119_ (_26406_, _26405_, _41806_);
  and _77120_ (_43591_, _26406_, _26404_);
  not _77121_ (_26407_, \oc8051_golden_model_1.SBUF [4]);
  nor _77122_ (_26409_, _05221_, _26407_);
  nor _77123_ (_26410_, _12816_, _10458_);
  nor _77124_ (_26411_, _26410_, _26409_);
  nor _77125_ (_26412_, _26411_, _07793_);
  and _77126_ (_26413_, _12817_, _05221_);
  nor _77127_ (_26414_, _26413_, _26409_);
  nor _77128_ (_26415_, _26414_, _07778_);
  and _77129_ (_26416_, _06298_, _05221_);
  nor _77130_ (_26417_, _26416_, _26409_);
  and _77131_ (_26418_, _26417_, _03601_);
  nor _77132_ (_26420_, _05777_, _10458_);
  nor _77133_ (_26421_, _26420_, _26409_);
  and _77134_ (_26422_, _26421_, _07390_);
  and _77135_ (_26423_, _05221_, \oc8051_golden_model_1.ACC [4]);
  nor _77136_ (_26424_, _26423_, _26409_);
  nor _77137_ (_26425_, _26424_, _03737_);
  nor _77138_ (_26426_, _26424_, _09029_);
  nor _77139_ (_26427_, _04409_, _26407_);
  or _77140_ (_26428_, _26427_, _26426_);
  and _77141_ (_26429_, _26428_, _04081_);
  nor _77142_ (_26431_, _12841_, _10458_);
  nor _77143_ (_26432_, _26431_, _26409_);
  nor _77144_ (_26433_, _26432_, _04081_);
  or _77145_ (_26434_, _26433_, _26429_);
  and _77146_ (_26435_, _26434_, _03996_);
  nor _77147_ (_26436_, _26421_, _03996_);
  nor _77148_ (_26437_, _26436_, _26435_);
  nor _77149_ (_26438_, _26437_, _03729_);
  or _77150_ (_26439_, _26438_, _07390_);
  nor _77151_ (_26440_, _26439_, _26425_);
  nor _77152_ (_26442_, _26440_, _26422_);
  nor _77153_ (_26443_, _26442_, _04481_);
  and _77154_ (_26444_, _06730_, _05221_);
  nor _77155_ (_26445_, _26409_, _07400_);
  not _77156_ (_26446_, _26445_);
  nor _77157_ (_26447_, _26446_, _26444_);
  or _77158_ (_26448_, _26447_, _03222_);
  nor _77159_ (_26449_, _26448_, _26443_);
  nor _77160_ (_26450_, _12933_, _10458_);
  nor _77161_ (_26451_, _26450_, _26409_);
  nor _77162_ (_26453_, _26451_, _03589_);
  or _77163_ (_26454_, _26453_, _03601_);
  nor _77164_ (_26455_, _26454_, _26449_);
  nor _77165_ (_26456_, _26455_, _26418_);
  or _77166_ (_26457_, _26456_, _03600_);
  and _77167_ (_26458_, _12821_, _05221_);
  or _77168_ (_26459_, _26458_, _26409_);
  or _77169_ (_26460_, _26459_, _07766_);
  and _77170_ (_26461_, _26460_, _07778_);
  and _77171_ (_26462_, _26461_, _26457_);
  nor _77172_ (_26464_, _26462_, _26415_);
  nor _77173_ (_26465_, _26464_, _03622_);
  nor _77174_ (_26466_, _26409_, _05825_);
  not _77175_ (_26467_, _26466_);
  nor _77176_ (_26468_, _26417_, _07777_);
  and _77177_ (_26469_, _26468_, _26467_);
  nor _77178_ (_26470_, _26469_, _26465_);
  nor _77179_ (_26471_, _26470_, _03790_);
  nor _77180_ (_26472_, _26424_, _06828_);
  and _77181_ (_26473_, _26472_, _26467_);
  nor _77182_ (_26475_, _26473_, _03624_);
  not _77183_ (_26476_, _26475_);
  nor _77184_ (_26477_, _26476_, _26471_);
  nor _77185_ (_26478_, _12819_, _10458_);
  or _77186_ (_26479_, _26409_, _07795_);
  nor _77187_ (_26480_, _26479_, _26478_);
  or _77188_ (_26481_, _26480_, _03785_);
  nor _77189_ (_26482_, _26481_, _26477_);
  nor _77190_ (_26483_, _26482_, _26412_);
  nor _77191_ (_26484_, _26483_, _03815_);
  nor _77192_ (_26486_, _26432_, _04246_);
  or _77193_ (_26487_, _26486_, _03447_);
  nor _77194_ (_26488_, _26487_, _26484_);
  and _77195_ (_26489_, _13003_, _05221_);
  or _77196_ (_26490_, _26409_, _03514_);
  nor _77197_ (_26491_, _26490_, _26489_);
  nor _77198_ (_26492_, _26491_, _26488_);
  or _77199_ (_26493_, _26492_, _43004_);
  or _77200_ (_26494_, _43000_, \oc8051_golden_model_1.SBUF [4]);
  and _77201_ (_26495_, _26494_, _41806_);
  and _77202_ (_43592_, _26495_, _26493_);
  not _77203_ (_26497_, \oc8051_golden_model_1.SBUF [5]);
  nor _77204_ (_26498_, _05221_, _26497_);
  nor _77205_ (_26499_, _13146_, _10458_);
  nor _77206_ (_26500_, _26499_, _26498_);
  nor _77207_ (_26501_, _26500_, _07793_);
  and _77208_ (_26502_, _13147_, _05221_);
  nor _77209_ (_26503_, _26502_, _26498_);
  nor _77210_ (_26504_, _26503_, _07778_);
  and _77211_ (_26505_, _06684_, _05221_);
  or _77212_ (_26507_, _26505_, _26498_);
  and _77213_ (_26508_, _26507_, _04481_);
  and _77214_ (_26509_, _05221_, \oc8051_golden_model_1.ACC [5]);
  nor _77215_ (_26510_, _26509_, _26498_);
  nor _77216_ (_26511_, _26510_, _03737_);
  nor _77217_ (_26512_, _26510_, _09029_);
  nor _77218_ (_26513_, _04409_, _26497_);
  or _77219_ (_26514_, _26513_, _26512_);
  and _77220_ (_26515_, _26514_, _04081_);
  nor _77221_ (_26516_, _13014_, _10458_);
  nor _77222_ (_26518_, _26516_, _26498_);
  nor _77223_ (_26519_, _26518_, _04081_);
  or _77224_ (_26520_, _26519_, _26515_);
  and _77225_ (_26521_, _26520_, _03996_);
  nor _77226_ (_26522_, _05469_, _10458_);
  nor _77227_ (_26523_, _26522_, _26498_);
  nor _77228_ (_26524_, _26523_, _03996_);
  nor _77229_ (_26525_, _26524_, _26521_);
  nor _77230_ (_26526_, _26525_, _03729_);
  or _77231_ (_26527_, _26526_, _07390_);
  nor _77232_ (_26529_, _26527_, _26511_);
  and _77233_ (_26530_, _26523_, _07390_);
  or _77234_ (_26531_, _26530_, _04481_);
  nor _77235_ (_26532_, _26531_, _26529_);
  or _77236_ (_26533_, _26532_, _26508_);
  and _77237_ (_26534_, _26533_, _03589_);
  nor _77238_ (_26535_, _13127_, _10458_);
  nor _77239_ (_26536_, _26535_, _26498_);
  nor _77240_ (_26537_, _26536_, _03589_);
  or _77241_ (_26538_, _26537_, _08828_);
  or _77242_ (_26540_, _26538_, _26534_);
  and _77243_ (_26541_, _13141_, _05221_);
  or _77244_ (_26542_, _26498_, _07766_);
  or _77245_ (_26543_, _26542_, _26541_);
  and _77246_ (_26544_, _06306_, _05221_);
  nor _77247_ (_26545_, _26544_, _26498_);
  and _77248_ (_26546_, _26545_, _03601_);
  nor _77249_ (_26547_, _26546_, _03780_);
  and _77250_ (_26548_, _26547_, _26543_);
  and _77251_ (_26549_, _26548_, _26540_);
  nor _77252_ (_26551_, _26549_, _26504_);
  nor _77253_ (_26552_, _26551_, _03622_);
  nor _77254_ (_26553_, _26498_, _05518_);
  not _77255_ (_26554_, _26553_);
  nor _77256_ (_26555_, _26545_, _07777_);
  and _77257_ (_26556_, _26555_, _26554_);
  nor _77258_ (_26557_, _26556_, _26552_);
  nor _77259_ (_26558_, _26557_, _03790_);
  nor _77260_ (_26559_, _26510_, _06828_);
  and _77261_ (_26560_, _26559_, _26554_);
  nor _77262_ (_26562_, _26560_, _03624_);
  not _77263_ (_26563_, _26562_);
  nor _77264_ (_26564_, _26563_, _26558_);
  nor _77265_ (_26565_, _13140_, _10458_);
  or _77266_ (_26566_, _26498_, _07795_);
  nor _77267_ (_26567_, _26566_, _26565_);
  or _77268_ (_26568_, _26567_, _03785_);
  nor _77269_ (_26569_, _26568_, _26564_);
  nor _77270_ (_26570_, _26569_, _26501_);
  nor _77271_ (_26571_, _26570_, _03815_);
  nor _77272_ (_26573_, _26518_, _04246_);
  or _77273_ (_26574_, _26573_, _03447_);
  nor _77274_ (_26575_, _26574_, _26571_);
  and _77275_ (_26576_, _13199_, _05221_);
  or _77276_ (_26577_, _26498_, _03514_);
  nor _77277_ (_26578_, _26577_, _26576_);
  nor _77278_ (_26579_, _26578_, _26575_);
  or _77279_ (_26580_, _26579_, _43004_);
  or _77280_ (_26581_, _43000_, \oc8051_golden_model_1.SBUF [5]);
  and _77281_ (_26582_, _26581_, _41806_);
  and _77282_ (_43594_, _26582_, _26580_);
  not _77283_ (_26584_, \oc8051_golden_model_1.SBUF [6]);
  nor _77284_ (_26585_, _05221_, _26584_);
  nor _77285_ (_26586_, _13352_, _10458_);
  nor _77286_ (_26587_, _26586_, _26585_);
  nor _77287_ (_26588_, _26587_, _07793_);
  and _77288_ (_26589_, _13353_, _05221_);
  nor _77289_ (_26590_, _26589_, _26585_);
  nor _77290_ (_26591_, _26590_, _07778_);
  and _77291_ (_26592_, _06455_, _05221_);
  or _77292_ (_26594_, _26592_, _26585_);
  and _77293_ (_26595_, _26594_, _04481_);
  and _77294_ (_26596_, _05221_, \oc8051_golden_model_1.ACC [6]);
  nor _77295_ (_26597_, _26596_, _26585_);
  nor _77296_ (_26598_, _26597_, _03737_);
  nor _77297_ (_26599_, _26597_, _09029_);
  nor _77298_ (_26600_, _04409_, _26584_);
  or _77299_ (_26601_, _26600_, _26599_);
  and _77300_ (_26602_, _26601_, _04081_);
  nor _77301_ (_26603_, _13242_, _10458_);
  nor _77302_ (_26605_, _26603_, _26585_);
  nor _77303_ (_26606_, _26605_, _04081_);
  or _77304_ (_26607_, _26606_, _26602_);
  and _77305_ (_26608_, _26607_, _03996_);
  nor _77306_ (_26609_, _05363_, _10458_);
  nor _77307_ (_26610_, _26609_, _26585_);
  nor _77308_ (_26611_, _26610_, _03996_);
  nor _77309_ (_26612_, _26611_, _26608_);
  nor _77310_ (_26613_, _26612_, _03729_);
  or _77311_ (_26614_, _26613_, _07390_);
  nor _77312_ (_26616_, _26614_, _26598_);
  and _77313_ (_26617_, _26610_, _07390_);
  or _77314_ (_26618_, _26617_, _04481_);
  nor _77315_ (_26619_, _26618_, _26616_);
  or _77316_ (_26620_, _26619_, _26595_);
  and _77317_ (_26621_, _26620_, _03589_);
  nor _77318_ (_26622_, _13332_, _10458_);
  nor _77319_ (_26623_, _26622_, _26585_);
  nor _77320_ (_26624_, _26623_, _03589_);
  or _77321_ (_26625_, _26624_, _08828_);
  or _77322_ (_26627_, _26625_, _26621_);
  and _77323_ (_26628_, _13347_, _05221_);
  or _77324_ (_26629_, _26585_, _07766_);
  or _77325_ (_26630_, _26629_, _26628_);
  and _77326_ (_26631_, _13339_, _05221_);
  nor _77327_ (_26632_, _26631_, _26585_);
  and _77328_ (_26633_, _26632_, _03601_);
  nor _77329_ (_26634_, _26633_, _03780_);
  and _77330_ (_26635_, _26634_, _26630_);
  and _77331_ (_26636_, _26635_, _26627_);
  nor _77332_ (_26637_, _26636_, _26591_);
  nor _77333_ (_26638_, _26637_, _03622_);
  nor _77334_ (_26639_, _26585_, _05412_);
  not _77335_ (_26640_, _26639_);
  nor _77336_ (_26641_, _26632_, _07777_);
  and _77337_ (_26642_, _26641_, _26640_);
  nor _77338_ (_26643_, _26642_, _26638_);
  nor _77339_ (_26644_, _26643_, _03790_);
  nor _77340_ (_26645_, _26597_, _06828_);
  and _77341_ (_26646_, _26645_, _26640_);
  nor _77342_ (_26649_, _26646_, _03624_);
  not _77343_ (_26650_, _26649_);
  nor _77344_ (_26651_, _26650_, _26644_);
  nor _77345_ (_26652_, _13346_, _10458_);
  or _77346_ (_26653_, _26585_, _07795_);
  nor _77347_ (_26654_, _26653_, _26652_);
  or _77348_ (_26655_, _26654_, _03785_);
  nor _77349_ (_26656_, _26655_, _26651_);
  nor _77350_ (_26657_, _26656_, _26588_);
  nor _77351_ (_26658_, _26657_, _03815_);
  nor _77352_ (_26660_, _26605_, _04246_);
  or _77353_ (_26661_, _26660_, _03447_);
  nor _77354_ (_26662_, _26661_, _26658_);
  and _77355_ (_26663_, _13402_, _05221_);
  or _77356_ (_26664_, _26585_, _03514_);
  nor _77357_ (_26665_, _26664_, _26663_);
  nor _77358_ (_26666_, _26665_, _26662_);
  or _77359_ (_26667_, _26666_, _43004_);
  or _77360_ (_26668_, _43000_, \oc8051_golden_model_1.SBUF [6]);
  and _77361_ (_26669_, _26668_, _41806_);
  and _77362_ (_43595_, _26669_, _26667_);
  not _77363_ (_26671_, \oc8051_golden_model_1.SCON [0]);
  nor _77364_ (_26672_, _05275_, _26671_);
  and _77365_ (_26673_, _12128_, _05275_);
  nor _77366_ (_26674_, _26673_, _26672_);
  nor _77367_ (_26675_, _26674_, _07778_);
  and _77368_ (_26676_, _05275_, _06274_);
  nor _77369_ (_26677_, _26676_, _26672_);
  and _77370_ (_26678_, _26677_, _03601_);
  and _77371_ (_26679_, _05275_, _04620_);
  nor _77372_ (_26681_, _26679_, _26672_);
  and _77373_ (_26682_, _26681_, _07390_);
  and _77374_ (_26683_, _05275_, \oc8051_golden_model_1.ACC [0]);
  nor _77375_ (_26684_, _26683_, _26672_);
  nor _77376_ (_26685_, _26684_, _09029_);
  nor _77377_ (_26686_, _04409_, _26671_);
  or _77378_ (_26687_, _26686_, _26685_);
  and _77379_ (_26688_, _26687_, _04081_);
  nor _77380_ (_26689_, _05666_, _10539_);
  nor _77381_ (_26690_, _26689_, _26672_);
  nor _77382_ (_26692_, _26690_, _04081_);
  or _77383_ (_26693_, _26692_, _26688_);
  and _77384_ (_26694_, _26693_, _04055_);
  nor _77385_ (_26695_, _05922_, _26671_);
  and _77386_ (_26696_, _12021_, _05922_);
  nor _77387_ (_26697_, _26696_, _26695_);
  nor _77388_ (_26698_, _26697_, _04055_);
  nor _77389_ (_26699_, _26698_, _26694_);
  nor _77390_ (_26700_, _26699_, _03723_);
  nor _77391_ (_26701_, _26681_, _03996_);
  or _77392_ (_26703_, _26701_, _26700_);
  and _77393_ (_26704_, _26703_, _03737_);
  nor _77394_ (_26705_, _26684_, _03737_);
  or _77395_ (_26706_, _26705_, _26704_);
  and _77396_ (_26707_, _26706_, _03736_);
  and _77397_ (_26708_, _26672_, _03714_);
  or _77398_ (_26709_, _26708_, _26707_);
  and _77399_ (_26710_, _26709_, _06840_);
  nor _77400_ (_26711_, _26690_, _06840_);
  or _77401_ (_26712_, _26711_, _26710_);
  and _77402_ (_26714_, _26712_, _03710_);
  nor _77403_ (_26715_, _12052_, _10576_);
  nor _77404_ (_26716_, _26715_, _26695_);
  nor _77405_ (_26717_, _26716_, _03710_);
  or _77406_ (_26718_, _26717_, _07390_);
  nor _77407_ (_26719_, _26718_, _26714_);
  nor _77408_ (_26720_, _26719_, _26682_);
  nor _77409_ (_26721_, _26720_, _04481_);
  and _77410_ (_26722_, _06546_, _05275_);
  nor _77411_ (_26723_, _26672_, _07400_);
  not _77412_ (_26725_, _26723_);
  nor _77413_ (_26726_, _26725_, _26722_);
  or _77414_ (_26727_, _26726_, _03222_);
  nor _77415_ (_26728_, _26727_, _26721_);
  nor _77416_ (_26729_, _12109_, _10539_);
  nor _77417_ (_26730_, _26729_, _26672_);
  nor _77418_ (_26731_, _26730_, _03589_);
  or _77419_ (_26732_, _26731_, _03601_);
  nor _77420_ (_26733_, _26732_, _26728_);
  nor _77421_ (_26734_, _26733_, _26678_);
  or _77422_ (_26736_, _26734_, _03600_);
  and _77423_ (_26737_, _12124_, _05275_);
  or _77424_ (_26738_, _26737_, _26672_);
  or _77425_ (_26739_, _26738_, _07766_);
  and _77426_ (_26740_, _26739_, _07778_);
  and _77427_ (_26741_, _26740_, _26736_);
  nor _77428_ (_26742_, _26741_, _26675_);
  nor _77429_ (_26743_, _26742_, _03622_);
  or _77430_ (_26744_, _26677_, _07777_);
  nor _77431_ (_26745_, _26744_, _26689_);
  nor _77432_ (_26747_, _26745_, _26743_);
  nor _77433_ (_26748_, _26747_, _03790_);
  and _77434_ (_26749_, _12005_, _05275_);
  or _77435_ (_26750_, _26749_, _26672_);
  and _77436_ (_26751_, _26750_, _03790_);
  or _77437_ (_26752_, _26751_, _26748_);
  and _77438_ (_26753_, _26752_, _07795_);
  nor _77439_ (_26754_, _12122_, _10539_);
  nor _77440_ (_26755_, _26754_, _26672_);
  nor _77441_ (_26756_, _26755_, _07795_);
  or _77442_ (_26758_, _26756_, _26753_);
  and _77443_ (_26759_, _26758_, _07793_);
  nor _77444_ (_26760_, _12003_, _10539_);
  nor _77445_ (_26761_, _26760_, _26672_);
  nor _77446_ (_26762_, _26761_, _07793_);
  or _77447_ (_26763_, _26762_, _26759_);
  and _77448_ (_26764_, _26763_, _04246_);
  nor _77449_ (_26765_, _26690_, _04246_);
  or _77450_ (_26766_, _26765_, _26764_);
  and _77451_ (_26767_, _26766_, _03823_);
  and _77452_ (_26769_, _26672_, _03453_);
  nor _77453_ (_26770_, _26769_, _03447_);
  not _77454_ (_26771_, _26770_);
  nor _77455_ (_26772_, _26771_, _26767_);
  and _77456_ (_26773_, _26690_, _03447_);
  or _77457_ (_26774_, _26773_, _26772_);
  nand _77458_ (_26775_, _26774_, _43000_);
  or _77459_ (_26776_, _43000_, \oc8051_golden_model_1.SCON [0]);
  and _77460_ (_26777_, _26776_, _41806_);
  and _77461_ (_43596_, _26777_, _26775_);
  not _77462_ (_26779_, \oc8051_golden_model_1.SCON [1]);
  nor _77463_ (_26780_, _05275_, _26779_);
  and _77464_ (_26781_, _06501_, _05275_);
  or _77465_ (_26782_, _26781_, _26780_);
  and _77466_ (_26783_, _26782_, _04481_);
  nor _77467_ (_26784_, _05275_, \oc8051_golden_model_1.SCON [1]);
  and _77468_ (_26785_, _05275_, _03274_);
  nor _77469_ (_26786_, _26785_, _26784_);
  and _77470_ (_26787_, _26786_, _04409_);
  nor _77471_ (_26788_, _04409_, _26779_);
  or _77472_ (_26790_, _26788_, _26787_);
  and _77473_ (_26791_, _26790_, _04081_);
  and _77474_ (_26792_, _12213_, _05275_);
  nor _77475_ (_26793_, _26792_, _26784_);
  and _77476_ (_26794_, _26793_, _03610_);
  or _77477_ (_26795_, _26794_, _26791_);
  and _77478_ (_26796_, _26795_, _04055_);
  and _77479_ (_26797_, _12224_, _05922_);
  nor _77480_ (_26798_, _05922_, _26779_);
  or _77481_ (_26799_, _26798_, _03723_);
  or _77482_ (_26801_, _26799_, _26797_);
  and _77483_ (_26802_, _26801_, _14265_);
  nor _77484_ (_26803_, _26802_, _26796_);
  and _77485_ (_26804_, _05275_, _06764_);
  nor _77486_ (_26805_, _26804_, _26780_);
  and _77487_ (_26806_, _26805_, _03723_);
  nor _77488_ (_26807_, _26806_, _26803_);
  and _77489_ (_26808_, _26807_, _03737_);
  and _77490_ (_26809_, _26786_, _03729_);
  or _77491_ (_26810_, _26809_, _26808_);
  and _77492_ (_26812_, _26810_, _03736_);
  and _77493_ (_26813_, _12211_, _05922_);
  nor _77494_ (_26814_, _26813_, _26798_);
  nor _77495_ (_26815_, _26814_, _03736_);
  or _77496_ (_26816_, _26815_, _26812_);
  and _77497_ (_26817_, _26816_, _06840_);
  and _77498_ (_26818_, _26797_, _12239_);
  or _77499_ (_26819_, _26818_, _26798_);
  and _77500_ (_26820_, _26819_, _03719_);
  or _77501_ (_26821_, _26820_, _26817_);
  and _77502_ (_26823_, _26821_, _03710_);
  nor _77503_ (_26824_, _12256_, _10576_);
  nor _77504_ (_26825_, _26798_, _26824_);
  nor _77505_ (_26826_, _26825_, _03710_);
  or _77506_ (_26827_, _26826_, _07390_);
  nor _77507_ (_26828_, _26827_, _26823_);
  and _77508_ (_26829_, _26805_, _07390_);
  or _77509_ (_26830_, _26829_, _04481_);
  nor _77510_ (_26831_, _26830_, _26828_);
  or _77511_ (_26832_, _26831_, _26783_);
  and _77512_ (_26834_, _26832_, _03589_);
  nor _77513_ (_26835_, _12313_, _10539_);
  nor _77514_ (_26836_, _26835_, _26780_);
  nor _77515_ (_26837_, _26836_, _03589_);
  nor _77516_ (_26838_, _26837_, _26834_);
  nor _77517_ (_26839_, _26838_, _08828_);
  not _77518_ (_26840_, _26784_);
  nor _77519_ (_26841_, _12327_, _10539_);
  nor _77520_ (_26842_, _26841_, _07766_);
  and _77521_ (_26843_, _05275_, _04303_);
  nor _77522_ (_26845_, _26843_, _05886_);
  or _77523_ (_26846_, _26845_, _26842_);
  and _77524_ (_26847_, _26846_, _26840_);
  nor _77525_ (_26848_, _26847_, _26839_);
  nor _77526_ (_26849_, _26848_, _03780_);
  nor _77527_ (_26850_, _12333_, _10539_);
  nor _77528_ (_26851_, _26850_, _07778_);
  and _77529_ (_26852_, _26851_, _26840_);
  nor _77530_ (_26853_, _26852_, _26849_);
  nor _77531_ (_26854_, _26853_, _03622_);
  nor _77532_ (_26856_, _12207_, _10539_);
  nor _77533_ (_26857_, _26856_, _07777_);
  and _77534_ (_26858_, _26857_, _26840_);
  nor _77535_ (_26859_, _26858_, _26854_);
  nor _77536_ (_26860_, _26859_, _03790_);
  nor _77537_ (_26861_, _26780_, _05618_);
  nor _77538_ (_26862_, _26861_, _06828_);
  and _77539_ (_26863_, _26862_, _26786_);
  nor _77540_ (_26864_, _26863_, _26860_);
  or _77541_ (_26865_, _26864_, _18499_);
  and _77542_ (_26867_, _26785_, _05617_);
  nor _77543_ (_26868_, _26867_, _07793_);
  and _77544_ (_26869_, _26868_, _26840_);
  nor _77545_ (_26870_, _26869_, _03815_);
  and _77546_ (_26871_, _26843_, _05617_);
  or _77547_ (_26872_, _26784_, _07795_);
  or _77548_ (_26873_, _26872_, _26871_);
  and _77549_ (_26874_, _26873_, _26870_);
  and _77550_ (_26875_, _26874_, _26865_);
  nor _77551_ (_26876_, _26793_, _04246_);
  or _77552_ (_26878_, _26876_, _03453_);
  nor _77553_ (_26879_, _26878_, _26875_);
  nor _77554_ (_26880_, _26814_, _03823_);
  or _77555_ (_26881_, _26880_, _03447_);
  nor _77556_ (_26882_, _26881_, _26879_);
  nor _77557_ (_26883_, _26792_, _26780_);
  and _77558_ (_26884_, _26883_, _03447_);
  nor _77559_ (_26885_, _26884_, _26882_);
  or _77560_ (_26886_, _26885_, _43004_);
  or _77561_ (_26887_, _43000_, \oc8051_golden_model_1.SCON [1]);
  and _77562_ (_26889_, _26887_, _41806_);
  and _77563_ (_43599_, _26889_, _26886_);
  not _77564_ (_26890_, \oc8051_golden_model_1.SCON [2]);
  nor _77565_ (_26891_, _05275_, _26890_);
  and _77566_ (_26892_, _05275_, _06332_);
  nor _77567_ (_26893_, _26892_, _26891_);
  and _77568_ (_26894_, _26893_, _03601_);
  nor _77569_ (_26895_, _10539_, _04875_);
  nor _77570_ (_26896_, _26895_, _26891_);
  and _77571_ (_26897_, _26896_, _07390_);
  nor _77572_ (_26899_, _26896_, _03996_);
  nor _77573_ (_26900_, _05922_, _26890_);
  and _77574_ (_26901_, _12411_, _05922_);
  nor _77575_ (_26902_, _26901_, _26900_);
  and _77576_ (_26903_, _26902_, _03715_);
  nor _77577_ (_26904_, _12416_, _10539_);
  nor _77578_ (_26905_, _26904_, _26891_);
  nor _77579_ (_26906_, _26905_, _04081_);
  nor _77580_ (_26907_, _04409_, _26890_);
  and _77581_ (_26908_, _05275_, \oc8051_golden_model_1.ACC [2]);
  nor _77582_ (_26910_, _26908_, _26891_);
  nor _77583_ (_26911_, _26910_, _09029_);
  nor _77584_ (_26912_, _26911_, _26907_);
  nor _77585_ (_26913_, _26912_, _03610_);
  or _77586_ (_26914_, _26913_, _03715_);
  nor _77587_ (_26915_, _26914_, _26906_);
  nor _77588_ (_26916_, _26915_, _26903_);
  and _77589_ (_26917_, _26916_, _03996_);
  or _77590_ (_26918_, _26917_, _26899_);
  and _77591_ (_26919_, _26918_, _03737_);
  nor _77592_ (_26921_, _26910_, _03737_);
  or _77593_ (_26922_, _26921_, _26919_);
  and _77594_ (_26923_, _26922_, _03736_);
  and _77595_ (_26924_, _12409_, _05922_);
  nor _77596_ (_26925_, _26924_, _26900_);
  nor _77597_ (_26926_, _26925_, _03736_);
  or _77598_ (_26927_, _26926_, _26923_);
  and _77599_ (_26928_, _26927_, _06840_);
  nor _77600_ (_26929_, _26900_, _12443_);
  nor _77601_ (_26930_, _26929_, _26902_);
  and _77602_ (_26931_, _26930_, _03719_);
  or _77603_ (_26932_, _26931_, _26928_);
  and _77604_ (_26933_, _26932_, _03710_);
  nor _77605_ (_26934_, _12461_, _10576_);
  nor _77606_ (_26935_, _26934_, _26900_);
  nor _77607_ (_26936_, _26935_, _03710_);
  nor _77608_ (_26937_, _26936_, _07390_);
  not _77609_ (_26938_, _26937_);
  nor _77610_ (_26939_, _26938_, _26933_);
  nor _77611_ (_26940_, _26939_, _26897_);
  nor _77612_ (_26943_, _26940_, _04481_);
  and _77613_ (_26944_, _06637_, _05275_);
  nor _77614_ (_26945_, _26891_, _07400_);
  not _77615_ (_26946_, _26945_);
  nor _77616_ (_26947_, _26946_, _26944_);
  or _77617_ (_26948_, _26947_, _03222_);
  nor _77618_ (_26949_, _26948_, _26943_);
  nor _77619_ (_26950_, _12519_, _10539_);
  nor _77620_ (_26951_, _26891_, _26950_);
  nor _77621_ (_26952_, _26951_, _03589_);
  or _77622_ (_26954_, _26952_, _03601_);
  nor _77623_ (_26955_, _26954_, _26949_);
  nor _77624_ (_26956_, _26955_, _26894_);
  or _77625_ (_26957_, _26956_, _03600_);
  and _77626_ (_26958_, _12533_, _05275_);
  or _77627_ (_26959_, _26958_, _26891_);
  or _77628_ (_26960_, _26959_, _07766_);
  and _77629_ (_26961_, _26960_, _07778_);
  and _77630_ (_26962_, _26961_, _26957_);
  and _77631_ (_26963_, _12539_, _05275_);
  nor _77632_ (_26965_, _26963_, _26891_);
  nor _77633_ (_26966_, _26965_, _07778_);
  nor _77634_ (_26967_, _26966_, _26962_);
  nor _77635_ (_26968_, _26967_, _03622_);
  nor _77636_ (_26969_, _26891_, _05718_);
  not _77637_ (_26970_, _26969_);
  nor _77638_ (_26971_, _26893_, _07777_);
  and _77639_ (_26972_, _26971_, _26970_);
  nor _77640_ (_26973_, _26972_, _26968_);
  nor _77641_ (_26974_, _26973_, _03790_);
  nor _77642_ (_26976_, _26910_, _06828_);
  and _77643_ (_26977_, _26976_, _26970_);
  or _77644_ (_26978_, _26977_, _26974_);
  and _77645_ (_26979_, _26978_, _07795_);
  nor _77646_ (_26980_, _12532_, _10539_);
  nor _77647_ (_26981_, _26980_, _26891_);
  nor _77648_ (_26982_, _26981_, _07795_);
  or _77649_ (_26983_, _26982_, _26979_);
  and _77650_ (_26984_, _26983_, _07793_);
  nor _77651_ (_26985_, _12538_, _10539_);
  nor _77652_ (_26987_, _26985_, _26891_);
  nor _77653_ (_26988_, _26987_, _07793_);
  or _77654_ (_26989_, _26988_, _26984_);
  and _77655_ (_26990_, _26989_, _04246_);
  nor _77656_ (_26991_, _26905_, _04246_);
  or _77657_ (_26992_, _26991_, _26990_);
  and _77658_ (_26993_, _26992_, _03823_);
  nor _77659_ (_26994_, _26925_, _03823_);
  or _77660_ (_26995_, _26994_, _26993_);
  and _77661_ (_26996_, _26995_, _03514_);
  and _77662_ (_26998_, _12592_, _05275_);
  nor _77663_ (_26999_, _26998_, _26891_);
  nor _77664_ (_27000_, _26999_, _03514_);
  or _77665_ (_27001_, _27000_, _26996_);
  or _77666_ (_27002_, _27001_, _43004_);
  or _77667_ (_27003_, _43000_, \oc8051_golden_model_1.SCON [2]);
  and _77668_ (_27004_, _27003_, _41806_);
  and _77669_ (_43600_, _27004_, _27002_);
  not _77670_ (_27005_, \oc8051_golden_model_1.SCON [3]);
  nor _77671_ (_27006_, _05275_, _27005_);
  and _77672_ (_27008_, _05275_, _06276_);
  nor _77673_ (_27009_, _27008_, _27006_);
  and _77674_ (_27010_, _27009_, _03601_);
  nor _77675_ (_27011_, _10539_, _05005_);
  nor _77676_ (_27012_, _27011_, _27006_);
  and _77677_ (_27013_, _27012_, _07390_);
  and _77678_ (_27014_, _05275_, \oc8051_golden_model_1.ACC [3]);
  nor _77679_ (_27015_, _27014_, _27006_);
  nor _77680_ (_27016_, _27015_, _09029_);
  nor _77681_ (_27017_, _04409_, _27005_);
  or _77682_ (_27019_, _27017_, _27016_);
  and _77683_ (_27020_, _27019_, _04081_);
  nor _77684_ (_27021_, _12627_, _10539_);
  nor _77685_ (_27022_, _27021_, _27006_);
  nor _77686_ (_27023_, _27022_, _04081_);
  or _77687_ (_27024_, _27023_, _27020_);
  and _77688_ (_27025_, _27024_, _04055_);
  nor _77689_ (_27026_, _05922_, _27005_);
  and _77690_ (_27027_, _12631_, _05922_);
  nor _77691_ (_27028_, _27027_, _27026_);
  nor _77692_ (_27030_, _27028_, _04055_);
  or _77693_ (_27031_, _27030_, _03723_);
  or _77694_ (_27032_, _27031_, _27025_);
  nand _77695_ (_27033_, _27012_, _03723_);
  and _77696_ (_27034_, _27033_, _27032_);
  and _77697_ (_27035_, _27034_, _03737_);
  nor _77698_ (_27036_, _27015_, _03737_);
  or _77699_ (_27037_, _27036_, _27035_);
  and _77700_ (_27038_, _27037_, _03736_);
  and _77701_ (_27039_, _12641_, _05922_);
  nor _77702_ (_27040_, _27039_, _27026_);
  nor _77703_ (_27041_, _27040_, _03736_);
  or _77704_ (_27042_, _27041_, _03719_);
  or _77705_ (_27043_, _27042_, _27038_);
  nor _77706_ (_27044_, _27026_, _12648_);
  nor _77707_ (_27045_, _27044_, _27028_);
  or _77708_ (_27046_, _27045_, _06840_);
  and _77709_ (_27047_, _27046_, _03710_);
  and _77710_ (_27048_, _27047_, _27043_);
  nor _77711_ (_27049_, _12612_, _10576_);
  nor _77712_ (_27052_, _27049_, _27026_);
  nor _77713_ (_27053_, _27052_, _03710_);
  nor _77714_ (_27054_, _27053_, _07390_);
  not _77715_ (_27055_, _27054_);
  nor _77716_ (_27056_, _27055_, _27048_);
  nor _77717_ (_27057_, _27056_, _27013_);
  nor _77718_ (_27058_, _27057_, _04481_);
  and _77719_ (_27059_, _06592_, _05275_);
  nor _77720_ (_27060_, _27006_, _07400_);
  not _77721_ (_27061_, _27060_);
  nor _77722_ (_27063_, _27061_, _27059_);
  or _77723_ (_27064_, _27063_, _03222_);
  nor _77724_ (_27065_, _27064_, _27058_);
  nor _77725_ (_27066_, _12718_, _10539_);
  nor _77726_ (_27067_, _27006_, _27066_);
  nor _77727_ (_27068_, _27067_, _03589_);
  or _77728_ (_27069_, _27068_, _03601_);
  nor _77729_ (_27070_, _27069_, _27065_);
  nor _77730_ (_27071_, _27070_, _27010_);
  or _77731_ (_27072_, _27071_, _03600_);
  and _77732_ (_27074_, _12733_, _05275_);
  or _77733_ (_27075_, _27074_, _27006_);
  or _77734_ (_27076_, _27075_, _07766_);
  and _77735_ (_27077_, _27076_, _07778_);
  and _77736_ (_27078_, _27077_, _27072_);
  and _77737_ (_27079_, _12739_, _05275_);
  nor _77738_ (_27080_, _27079_, _27006_);
  nor _77739_ (_27081_, _27080_, _07778_);
  nor _77740_ (_27082_, _27081_, _27078_);
  nor _77741_ (_27083_, _27082_, _03622_);
  nor _77742_ (_27085_, _27006_, _05567_);
  not _77743_ (_27086_, _27085_);
  nor _77744_ (_27087_, _27009_, _07777_);
  and _77745_ (_27088_, _27087_, _27086_);
  nor _77746_ (_27089_, _27088_, _27083_);
  nor _77747_ (_27090_, _27089_, _03790_);
  nor _77748_ (_27091_, _27015_, _06828_);
  and _77749_ (_27092_, _27091_, _27086_);
  nor _77750_ (_27093_, _27092_, _03624_);
  not _77751_ (_27094_, _27093_);
  nor _77752_ (_27096_, _27094_, _27090_);
  nor _77753_ (_27097_, _12732_, _10539_);
  or _77754_ (_27098_, _27006_, _07795_);
  nor _77755_ (_27099_, _27098_, _27097_);
  or _77756_ (_27100_, _27099_, _03785_);
  nor _77757_ (_27101_, _27100_, _27096_);
  nor _77758_ (_27102_, _12738_, _10539_);
  nor _77759_ (_27103_, _27102_, _27006_);
  nor _77760_ (_27104_, _27103_, _07793_);
  or _77761_ (_27105_, _27104_, _27101_);
  and _77762_ (_27107_, _27105_, _04246_);
  nor _77763_ (_27108_, _27022_, _04246_);
  or _77764_ (_27109_, _27108_, _27107_);
  and _77765_ (_27110_, _27109_, _03823_);
  nor _77766_ (_27111_, _27040_, _03823_);
  or _77767_ (_27112_, _27111_, _27110_);
  and _77768_ (_27113_, _27112_, _03514_);
  and _77769_ (_27114_, _12794_, _05275_);
  nor _77770_ (_27115_, _27114_, _27006_);
  nor _77771_ (_27116_, _27115_, _03514_);
  or _77772_ (_27118_, _27116_, _27113_);
  or _77773_ (_27119_, _27118_, _43004_);
  or _77774_ (_27120_, _43000_, \oc8051_golden_model_1.SCON [3]);
  and _77775_ (_27121_, _27120_, _41806_);
  and _77776_ (_43601_, _27121_, _27119_);
  not _77777_ (_27122_, \oc8051_golden_model_1.SCON [4]);
  nor _77778_ (_27123_, _05275_, _27122_);
  nor _77779_ (_27124_, _05777_, _10539_);
  nor _77780_ (_27125_, _27124_, _27123_);
  and _77781_ (_27126_, _27125_, _07390_);
  nor _77782_ (_27128_, _05922_, _27122_);
  and _77783_ (_27129_, _12827_, _05922_);
  nor _77784_ (_27130_, _27129_, _27128_);
  nor _77785_ (_27131_, _27130_, _03736_);
  and _77786_ (_27132_, _05275_, \oc8051_golden_model_1.ACC [4]);
  nor _77787_ (_27133_, _27132_, _27123_);
  nor _77788_ (_27134_, _27133_, _09029_);
  nor _77789_ (_27135_, _04409_, _27122_);
  or _77790_ (_27136_, _27135_, _27134_);
  and _77791_ (_27137_, _27136_, _04081_);
  nor _77792_ (_27139_, _12841_, _10539_);
  nor _77793_ (_27140_, _27139_, _27123_);
  nor _77794_ (_27141_, _27140_, _04081_);
  or _77795_ (_27142_, _27141_, _27137_);
  and _77796_ (_27143_, _27142_, _04055_);
  and _77797_ (_27144_, _12845_, _05922_);
  nor _77798_ (_27145_, _27144_, _27128_);
  nor _77799_ (_27146_, _27145_, _04055_);
  or _77800_ (_27147_, _27146_, _03723_);
  or _77801_ (_27148_, _27147_, _27143_);
  nand _77802_ (_27150_, _27125_, _03723_);
  and _77803_ (_27151_, _27150_, _27148_);
  and _77804_ (_27152_, _27151_, _03737_);
  nor _77805_ (_27153_, _27133_, _03737_);
  or _77806_ (_27154_, _27153_, _27152_);
  and _77807_ (_27155_, _27154_, _03736_);
  nor _77808_ (_27156_, _27155_, _27131_);
  nor _77809_ (_27157_, _27156_, _03719_);
  nor _77810_ (_27158_, _27128_, _12860_);
  or _77811_ (_27159_, _27145_, _06840_);
  nor _77812_ (_27161_, _27159_, _27158_);
  nor _77813_ (_27162_, _27161_, _27157_);
  nor _77814_ (_27163_, _27162_, _03505_);
  nor _77815_ (_27164_, _12825_, _10576_);
  nor _77816_ (_27165_, _27164_, _27128_);
  nor _77817_ (_27166_, _27165_, _03710_);
  nor _77818_ (_27167_, _27166_, _07390_);
  not _77819_ (_27168_, _27167_);
  nor _77820_ (_27169_, _27168_, _27163_);
  nor _77821_ (_27170_, _27169_, _27126_);
  nor _77822_ (_27172_, _27170_, _04481_);
  and _77823_ (_27173_, _06730_, _05275_);
  nor _77824_ (_27174_, _27123_, _07400_);
  not _77825_ (_27175_, _27174_);
  nor _77826_ (_27176_, _27175_, _27173_);
  nor _77827_ (_27177_, _27176_, _03222_);
  not _77828_ (_27178_, _27177_);
  nor _77829_ (_27179_, _27178_, _27172_);
  nor _77830_ (_27180_, _12933_, _10539_);
  nor _77831_ (_27181_, _27180_, _27123_);
  nor _77832_ (_27183_, _27181_, _03589_);
  or _77833_ (_27184_, _27183_, _08828_);
  or _77834_ (_27185_, _27184_, _27179_);
  and _77835_ (_27186_, _12821_, _05275_);
  or _77836_ (_27187_, _27123_, _07766_);
  or _77837_ (_27188_, _27187_, _27186_);
  and _77838_ (_27189_, _06298_, _05275_);
  nor _77839_ (_27190_, _27189_, _27123_);
  and _77840_ (_27191_, _27190_, _03601_);
  nor _77841_ (_27192_, _27191_, _03780_);
  and _77842_ (_27194_, _27192_, _27188_);
  and _77843_ (_27195_, _27194_, _27185_);
  and _77844_ (_27196_, _12817_, _05275_);
  nor _77845_ (_27197_, _27196_, _27123_);
  nor _77846_ (_27198_, _27197_, _07778_);
  nor _77847_ (_27199_, _27198_, _27195_);
  nor _77848_ (_27200_, _27199_, _03622_);
  nor _77849_ (_27201_, _27123_, _05825_);
  not _77850_ (_27202_, _27201_);
  nor _77851_ (_27203_, _27190_, _07777_);
  and _77852_ (_27205_, _27203_, _27202_);
  nor _77853_ (_27206_, _27205_, _27200_);
  nor _77854_ (_27207_, _27206_, _03790_);
  nor _77855_ (_27208_, _27133_, _06828_);
  and _77856_ (_27209_, _27208_, _27202_);
  nor _77857_ (_27210_, _27209_, _03624_);
  not _77858_ (_27211_, _27210_);
  nor _77859_ (_27212_, _27211_, _27207_);
  nor _77860_ (_27213_, _12819_, _10539_);
  or _77861_ (_27214_, _27123_, _07795_);
  nor _77862_ (_27216_, _27214_, _27213_);
  or _77863_ (_27217_, _27216_, _03785_);
  nor _77864_ (_27218_, _27217_, _27212_);
  nor _77865_ (_27219_, _12816_, _10539_);
  nor _77866_ (_27220_, _27219_, _27123_);
  nor _77867_ (_27221_, _27220_, _07793_);
  or _77868_ (_27222_, _27221_, _27218_);
  and _77869_ (_27223_, _27222_, _04246_);
  nor _77870_ (_27224_, _27140_, _04246_);
  or _77871_ (_27225_, _27224_, _27223_);
  and _77872_ (_27227_, _27225_, _03823_);
  nor _77873_ (_27228_, _27130_, _03823_);
  or _77874_ (_27229_, _27228_, _27227_);
  and _77875_ (_27230_, _27229_, _03514_);
  and _77876_ (_27231_, _13003_, _05275_);
  nor _77877_ (_27232_, _27231_, _27123_);
  nor _77878_ (_27233_, _27232_, _03514_);
  or _77879_ (_27234_, _27233_, _27230_);
  or _77880_ (_27235_, _27234_, _43004_);
  or _77881_ (_27236_, _43000_, \oc8051_golden_model_1.SCON [4]);
  and _77882_ (_27238_, _27236_, _41806_);
  and _77883_ (_43602_, _27238_, _27235_);
  not _77884_ (_27239_, \oc8051_golden_model_1.SCON [5]);
  nor _77885_ (_27240_, _05275_, _27239_);
  and _77886_ (_27241_, _06684_, _05275_);
  or _77887_ (_27242_, _27241_, _27240_);
  and _77888_ (_27243_, _27242_, _04481_);
  and _77889_ (_27244_, _05275_, \oc8051_golden_model_1.ACC [5]);
  nor _77890_ (_27245_, _27244_, _27240_);
  nor _77891_ (_27246_, _27245_, _09029_);
  nor _77892_ (_27248_, _04409_, _27239_);
  or _77893_ (_27249_, _27248_, _27246_);
  and _77894_ (_27250_, _27249_, _04081_);
  nor _77895_ (_27251_, _13014_, _10539_);
  nor _77896_ (_27252_, _27251_, _27240_);
  nor _77897_ (_27253_, _27252_, _04081_);
  or _77898_ (_27254_, _27253_, _27250_);
  and _77899_ (_27255_, _27254_, _04055_);
  nor _77900_ (_27256_, _05922_, _27239_);
  and _77901_ (_27257_, _13037_, _05922_);
  nor _77902_ (_27258_, _27257_, _27256_);
  nor _77903_ (_27259_, _27258_, _04055_);
  or _77904_ (_27260_, _27259_, _03723_);
  or _77905_ (_27261_, _27260_, _27255_);
  nor _77906_ (_27262_, _05469_, _10539_);
  nor _77907_ (_27263_, _27262_, _27240_);
  nand _77908_ (_27264_, _27263_, _03723_);
  and _77909_ (_27265_, _27264_, _27261_);
  and _77910_ (_27266_, _27265_, _03737_);
  nor _77911_ (_27267_, _27245_, _03737_);
  or _77912_ (_27270_, _27267_, _27266_);
  and _77913_ (_27271_, _27270_, _03736_);
  and _77914_ (_27272_, _13047_, _05922_);
  nor _77915_ (_27273_, _27272_, _27256_);
  nor _77916_ (_27274_, _27273_, _03736_);
  or _77917_ (_27275_, _27274_, _27271_);
  and _77918_ (_27276_, _27275_, _06840_);
  nor _77919_ (_27277_, _27256_, _13054_);
  nor _77920_ (_27278_, _27277_, _27258_);
  and _77921_ (_27279_, _27278_, _03719_);
  or _77922_ (_27281_, _27279_, _27276_);
  and _77923_ (_27282_, _27281_, _03710_);
  nor _77924_ (_27283_, _13020_, _10576_);
  nor _77925_ (_27284_, _27283_, _27256_);
  nor _77926_ (_27285_, _27284_, _03710_);
  nor _77927_ (_27286_, _27285_, _07390_);
  not _77928_ (_27287_, _27286_);
  nor _77929_ (_27288_, _27287_, _27282_);
  and _77930_ (_27289_, _27263_, _07390_);
  or _77931_ (_27290_, _27289_, _04481_);
  nor _77932_ (_27292_, _27290_, _27288_);
  or _77933_ (_27293_, _27292_, _27243_);
  and _77934_ (_27294_, _27293_, _03589_);
  nor _77935_ (_27295_, _13127_, _10539_);
  nor _77936_ (_27296_, _27295_, _27240_);
  nor _77937_ (_27297_, _27296_, _03589_);
  or _77938_ (_27298_, _27297_, _08828_);
  or _77939_ (_27299_, _27298_, _27294_);
  and _77940_ (_27300_, _13141_, _05275_);
  or _77941_ (_27301_, _27240_, _07766_);
  or _77942_ (_27303_, _27301_, _27300_);
  and _77943_ (_27304_, _06306_, _05275_);
  nor _77944_ (_27305_, _27304_, _27240_);
  and _77945_ (_27306_, _27305_, _03601_);
  nor _77946_ (_27307_, _27306_, _03780_);
  and _77947_ (_27308_, _27307_, _27303_);
  and _77948_ (_27309_, _27308_, _27299_);
  and _77949_ (_27310_, _13147_, _05275_);
  nor _77950_ (_27311_, _27310_, _27240_);
  nor _77951_ (_27312_, _27311_, _07778_);
  nor _77952_ (_27314_, _27312_, _27309_);
  nor _77953_ (_27315_, _27314_, _03622_);
  nor _77954_ (_27316_, _27240_, _05518_);
  not _77955_ (_27317_, _27316_);
  nor _77956_ (_27318_, _27305_, _07777_);
  and _77957_ (_27319_, _27318_, _27317_);
  nor _77958_ (_27320_, _27319_, _27315_);
  nor _77959_ (_27321_, _27320_, _03790_);
  nor _77960_ (_27322_, _27245_, _06828_);
  and _77961_ (_27323_, _27322_, _27317_);
  nor _77962_ (_27325_, _27323_, _03624_);
  not _77963_ (_27326_, _27325_);
  nor _77964_ (_27327_, _27326_, _27321_);
  nor _77965_ (_27328_, _13140_, _10539_);
  or _77966_ (_27329_, _27240_, _07795_);
  nor _77967_ (_27330_, _27329_, _27328_);
  or _77968_ (_27331_, _27330_, _03785_);
  nor _77969_ (_27332_, _27331_, _27327_);
  nor _77970_ (_27333_, _13146_, _10539_);
  nor _77971_ (_27334_, _27333_, _27240_);
  nor _77972_ (_27336_, _27334_, _07793_);
  or _77973_ (_27337_, _27336_, _27332_);
  and _77974_ (_27338_, _27337_, _04246_);
  nor _77975_ (_27339_, _27252_, _04246_);
  or _77976_ (_27340_, _27339_, _27338_);
  and _77977_ (_27341_, _27340_, _03823_);
  nor _77978_ (_27342_, _27273_, _03823_);
  or _77979_ (_27343_, _27342_, _27341_);
  and _77980_ (_27344_, _27343_, _03514_);
  and _77981_ (_27345_, _13199_, _05275_);
  nor _77982_ (_27347_, _27345_, _27240_);
  nor _77983_ (_27348_, _27347_, _03514_);
  or _77984_ (_27349_, _27348_, _27344_);
  or _77985_ (_27350_, _27349_, _43004_);
  or _77986_ (_27351_, _43000_, \oc8051_golden_model_1.SCON [5]);
  and _77987_ (_27352_, _27351_, _41806_);
  and _77988_ (_43603_, _27352_, _27350_);
  not _77989_ (_27353_, \oc8051_golden_model_1.SCON [6]);
  nor _77990_ (_27354_, _05275_, _27353_);
  and _77991_ (_27355_, _06455_, _05275_);
  or _77992_ (_27357_, _27355_, _27354_);
  and _77993_ (_27358_, _27357_, _04481_);
  and _77994_ (_27359_, _05275_, \oc8051_golden_model_1.ACC [6]);
  nor _77995_ (_27360_, _27359_, _27354_);
  nor _77996_ (_27361_, _27360_, _09029_);
  nor _77997_ (_27362_, _04409_, _27353_);
  or _77998_ (_27363_, _27362_, _27361_);
  and _77999_ (_27364_, _27363_, _04081_);
  nor _78000_ (_27365_, _13242_, _10539_);
  nor _78001_ (_27366_, _27365_, _27354_);
  nor _78002_ (_27368_, _27366_, _04081_);
  or _78003_ (_27369_, _27368_, _27364_);
  and _78004_ (_27370_, _27369_, _04055_);
  nor _78005_ (_27371_, _05922_, _27353_);
  and _78006_ (_27372_, _13229_, _05922_);
  nor _78007_ (_27373_, _27372_, _27371_);
  nor _78008_ (_27374_, _27373_, _04055_);
  or _78009_ (_27375_, _27374_, _03723_);
  or _78010_ (_27376_, _27375_, _27370_);
  nor _78011_ (_27377_, _05363_, _10539_);
  nor _78012_ (_27379_, _27377_, _27354_);
  nand _78013_ (_27380_, _27379_, _03723_);
  and _78014_ (_27381_, _27380_, _27376_);
  and _78015_ (_27382_, _27381_, _03737_);
  nor _78016_ (_27383_, _27360_, _03737_);
  or _78017_ (_27384_, _27383_, _27382_);
  and _78018_ (_27385_, _27384_, _03736_);
  and _78019_ (_27386_, _13253_, _05922_);
  nor _78020_ (_27387_, _27386_, _27371_);
  nor _78021_ (_27388_, _27387_, _03736_);
  or _78022_ (_27390_, _27388_, _03719_);
  or _78023_ (_27391_, _27390_, _27385_);
  nor _78024_ (_27392_, _27371_, _13260_);
  nor _78025_ (_27393_, _27392_, _27373_);
  or _78026_ (_27394_, _27393_, _06840_);
  and _78027_ (_27395_, _27394_, _03710_);
  and _78028_ (_27396_, _27395_, _27391_);
  nor _78029_ (_27397_, _13226_, _10576_);
  nor _78030_ (_27398_, _27397_, _27371_);
  nor _78031_ (_27399_, _27398_, _03710_);
  nor _78032_ (_27401_, _27399_, _07390_);
  not _78033_ (_27402_, _27401_);
  nor _78034_ (_27403_, _27402_, _27396_);
  and _78035_ (_27404_, _27379_, _07390_);
  or _78036_ (_27405_, _27404_, _04481_);
  nor _78037_ (_27406_, _27405_, _27403_);
  or _78038_ (_27407_, _27406_, _27358_);
  and _78039_ (_27408_, _27407_, _03589_);
  nor _78040_ (_27409_, _13332_, _10539_);
  nor _78041_ (_27410_, _27409_, _27354_);
  nor _78042_ (_27412_, _27410_, _03589_);
  or _78043_ (_27413_, _27412_, _08828_);
  or _78044_ (_27414_, _27413_, _27408_);
  and _78045_ (_27415_, _13347_, _05275_);
  or _78046_ (_27416_, _27354_, _07766_);
  or _78047_ (_27417_, _27416_, _27415_);
  and _78048_ (_27418_, _13339_, _05275_);
  nor _78049_ (_27419_, _27418_, _27354_);
  and _78050_ (_27420_, _27419_, _03601_);
  nor _78051_ (_27421_, _27420_, _03780_);
  and _78052_ (_27423_, _27421_, _27417_);
  and _78053_ (_27424_, _27423_, _27414_);
  and _78054_ (_27425_, _13353_, _05275_);
  nor _78055_ (_27426_, _27425_, _27354_);
  nor _78056_ (_27427_, _27426_, _07778_);
  nor _78057_ (_27428_, _27427_, _27424_);
  nor _78058_ (_27429_, _27428_, _03622_);
  nor _78059_ (_27430_, _27354_, _05412_);
  not _78060_ (_27431_, _27430_);
  nor _78061_ (_27432_, _27419_, _07777_);
  and _78062_ (_27434_, _27432_, _27431_);
  nor _78063_ (_27435_, _27434_, _27429_);
  nor _78064_ (_27436_, _27435_, _03790_);
  nor _78065_ (_27437_, _27360_, _06828_);
  and _78066_ (_27438_, _27437_, _27431_);
  nor _78067_ (_27439_, _27438_, _03624_);
  not _78068_ (_27440_, _27439_);
  nor _78069_ (_27441_, _27440_, _27436_);
  nor _78070_ (_27442_, _13346_, _10539_);
  or _78071_ (_27443_, _27354_, _07795_);
  nor _78072_ (_27445_, _27443_, _27442_);
  or _78073_ (_27446_, _27445_, _03785_);
  nor _78074_ (_27447_, _27446_, _27441_);
  nor _78075_ (_27448_, _13352_, _10539_);
  nor _78076_ (_27449_, _27448_, _27354_);
  nor _78077_ (_27450_, _27449_, _07793_);
  or _78078_ (_27451_, _27450_, _27447_);
  and _78079_ (_27452_, _27451_, _04246_);
  nor _78080_ (_27453_, _27366_, _04246_);
  or _78081_ (_27454_, _27453_, _27452_);
  and _78082_ (_27456_, _27454_, _03823_);
  nor _78083_ (_27457_, _27387_, _03823_);
  or _78084_ (_27458_, _27457_, _27456_);
  and _78085_ (_27459_, _27458_, _03514_);
  and _78086_ (_27460_, _13402_, _05275_);
  nor _78087_ (_27461_, _27460_, _27354_);
  nor _78088_ (_27462_, _27461_, _03514_);
  or _78089_ (_27463_, _27462_, _27459_);
  or _78090_ (_27464_, _27463_, _43004_);
  or _78091_ (_27465_, _43000_, \oc8051_golden_model_1.SCON [6]);
  and _78092_ (_27467_, _27465_, _41806_);
  and _78093_ (_43604_, _27467_, _27464_);
  nor _78094_ (_27468_, _05300_, _03498_);
  nor _78095_ (_27469_, _05666_, _10706_);
  nor _78096_ (_27470_, _27469_, _27468_);
  and _78097_ (_27471_, _27470_, _17166_);
  and _78098_ (_27472_, _05300_, \oc8051_golden_model_1.ACC [0]);
  nor _78099_ (_27473_, _27472_, _27468_);
  nor _78100_ (_27474_, _27473_, _09029_);
  nor _78101_ (_27475_, _04409_, _03498_);
  or _78102_ (_27477_, _27475_, _27474_);
  and _78103_ (_27478_, _27477_, _04081_);
  nor _78104_ (_27479_, _27470_, _04081_);
  or _78105_ (_27480_, _27479_, _27478_);
  and _78106_ (_27481_, _27480_, _03996_);
  nor _78107_ (_27482_, _27481_, _04089_);
  and _78108_ (_27483_, _27473_, _03729_);
  nor _78109_ (_27484_, _27483_, _03508_);
  not _78110_ (_27485_, _27484_);
  nor _78111_ (_27486_, _27485_, _27482_);
  nor _78112_ (_27488_, _07390_, _04657_);
  not _78113_ (_27489_, _27488_);
  nor _78114_ (_27490_, _27489_, _27486_);
  not _78115_ (_27491_, _27468_);
  and _78116_ (_27492_, _05300_, _04620_);
  nor _78117_ (_27493_, _27492_, _06838_);
  and _78118_ (_27494_, _27493_, _27491_);
  nor _78119_ (_27495_, _27494_, _27490_);
  nor _78120_ (_27496_, _27495_, _04481_);
  and _78121_ (_27497_, _06546_, _05300_);
  nor _78122_ (_27499_, _27468_, _07400_);
  not _78123_ (_27500_, _27499_);
  nor _78124_ (_27501_, _27500_, _27497_);
  nor _78125_ (_27502_, _27501_, _27496_);
  nor _78126_ (_27503_, _27502_, _03222_);
  nor _78127_ (_27504_, _12109_, _10706_);
  or _78128_ (_27505_, _27468_, _03589_);
  nor _78129_ (_27506_, _27505_, _27504_);
  or _78130_ (_27507_, _27506_, _03601_);
  nor _78131_ (_27508_, _27507_, _27503_);
  and _78132_ (_27510_, _05300_, _06274_);
  nor _78133_ (_27511_, _27510_, _27468_);
  nand _78134_ (_27512_, _27511_, _07766_);
  and _78135_ (_27513_, _27512_, _08828_);
  nor _78136_ (_27514_, _27513_, _27508_);
  and _78137_ (_27515_, _12124_, _05300_);
  nor _78138_ (_27516_, _27515_, _27468_);
  and _78139_ (_27517_, _27516_, _03600_);
  nor _78140_ (_27518_, _27517_, _27514_);
  nor _78141_ (_27519_, _27518_, _03780_);
  and _78142_ (_27520_, _12128_, _05300_);
  or _78143_ (_27521_, _27468_, _07778_);
  nor _78144_ (_27522_, _27521_, _27520_);
  or _78145_ (_27523_, _27522_, _03622_);
  nor _78146_ (_27524_, _27523_, _27519_);
  or _78147_ (_27525_, _27511_, _07777_);
  nor _78148_ (_27526_, _27525_, _27469_);
  nor _78149_ (_27527_, _27526_, _27524_);
  nor _78150_ (_27528_, _27527_, _03790_);
  and _78151_ (_27529_, _12005_, _05300_);
  or _78152_ (_27532_, _27529_, _27468_);
  and _78153_ (_27533_, _27532_, _03790_);
  or _78154_ (_27534_, _27533_, _27528_);
  and _78155_ (_27535_, _27534_, _07795_);
  nor _78156_ (_27536_, _12122_, _10706_);
  nor _78157_ (_27537_, _27536_, _27468_);
  nor _78158_ (_27538_, _27537_, _07795_);
  or _78159_ (_27539_, _27538_, _27535_);
  and _78160_ (_27540_, _27539_, _07793_);
  nor _78161_ (_27541_, _12003_, _10706_);
  nor _78162_ (_27543_, _27541_, _27468_);
  nor _78163_ (_27544_, _27543_, _07793_);
  nor _78164_ (_27545_, _27544_, _17166_);
  not _78165_ (_27546_, _27545_);
  nor _78166_ (_27547_, _27546_, _27540_);
  nor _78167_ (_27548_, _27547_, _27471_);
  and _78168_ (_27549_, _27548_, _43000_);
  nor _78169_ (_27550_, \oc8051_golden_model_1.SP [0], rst);
  nor _78170_ (_27551_, _27550_, _00000_);
  or _78171_ (_43606_, _27551_, _27549_);
  nor _78172_ (_27553_, _05300_, _03496_);
  and _78173_ (_27554_, _12213_, _05300_);
  nor _78174_ (_27555_, _27554_, _27553_);
  nor _78175_ (_27556_, _27555_, _03514_);
  nor _78176_ (_27557_, _10774_, _03496_);
  and _78177_ (_27558_, _03178_, _03496_);
  nor _78178_ (_27559_, _05300_, \oc8051_golden_model_1.SP [1]);
  and _78179_ (_27560_, _05300_, _03274_);
  nor _78180_ (_27561_, _27560_, _27559_);
  and _78181_ (_27562_, _27561_, _04409_);
  nor _78182_ (_27564_, _04409_, _03496_);
  or _78183_ (_27565_, _27564_, _27562_);
  and _78184_ (_27566_, _27565_, _04763_);
  and _78185_ (_27567_, _03980_, _03496_);
  or _78186_ (_27568_, _27567_, _27566_);
  and _78187_ (_27569_, _27568_, _04081_);
  nor _78188_ (_27570_, _27559_, _27554_);
  and _78189_ (_27571_, _27570_, _03610_);
  or _78190_ (_27572_, _27571_, _27569_);
  and _78191_ (_27573_, _27572_, _03230_);
  nor _78192_ (_27575_, _03230_, \oc8051_golden_model_1.SP [1]);
  or _78193_ (_27576_, _27575_, _03723_);
  or _78194_ (_27577_, _27576_, _27573_);
  nand _78195_ (_27578_, _03501_, _03723_);
  and _78196_ (_27579_, _27578_, _27577_);
  and _78197_ (_27580_, _27579_, _03737_);
  and _78198_ (_27581_, _27561_, _03729_);
  or _78199_ (_27582_, _27581_, _27580_);
  and _78200_ (_27583_, _27582_, _03510_);
  or _78201_ (_27584_, _27583_, _10694_);
  nor _78202_ (_27586_, _27584_, _03509_);
  nor _78203_ (_27587_, _04767_, _03496_);
  or _78204_ (_27588_, _27587_, _07390_);
  nor _78205_ (_27589_, _27588_, _27586_);
  or _78206_ (_27590_, _10706_, _06764_);
  nor _78207_ (_27591_, _27559_, _06838_);
  and _78208_ (_27592_, _27591_, _27590_);
  nor _78209_ (_27593_, _27592_, _04481_);
  not _78210_ (_27594_, _27593_);
  nor _78211_ (_27595_, _27594_, _27589_);
  and _78212_ (_27597_, _06501_, _05300_);
  nor _78213_ (_27598_, _27553_, _07400_);
  not _78214_ (_27599_, _27598_);
  nor _78215_ (_27600_, _27599_, _27597_);
  nor _78216_ (_27601_, _27600_, _03222_);
  not _78217_ (_27602_, _27601_);
  nor _78218_ (_27603_, _27602_, _27595_);
  nor _78219_ (_27604_, _12313_, _10706_);
  or _78220_ (_27605_, _27604_, _27553_);
  and _78221_ (_27606_, _27605_, _03222_);
  nor _78222_ (_27608_, _27606_, _27603_);
  nor _78223_ (_27609_, _27608_, _03601_);
  and _78224_ (_27610_, _05300_, _06282_);
  or _78225_ (_27611_, _27610_, _27553_);
  and _78226_ (_27612_, _27611_, _03601_);
  or _78227_ (_27613_, _27612_, _27609_);
  and _78228_ (_27614_, _27613_, _10736_);
  or _78229_ (_27615_, _27614_, _27558_);
  and _78230_ (_27616_, _27615_, _07766_);
  nor _78231_ (_27617_, _12327_, _10706_);
  or _78232_ (_27619_, _27617_, _07766_);
  nor _78233_ (_27620_, _27619_, _27559_);
  nor _78234_ (_27621_, _27620_, _27616_);
  nor _78235_ (_27622_, _27621_, _03780_);
  nor _78236_ (_27623_, _12333_, _10706_);
  or _78237_ (_27624_, _27623_, _07778_);
  nor _78238_ (_27625_, _27624_, _27559_);
  nor _78239_ (_27626_, _27625_, _27622_);
  nor _78240_ (_27627_, _27626_, _03622_);
  nor _78241_ (_27628_, _12207_, _10706_);
  or _78242_ (_27630_, _27628_, _07777_);
  nor _78243_ (_27631_, _27630_, _27559_);
  nor _78244_ (_27632_, _27631_, _27627_);
  nor _78245_ (_27633_, _27632_, _10754_);
  and _78246_ (_27634_, _03192_, _03496_);
  nor _78247_ (_27635_, _27553_, _05618_);
  nor _78248_ (_27636_, _27635_, _06828_);
  and _78249_ (_27637_, _27636_, _27561_);
  nor _78250_ (_27638_, _27637_, _27634_);
  not _78251_ (_27639_, _27638_);
  nor _78252_ (_27641_, _27639_, _27633_);
  or _78253_ (_27642_, _27641_, _18499_);
  nor _78254_ (_27643_, _12332_, _10706_);
  or _78255_ (_27644_, _27643_, _27553_);
  and _78256_ (_27645_, _27644_, _03785_);
  not _78257_ (_27646_, _10774_);
  nor _78258_ (_27647_, _12326_, _10706_);
  or _78259_ (_27648_, _27647_, _27553_);
  and _78260_ (_27649_, _27648_, _03624_);
  or _78261_ (_27650_, _27649_, _27646_);
  nor _78262_ (_27652_, _27650_, _27645_);
  and _78263_ (_27653_, _27652_, _27642_);
  nor _78264_ (_27654_, _27653_, _27557_);
  and _78265_ (_27655_, _27654_, _03516_);
  and _78266_ (_27656_, _03515_, _03496_);
  or _78267_ (_27657_, _27656_, _27655_);
  and _78268_ (_27658_, _27657_, _04246_);
  and _78269_ (_27659_, _27570_, _03815_);
  nor _78270_ (_27660_, _27659_, _05103_);
  not _78271_ (_27661_, _27660_);
  nor _78272_ (_27663_, _27661_, _27658_);
  nor _78273_ (_27664_, _04540_, _03496_);
  nor _78274_ (_27665_, _27664_, _03447_);
  not _78275_ (_27666_, _27665_);
  nor _78276_ (_27667_, _27666_, _27663_);
  nor _78277_ (_27668_, _27667_, _27556_);
  nor _78278_ (_27669_, _27668_, _43004_);
  nor _78279_ (_27670_, \oc8051_golden_model_1.SP [1], rst);
  nor _78280_ (_27671_, _27670_, _00000_);
  or _78281_ (_43607_, _27671_, _27669_);
  and _78282_ (_27673_, _05129_, _03188_);
  nor _78283_ (_27674_, _05300_, _03995_);
  and _78284_ (_27675_, _12539_, _05300_);
  nor _78285_ (_27676_, _27675_, _27674_);
  nor _78286_ (_27677_, _27676_, _07778_);
  and _78287_ (_27678_, _12192_, _03178_);
  not _78288_ (_27679_, _27674_);
  nor _78289_ (_27680_, _10706_, _04875_);
  nor _78290_ (_27681_, _27680_, _06838_);
  and _78291_ (_27682_, _27681_, _27679_);
  nor _78292_ (_27684_, _12416_, _10706_);
  nor _78293_ (_27685_, _27684_, _27674_);
  nor _78294_ (_27686_, _27685_, _04081_);
  nor _78295_ (_27687_, _04409_, _03995_);
  and _78296_ (_27688_, _05300_, \oc8051_golden_model_1.ACC [2]);
  nor _78297_ (_27689_, _27688_, _27674_);
  nor _78298_ (_27690_, _27689_, _09029_);
  nor _78299_ (_27691_, _27690_, _27687_);
  nor _78300_ (_27692_, _27691_, _03980_);
  and _78301_ (_27693_, _05129_, _03980_);
  nor _78302_ (_27695_, _27693_, _27692_);
  nor _78303_ (_27696_, _27695_, _03610_);
  or _78304_ (_27697_, _27696_, _04768_);
  nor _78305_ (_27698_, _27697_, _27686_);
  nor _78306_ (_27699_, _05129_, _03230_);
  or _78307_ (_27700_, _27699_, _03723_);
  nor _78308_ (_27701_, _27700_, _27698_);
  nor _78309_ (_27702_, _05984_, _03996_);
  or _78310_ (_27703_, _27702_, _27701_);
  and _78311_ (_27704_, _27703_, _03737_);
  nor _78312_ (_27706_, _27689_, _03737_);
  or _78313_ (_27707_, _27706_, _27704_);
  and _78314_ (_27708_, _27707_, _03510_);
  nor _78315_ (_27709_, _27708_, _04811_);
  nor _78316_ (_27710_, _27709_, _10694_);
  nor _78317_ (_27711_, _12192_, _04767_);
  nor _78318_ (_27712_, _27711_, _07390_);
  not _78319_ (_27713_, _27712_);
  nor _78320_ (_27714_, _27713_, _27710_);
  nor _78321_ (_27715_, _27714_, _27682_);
  nor _78322_ (_27717_, _27715_, _04481_);
  and _78323_ (_27718_, _06637_, _05300_);
  nor _78324_ (_27719_, _27674_, _07400_);
  not _78325_ (_27720_, _27719_);
  nor _78326_ (_27721_, _27720_, _27718_);
  or _78327_ (_27722_, _27721_, _03222_);
  nor _78328_ (_27723_, _27722_, _27717_);
  nor _78329_ (_27724_, _12519_, _10706_);
  nor _78330_ (_27725_, _27724_, _27674_);
  nor _78331_ (_27726_, _27725_, _03589_);
  or _78332_ (_27728_, _27726_, _03601_);
  or _78333_ (_27729_, _27728_, _27723_);
  and _78334_ (_27730_, _05300_, _06332_);
  nor _78335_ (_27731_, _27730_, _27674_);
  nand _78336_ (_27732_, _27731_, _03601_);
  and _78337_ (_27733_, _27732_, _27729_);
  nor _78338_ (_27734_, _27733_, _03178_);
  nor _78339_ (_27735_, _27734_, _27678_);
  nor _78340_ (_27736_, _27735_, _03600_);
  and _78341_ (_27737_, _12533_, _05300_);
  or _78342_ (_27739_, _27674_, _07766_);
  nor _78343_ (_27740_, _27739_, _27737_);
  or _78344_ (_27741_, _27740_, _03780_);
  nor _78345_ (_27742_, _27741_, _27736_);
  nor _78346_ (_27743_, _27742_, _27677_);
  nor _78347_ (_27744_, _27743_, _03622_);
  and _78348_ (_27745_, _27679_, _05717_);
  not _78349_ (_27746_, _27745_);
  nor _78350_ (_27747_, _27731_, _07777_);
  and _78351_ (_27748_, _27747_, _27746_);
  nor _78352_ (_27750_, _27748_, _27744_);
  nor _78353_ (_27751_, _27750_, _10754_);
  nor _78354_ (_27752_, _27689_, _06828_);
  and _78355_ (_27753_, _27752_, _27746_);
  and _78356_ (_27754_, _05129_, _03192_);
  nor _78357_ (_27755_, _27754_, _27753_);
  and _78358_ (_27756_, _27755_, _07795_);
  not _78359_ (_27757_, _27756_);
  nor _78360_ (_27758_, _27757_, _27751_);
  nor _78361_ (_27759_, _12532_, _10706_);
  nor _78362_ (_27761_, _27759_, _27674_);
  and _78363_ (_27762_, _27761_, _03624_);
  nor _78364_ (_27763_, _27762_, _27758_);
  nor _78365_ (_27764_, _27763_, _03785_);
  nor _78366_ (_27765_, _12538_, _10706_);
  or _78367_ (_27766_, _27674_, _07793_);
  nor _78368_ (_27767_, _27766_, _27765_);
  or _78369_ (_27768_, _27767_, _03798_);
  nor _78370_ (_27769_, _27768_, _27764_);
  and _78371_ (_27770_, _12192_, _03798_);
  or _78372_ (_27772_, _27770_, _27769_);
  and _78373_ (_27773_, _27772_, _06399_);
  or _78374_ (_27774_, _27773_, _27673_);
  and _78375_ (_27775_, _27774_, _03516_);
  and _78376_ (_27776_, _12192_, _03515_);
  or _78377_ (_27777_, _27776_, _03815_);
  nor _78378_ (_27778_, _27777_, _27775_);
  and _78379_ (_27779_, _27685_, _03815_);
  or _78380_ (_27780_, _27779_, _05103_);
  nor _78381_ (_27781_, _27780_, _27778_);
  nor _78382_ (_27783_, _12192_, _04540_);
  nor _78383_ (_27784_, _27783_, _03447_);
  not _78384_ (_27785_, _27784_);
  nor _78385_ (_27786_, _27785_, _27781_);
  and _78386_ (_27787_, _12592_, _05300_);
  nor _78387_ (_27788_, _27787_, _27674_);
  and _78388_ (_27789_, _27788_, _03447_);
  nor _78389_ (_27790_, _27789_, _27786_);
  and _78390_ (_27791_, _27790_, _43000_);
  nor _78391_ (_27792_, \oc8051_golden_model_1.SP [2], rst);
  nor _78392_ (_27794_, _27792_, _00000_);
  or _78393_ (_43608_, _27794_, _27791_);
  nor _78394_ (_27795_, _05133_, _04540_);
  and _78395_ (_27796_, _05133_, _03188_);
  and _78396_ (_27797_, _05133_, _03192_);
  nor _78397_ (_27798_, _27797_, _03624_);
  nor _78398_ (_27799_, _05300_, _03722_);
  and _78399_ (_27800_, _12739_, _05300_);
  nor _78400_ (_27801_, _27800_, _27799_);
  nor _78401_ (_27802_, _27801_, _07778_);
  and _78402_ (_27803_, _05132_, _03178_);
  nor _78403_ (_27804_, _04409_, _03722_);
  and _78404_ (_27805_, _05300_, \oc8051_golden_model_1.ACC [3]);
  nor _78405_ (_27806_, _27805_, _27799_);
  nor _78406_ (_27807_, _27806_, _09029_);
  or _78407_ (_27808_, _27807_, _27804_);
  and _78408_ (_27809_, _27808_, _04763_);
  and _78409_ (_27810_, _05133_, _03980_);
  nor _78410_ (_27811_, _27810_, _27809_);
  nor _78411_ (_27812_, _27811_, _03610_);
  nor _78412_ (_27815_, _12627_, _10706_);
  nor _78413_ (_27816_, _27815_, _27799_);
  nor _78414_ (_27817_, _27816_, _04081_);
  or _78415_ (_27818_, _27817_, _27812_);
  and _78416_ (_27819_, _27818_, _03230_);
  nor _78417_ (_27820_, _05132_, _03230_);
  or _78418_ (_27821_, _27820_, _03723_);
  or _78419_ (_27822_, _27821_, _27819_);
  nand _78420_ (_27823_, _05973_, _03723_);
  and _78421_ (_27824_, _27823_, _27822_);
  and _78422_ (_27826_, _27824_, _03737_);
  nor _78423_ (_27827_, _27806_, _03737_);
  or _78424_ (_27828_, _27827_, _27826_);
  and _78425_ (_27829_, _27828_, _03510_);
  or _78426_ (_27830_, _27829_, _10694_);
  nor _78427_ (_27831_, _27830_, _05053_);
  nor _78428_ (_27832_, _05133_, _04767_);
  or _78429_ (_27833_, _27832_, _07390_);
  nor _78430_ (_27834_, _27833_, _27831_);
  nor _78431_ (_27835_, _10706_, _05005_);
  nor _78432_ (_27837_, _27835_, _27799_);
  nor _78433_ (_27838_, _27837_, _06838_);
  nor _78434_ (_27839_, _27838_, _04481_);
  not _78435_ (_27840_, _27839_);
  nor _78436_ (_27841_, _27840_, _27834_);
  and _78437_ (_27842_, _06592_, _05300_);
  nor _78438_ (_27843_, _27799_, _07400_);
  not _78439_ (_27844_, _27843_);
  nor _78440_ (_27845_, _27844_, _27842_);
  or _78441_ (_27846_, _27845_, _03222_);
  nor _78442_ (_27848_, _27846_, _27841_);
  nor _78443_ (_27849_, _12718_, _10706_);
  nor _78444_ (_27850_, _27849_, _27799_);
  nor _78445_ (_27851_, _27850_, _03589_);
  or _78446_ (_27852_, _27851_, _03601_);
  or _78447_ (_27853_, _27852_, _27848_);
  and _78448_ (_27854_, _05300_, _06276_);
  nor _78449_ (_27855_, _27854_, _27799_);
  nand _78450_ (_27856_, _27855_, _03601_);
  and _78451_ (_27857_, _27856_, _27853_);
  nor _78452_ (_27859_, _27857_, _03178_);
  nor _78453_ (_27860_, _27859_, _27803_);
  nor _78454_ (_27861_, _27860_, _03600_);
  and _78455_ (_27862_, _12733_, _05300_);
  or _78456_ (_27863_, _27799_, _07766_);
  nor _78457_ (_27864_, _27863_, _27862_);
  or _78458_ (_27865_, _27864_, _03780_);
  nor _78459_ (_27866_, _27865_, _27861_);
  nor _78460_ (_27867_, _27866_, _27802_);
  nor _78461_ (_27868_, _27867_, _03622_);
  nor _78462_ (_27870_, _27799_, _05567_);
  not _78463_ (_27871_, _27870_);
  nor _78464_ (_27872_, _27855_, _07777_);
  and _78465_ (_27873_, _27872_, _27871_);
  nor _78466_ (_27874_, _27873_, _27868_);
  nor _78467_ (_27875_, _27874_, _10754_);
  nor _78468_ (_27876_, _27806_, _06828_);
  and _78469_ (_27877_, _27876_, _27871_);
  nor _78470_ (_27878_, _27877_, _27875_);
  and _78471_ (_27879_, _27878_, _27798_);
  nor _78472_ (_27881_, _12732_, _10706_);
  nor _78473_ (_27882_, _27881_, _27799_);
  and _78474_ (_27883_, _27882_, _03624_);
  nor _78475_ (_27884_, _27883_, _27879_);
  nor _78476_ (_27885_, _27884_, _03785_);
  nor _78477_ (_27886_, _12738_, _10706_);
  or _78478_ (_27887_, _27799_, _07793_);
  nor _78479_ (_27888_, _27887_, _27886_);
  or _78480_ (_27889_, _27888_, _03798_);
  nor _78481_ (_27890_, _27889_, _27885_);
  nor _78482_ (_27892_, _05970_, _03722_);
  nor _78483_ (_27893_, _27892_, _05971_);
  nor _78484_ (_27894_, _27893_, _10652_);
  or _78485_ (_27895_, _27894_, _27890_);
  and _78486_ (_27896_, _27895_, _06399_);
  or _78487_ (_27897_, _27896_, _27796_);
  and _78488_ (_27898_, _27897_, _03516_);
  nor _78489_ (_27899_, _27893_, _03516_);
  or _78490_ (_27900_, _27899_, _27898_);
  and _78491_ (_27901_, _27900_, _04246_);
  nor _78492_ (_27903_, _27816_, _04246_);
  nor _78493_ (_27904_, _27903_, _05103_);
  not _78494_ (_27905_, _27904_);
  nor _78495_ (_27906_, _27905_, _27901_);
  nor _78496_ (_27907_, _27906_, _27795_);
  and _78497_ (_27908_, _27907_, _03514_);
  and _78498_ (_27909_, _12794_, _05300_);
  nor _78499_ (_27910_, _27909_, _27799_);
  nor _78500_ (_27911_, _27910_, _03514_);
  or _78501_ (_27912_, _27911_, _27908_);
  or _78502_ (_27914_, _27912_, _43004_);
  or _78503_ (_27915_, _43000_, \oc8051_golden_model_1.SP [3]);
  and _78504_ (_27916_, _27915_, _41806_);
  and _78505_ (_43609_, _27916_, _27914_);
  nor _78506_ (_27917_, _05010_, \oc8051_golden_model_1.SP [4]);
  nor _78507_ (_27918_, _27917_, _10645_);
  nor _78508_ (_27919_, _27918_, _04540_);
  and _78509_ (_27920_, _27918_, _03192_);
  nor _78510_ (_27921_, _27920_, _03624_);
  nor _78511_ (_27922_, _05300_, _10679_);
  and _78512_ (_27924_, _12817_, _05300_);
  nor _78513_ (_27925_, _27924_, _27922_);
  nor _78514_ (_27926_, _27925_, _07778_);
  and _78515_ (_27927_, _05011_, \oc8051_golden_model_1.SP [4]);
  nor _78516_ (_27928_, _05011_, \oc8051_golden_model_1.SP [4]);
  nor _78517_ (_27929_, _27928_, _27927_);
  and _78518_ (_27930_, _27929_, _03508_);
  nor _78519_ (_27931_, _04409_, _10679_);
  and _78520_ (_27932_, _05300_, \oc8051_golden_model_1.ACC [4]);
  nor _78521_ (_27933_, _27932_, _27922_);
  nor _78522_ (_27935_, _27933_, _09029_);
  or _78523_ (_27936_, _27935_, _27931_);
  and _78524_ (_27937_, _27936_, _04763_);
  and _78525_ (_27938_, _27918_, _03980_);
  nor _78526_ (_27939_, _27938_, _27937_);
  nor _78527_ (_27940_, _27939_, _03610_);
  nor _78528_ (_27941_, _12841_, _10706_);
  nor _78529_ (_27942_, _27941_, _27922_);
  nor _78530_ (_27943_, _27942_, _04081_);
  or _78531_ (_27944_, _27943_, _27940_);
  and _78532_ (_27946_, _27944_, _03230_);
  and _78533_ (_27947_, _27918_, _04768_);
  or _78534_ (_27948_, _27947_, _27946_);
  and _78535_ (_27949_, _27948_, _03996_);
  and _78536_ (_27950_, _10680_, _03498_);
  nor _78537_ (_27951_, _05972_, _10679_);
  nor _78538_ (_27952_, _27951_, _27950_);
  nor _78539_ (_27953_, _27952_, _03996_);
  or _78540_ (_27954_, _27953_, _27949_);
  and _78541_ (_27955_, _27954_, _03737_);
  nor _78542_ (_27957_, _27933_, _03737_);
  or _78543_ (_27958_, _27957_, _27955_);
  and _78544_ (_27959_, _27958_, _03510_);
  or _78545_ (_27960_, _27959_, _10694_);
  nor _78546_ (_27961_, _27960_, _27930_);
  nor _78547_ (_27962_, _27918_, _04767_);
  or _78548_ (_27963_, _27962_, _07390_);
  nor _78549_ (_27964_, _27963_, _27961_);
  nor _78550_ (_27965_, _05777_, _10706_);
  nor _78551_ (_27966_, _27965_, _27922_);
  nor _78552_ (_27968_, _27966_, _06838_);
  nor _78553_ (_27969_, _27968_, _04481_);
  not _78554_ (_27970_, _27969_);
  nor _78555_ (_27971_, _27970_, _27964_);
  and _78556_ (_27972_, _06730_, _05300_);
  nor _78557_ (_27973_, _27922_, _07400_);
  not _78558_ (_27974_, _27973_);
  nor _78559_ (_27975_, _27974_, _27972_);
  nor _78560_ (_27976_, _27975_, _03222_);
  not _78561_ (_27977_, _27976_);
  nor _78562_ (_27979_, _27977_, _27971_);
  nor _78563_ (_27980_, _12933_, _10706_);
  nor _78564_ (_27981_, _27980_, _27922_);
  nor _78565_ (_27982_, _27981_, _03589_);
  or _78566_ (_27983_, _27982_, _27979_);
  and _78567_ (_27984_, _27983_, _05886_);
  and _78568_ (_27985_, _06298_, _05300_);
  nor _78569_ (_27986_, _27985_, _27922_);
  nor _78570_ (_27987_, _27986_, _05886_);
  or _78571_ (_27988_, _27987_, _27984_);
  and _78572_ (_27990_, _27988_, _10736_);
  and _78573_ (_27991_, _27918_, _03178_);
  or _78574_ (_27992_, _27991_, _03600_);
  nor _78575_ (_27993_, _27992_, _27990_);
  and _78576_ (_27994_, _12821_, _05300_);
  or _78577_ (_27995_, _27922_, _07766_);
  nor _78578_ (_27996_, _27995_, _27994_);
  or _78579_ (_27997_, _27996_, _03780_);
  nor _78580_ (_27998_, _27997_, _27993_);
  nor _78581_ (_27999_, _27998_, _27926_);
  nor _78582_ (_28001_, _27999_, _03622_);
  nor _78583_ (_28002_, _27922_, _05825_);
  not _78584_ (_28003_, _28002_);
  nor _78585_ (_28004_, _27986_, _07777_);
  and _78586_ (_28005_, _28004_, _28003_);
  nor _78587_ (_28006_, _28005_, _28001_);
  nor _78588_ (_28007_, _28006_, _10754_);
  nor _78589_ (_28008_, _27933_, _06828_);
  and _78590_ (_28009_, _28008_, _28003_);
  nor _78591_ (_28010_, _28009_, _28007_);
  and _78592_ (_28012_, _28010_, _27921_);
  nor _78593_ (_28013_, _12819_, _10706_);
  nor _78594_ (_28014_, _28013_, _27922_);
  and _78595_ (_28015_, _28014_, _03624_);
  nor _78596_ (_28016_, _28015_, _28012_);
  nor _78597_ (_28017_, _28016_, _03785_);
  nor _78598_ (_28018_, _12816_, _10706_);
  or _78599_ (_28019_, _27922_, _07793_);
  nor _78600_ (_28020_, _28019_, _28018_);
  or _78601_ (_28021_, _28020_, _03798_);
  nor _78602_ (_28023_, _28021_, _28017_);
  nor _78603_ (_28024_, _05971_, _10679_);
  nor _78604_ (_28025_, _28024_, _10680_);
  nor _78605_ (_28026_, _28025_, _10652_);
  or _78606_ (_28027_, _28026_, _28023_);
  and _78607_ (_28028_, _28027_, _06399_);
  and _78608_ (_28029_, _27918_, _03188_);
  or _78609_ (_28030_, _28029_, _28028_);
  and _78610_ (_28031_, _28030_, _03516_);
  nor _78611_ (_28032_, _28025_, _03516_);
  or _78612_ (_28034_, _28032_, _28031_);
  and _78613_ (_28035_, _28034_, _04246_);
  nor _78614_ (_28036_, _27942_, _04246_);
  nor _78615_ (_28037_, _28036_, _05103_);
  not _78616_ (_28038_, _28037_);
  nor _78617_ (_28039_, _28038_, _28035_);
  nor _78618_ (_28040_, _28039_, _27919_);
  and _78619_ (_28041_, _28040_, _03514_);
  and _78620_ (_28042_, _13003_, _05300_);
  nor _78621_ (_28043_, _28042_, _27922_);
  nor _78622_ (_28045_, _28043_, _03514_);
  or _78623_ (_28046_, _28045_, _28041_);
  or _78624_ (_28047_, _28046_, _43004_);
  or _78625_ (_28048_, _43000_, \oc8051_golden_model_1.SP [4]);
  and _78626_ (_28049_, _28048_, _41806_);
  and _78627_ (_43610_, _28049_, _28047_);
  nor _78628_ (_28050_, _10645_, \oc8051_golden_model_1.SP [5]);
  nor _78629_ (_28051_, _28050_, _10646_);
  nor _78630_ (_28052_, _28051_, _04540_);
  nor _78631_ (_28053_, _05300_, _10678_);
  and _78632_ (_28055_, _13147_, _05300_);
  nor _78633_ (_28056_, _28055_, _28053_);
  nor _78634_ (_28057_, _28056_, _07778_);
  nor _78635_ (_28058_, _04409_, _10678_);
  and _78636_ (_28059_, _05300_, \oc8051_golden_model_1.ACC [5]);
  nor _78637_ (_28060_, _28059_, _28053_);
  nor _78638_ (_28061_, _28060_, _09029_);
  or _78639_ (_28062_, _28061_, _28058_);
  and _78640_ (_28063_, _28062_, _04763_);
  and _78641_ (_28064_, _28051_, _03980_);
  nor _78642_ (_28066_, _28064_, _28063_);
  nor _78643_ (_28067_, _28066_, _03610_);
  nor _78644_ (_28068_, _13014_, _10706_);
  nor _78645_ (_28069_, _28068_, _28053_);
  nor _78646_ (_28070_, _28069_, _04081_);
  or _78647_ (_28071_, _28070_, _28067_);
  and _78648_ (_28072_, _28071_, _03230_);
  and _78649_ (_28073_, _28051_, _04768_);
  or _78650_ (_28074_, _28073_, _28072_);
  and _78651_ (_28075_, _28074_, _03996_);
  and _78652_ (_28077_, _10681_, _03498_);
  nor _78653_ (_28078_, _27950_, _10678_);
  nor _78654_ (_28079_, _28078_, _28077_);
  nor _78655_ (_28080_, _28079_, _03996_);
  or _78656_ (_28081_, _28080_, _28075_);
  and _78657_ (_28082_, _28081_, _03737_);
  nor _78658_ (_28083_, _28060_, _03737_);
  or _78659_ (_28084_, _28083_, _28082_);
  and _78660_ (_28085_, _28084_, _03510_);
  and _78661_ (_28086_, _10646_, \oc8051_golden_model_1.SP [0]);
  nor _78662_ (_28088_, _27927_, \oc8051_golden_model_1.SP [5]);
  nor _78663_ (_28089_, _28088_, _28086_);
  and _78664_ (_28090_, _28089_, _03508_);
  nor _78665_ (_28091_, _28090_, _10694_);
  not _78666_ (_28092_, _28091_);
  nor _78667_ (_28093_, _28092_, _28085_);
  nor _78668_ (_28094_, _28051_, _04767_);
  or _78669_ (_28095_, _28094_, _07390_);
  nor _78670_ (_28096_, _28095_, _28093_);
  nor _78671_ (_28097_, _05469_, _10706_);
  nor _78672_ (_28099_, _28097_, _28053_);
  nor _78673_ (_28100_, _28099_, _06838_);
  nor _78674_ (_28101_, _28100_, _04481_);
  not _78675_ (_28102_, _28101_);
  nor _78676_ (_28103_, _28102_, _28096_);
  and _78677_ (_28104_, _06684_, _05300_);
  nor _78678_ (_28105_, _28053_, _07400_);
  not _78679_ (_28106_, _28105_);
  nor _78680_ (_28107_, _28106_, _28104_);
  nor _78681_ (_28108_, _28107_, _03222_);
  not _78682_ (_28110_, _28108_);
  nor _78683_ (_28111_, _28110_, _28103_);
  nor _78684_ (_28112_, _13127_, _10706_);
  nor _78685_ (_28113_, _28112_, _28053_);
  nor _78686_ (_28114_, _28113_, _03589_);
  or _78687_ (_28115_, _28114_, _28111_);
  and _78688_ (_28116_, _28115_, _05886_);
  and _78689_ (_28117_, _06306_, _05300_);
  nor _78690_ (_28118_, _28117_, _28053_);
  nor _78691_ (_28119_, _28118_, _05886_);
  or _78692_ (_28121_, _28119_, _28116_);
  and _78693_ (_28122_, _28121_, _10736_);
  and _78694_ (_28123_, _28051_, _03178_);
  or _78695_ (_28124_, _28123_, _03600_);
  nor _78696_ (_28125_, _28124_, _28122_);
  and _78697_ (_28126_, _13141_, _05300_);
  or _78698_ (_28127_, _28053_, _07766_);
  nor _78699_ (_28128_, _28127_, _28126_);
  or _78700_ (_28129_, _28128_, _03780_);
  nor _78701_ (_28130_, _28129_, _28125_);
  nor _78702_ (_28132_, _28130_, _28057_);
  nor _78703_ (_28133_, _28132_, _03622_);
  nor _78704_ (_28134_, _28053_, _05518_);
  not _78705_ (_28135_, _28134_);
  nor _78706_ (_28136_, _28118_, _07777_);
  and _78707_ (_28137_, _28136_, _28135_);
  nor _78708_ (_28138_, _28137_, _28133_);
  nor _78709_ (_28139_, _28138_, _10754_);
  nor _78710_ (_28140_, _28060_, _06828_);
  and _78711_ (_28141_, _28140_, _28135_);
  and _78712_ (_28143_, _28051_, _03192_);
  nor _78713_ (_28144_, _28143_, _28141_);
  and _78714_ (_28145_, _28144_, _07795_);
  not _78715_ (_28146_, _28145_);
  nor _78716_ (_28147_, _28146_, _28139_);
  nor _78717_ (_28148_, _13140_, _10706_);
  nor _78718_ (_28149_, _28148_, _28053_);
  and _78719_ (_28150_, _28149_, _03624_);
  nor _78720_ (_28151_, _28150_, _28147_);
  nor _78721_ (_28152_, _28151_, _03785_);
  nor _78722_ (_28154_, _13146_, _10706_);
  or _78723_ (_28155_, _28053_, _07793_);
  nor _78724_ (_28156_, _28155_, _28154_);
  or _78725_ (_28157_, _28156_, _03798_);
  nor _78726_ (_28158_, _28157_, _28152_);
  nor _78727_ (_28159_, _10680_, _10678_);
  nor _78728_ (_28160_, _28159_, _10681_);
  nor _78729_ (_28161_, _28160_, _10652_);
  or _78730_ (_28162_, _28161_, _28158_);
  and _78731_ (_28163_, _28162_, _06399_);
  and _78732_ (_28165_, _28051_, _03188_);
  or _78733_ (_28166_, _28165_, _28163_);
  and _78734_ (_28167_, _28166_, _03516_);
  nor _78735_ (_28168_, _28160_, _03516_);
  or _78736_ (_28169_, _28168_, _28167_);
  and _78737_ (_28170_, _28169_, _04246_);
  nor _78738_ (_28171_, _28069_, _04246_);
  nor _78739_ (_28172_, _28171_, _05103_);
  not _78740_ (_28173_, _28172_);
  nor _78741_ (_28174_, _28173_, _28170_);
  nor _78742_ (_28176_, _28174_, _28052_);
  nor _78743_ (_28177_, _28176_, _03447_);
  and _78744_ (_28178_, _13199_, _05300_);
  nor _78745_ (_28179_, _28178_, _28053_);
  and _78746_ (_28180_, _28179_, _03447_);
  nor _78747_ (_28181_, _28180_, _28177_);
  or _78748_ (_28182_, _28181_, _43004_);
  or _78749_ (_28183_, _43000_, \oc8051_golden_model_1.SP [5]);
  and _78750_ (_28184_, _28183_, _41806_);
  and _78751_ (_43611_, _28184_, _28182_);
  nor _78752_ (_28186_, _05300_, _10677_);
  and _78753_ (_28187_, _13353_, _05300_);
  nor _78754_ (_28188_, _28187_, _28186_);
  nor _78755_ (_28189_, _28188_, _07778_);
  and _78756_ (_28190_, _06455_, _05300_);
  or _78757_ (_28191_, _28190_, _28186_);
  and _78758_ (_28192_, _28191_, _04481_);
  and _78759_ (_28193_, _05300_, \oc8051_golden_model_1.ACC [6]);
  nor _78760_ (_28194_, _28193_, _28186_);
  nor _78761_ (_28195_, _28194_, _09029_);
  nor _78762_ (_28197_, _04409_, _10677_);
  or _78763_ (_28198_, _28197_, _03980_);
  nor _78764_ (_28199_, _28198_, _28195_);
  nor _78765_ (_28200_, _10646_, \oc8051_golden_model_1.SP [6]);
  nor _78766_ (_28201_, _28200_, _10647_);
  not _78767_ (_28202_, _28201_);
  and _78768_ (_28203_, _28202_, _03980_);
  nor _78769_ (_28204_, _28203_, _28199_);
  and _78770_ (_28205_, _28204_, _04081_);
  nor _78771_ (_28206_, _13242_, _10706_);
  nor _78772_ (_28208_, _28206_, _28186_);
  nor _78773_ (_28209_, _28208_, _04081_);
  or _78774_ (_28210_, _28209_, _28205_);
  and _78775_ (_28211_, _28210_, _03230_);
  nor _78776_ (_28212_, _28202_, _03230_);
  or _78777_ (_28213_, _28212_, _28211_);
  and _78778_ (_28214_, _28213_, _03996_);
  nor _78779_ (_28215_, _28077_, _10677_);
  nor _78780_ (_28216_, _28215_, _10683_);
  nor _78781_ (_28217_, _28216_, _03996_);
  or _78782_ (_28219_, _28217_, _28214_);
  and _78783_ (_28220_, _28219_, _03737_);
  nor _78784_ (_28221_, _28194_, _03737_);
  or _78785_ (_28222_, _28221_, _28220_);
  and _78786_ (_28223_, _28222_, _03510_);
  nor _78787_ (_28224_, _28086_, \oc8051_golden_model_1.SP [6]);
  nor _78788_ (_28225_, _28224_, _10695_);
  and _78789_ (_28226_, _28225_, _03508_);
  nor _78790_ (_28227_, _28226_, _28223_);
  nor _78791_ (_28228_, _28227_, _10694_);
  nor _78792_ (_28230_, _28202_, _04767_);
  nor _78793_ (_28231_, _28230_, _07390_);
  not _78794_ (_28232_, _28231_);
  nor _78795_ (_28233_, _28232_, _28228_);
  not _78796_ (_28234_, _28186_);
  nor _78797_ (_28235_, _05363_, _10706_);
  nor _78798_ (_28236_, _28235_, _06838_);
  and _78799_ (_28237_, _28236_, _28234_);
  or _78800_ (_28238_, _28237_, _04481_);
  nor _78801_ (_28239_, _28238_, _28233_);
  or _78802_ (_28240_, _28239_, _28192_);
  and _78803_ (_28241_, _28240_, _03589_);
  nor _78804_ (_28242_, _13332_, _10706_);
  nor _78805_ (_28243_, _28242_, _28186_);
  nor _78806_ (_28244_, _28243_, _03589_);
  or _78807_ (_28245_, _28244_, _03601_);
  or _78808_ (_28246_, _28245_, _28241_);
  and _78809_ (_28247_, _13339_, _05300_);
  nor _78810_ (_28248_, _28247_, _28186_);
  nand _78811_ (_28249_, _28248_, _03601_);
  and _78812_ (_28252_, _28249_, _28246_);
  nor _78813_ (_28253_, _28252_, _03178_);
  and _78814_ (_28254_, _28202_, _03178_);
  nor _78815_ (_28255_, _28254_, _28253_);
  nor _78816_ (_28256_, _28255_, _03600_);
  and _78817_ (_28257_, _13347_, _05300_);
  or _78818_ (_28258_, _28186_, _07766_);
  nor _78819_ (_28259_, _28258_, _28257_);
  or _78820_ (_28260_, _28259_, _03780_);
  nor _78821_ (_28261_, _28260_, _28256_);
  nor _78822_ (_28263_, _28261_, _28189_);
  nor _78823_ (_28264_, _28263_, _03622_);
  and _78824_ (_28265_, _28234_, _05411_);
  not _78825_ (_28266_, _28265_);
  nor _78826_ (_28267_, _28248_, _07777_);
  and _78827_ (_28268_, _28267_, _28266_);
  nor _78828_ (_28269_, _28268_, _28264_);
  nor _78829_ (_28270_, _28269_, _10754_);
  and _78830_ (_28271_, _28201_, _03192_);
  or _78831_ (_28272_, _28265_, _06828_);
  nor _78832_ (_28274_, _28272_, _28194_);
  nor _78833_ (_28275_, _28274_, _28271_);
  and _78834_ (_28276_, _28275_, _07795_);
  not _78835_ (_28277_, _28276_);
  nor _78836_ (_28278_, _28277_, _28270_);
  nor _78837_ (_28279_, _13346_, _10706_);
  nor _78838_ (_28280_, _28279_, _28186_);
  and _78839_ (_28281_, _28280_, _03624_);
  nor _78840_ (_28282_, _28281_, _28278_);
  and _78841_ (_28283_, _28282_, _07793_);
  nor _78842_ (_28285_, _13352_, _10706_);
  nor _78843_ (_28286_, _28285_, _28186_);
  nor _78844_ (_28287_, _28286_, _07793_);
  or _78845_ (_28288_, _28287_, _28283_);
  and _78846_ (_28289_, _28288_, _10652_);
  nor _78847_ (_28290_, _10681_, _10677_);
  nor _78848_ (_28291_, _28290_, _10682_);
  not _78849_ (_28292_, _28291_);
  nor _78850_ (_28293_, _28292_, _03188_);
  nor _78851_ (_28294_, _28293_, _10774_);
  nor _78852_ (_28296_, _28294_, _28289_);
  and _78853_ (_28297_, _28202_, _03188_);
  or _78854_ (_28298_, _28297_, _03515_);
  nor _78855_ (_28299_, _28298_, _28296_);
  and _78856_ (_28300_, _28292_, _03515_);
  or _78857_ (_28301_, _28300_, _03815_);
  nor _78858_ (_28302_, _28301_, _28299_);
  and _78859_ (_28303_, _28208_, _03815_);
  nor _78860_ (_28304_, _28303_, _05103_);
  not _78861_ (_28305_, _28304_);
  nor _78862_ (_28307_, _28305_, _28302_);
  nor _78863_ (_28308_, _28202_, _04540_);
  nor _78864_ (_28309_, _28308_, _03447_);
  not _78865_ (_28310_, _28309_);
  nor _78866_ (_28311_, _28310_, _28307_);
  and _78867_ (_28312_, _13402_, _05300_);
  or _78868_ (_28313_, _28186_, _03514_);
  nor _78869_ (_28314_, _28313_, _28312_);
  nor _78870_ (_28315_, _28314_, _28311_);
  or _78871_ (_28316_, _28315_, _43004_);
  or _78872_ (_28318_, _43000_, \oc8051_golden_model_1.SP [6]);
  and _78873_ (_28319_, _28318_, _41806_);
  and _78874_ (_43612_, _28319_, _28316_);
  not _78875_ (_28320_, \oc8051_golden_model_1.TCON [0]);
  nor _78876_ (_28321_, _05258_, _28320_);
  and _78877_ (_28322_, _12128_, _05258_);
  nor _78878_ (_28323_, _28322_, _28321_);
  nor _78879_ (_28324_, _28323_, _07778_);
  and _78880_ (_28325_, _05258_, _06274_);
  nor _78881_ (_28326_, _28325_, _28321_);
  and _78882_ (_28328_, _28326_, _03601_);
  and _78883_ (_28329_, _05258_, _04620_);
  nor _78884_ (_28330_, _28329_, _28321_);
  and _78885_ (_28331_, _28330_, _07390_);
  and _78886_ (_28332_, _05258_, \oc8051_golden_model_1.ACC [0]);
  nor _78887_ (_28333_, _28332_, _28321_);
  nor _78888_ (_28334_, _28333_, _09029_);
  nor _78889_ (_28335_, _04409_, _28320_);
  or _78890_ (_28336_, _28335_, _28334_);
  and _78891_ (_28337_, _28336_, _04081_);
  nor _78892_ (_28339_, _05666_, _10802_);
  nor _78893_ (_28340_, _28339_, _28321_);
  nor _78894_ (_28341_, _28340_, _04081_);
  or _78895_ (_28342_, _28341_, _28337_);
  and _78896_ (_28343_, _28342_, _04055_);
  nor _78897_ (_28344_, _05927_, _28320_);
  and _78898_ (_28345_, _12021_, _05927_);
  nor _78899_ (_28346_, _28345_, _28344_);
  nor _78900_ (_28347_, _28346_, _04055_);
  nor _78901_ (_28348_, _28347_, _28343_);
  nor _78902_ (_28350_, _28348_, _03723_);
  nor _78903_ (_28351_, _28330_, _03996_);
  or _78904_ (_28352_, _28351_, _28350_);
  and _78905_ (_28353_, _28352_, _03737_);
  nor _78906_ (_28354_, _28333_, _03737_);
  or _78907_ (_28355_, _28354_, _28353_);
  and _78908_ (_28356_, _28355_, _03736_);
  and _78909_ (_28357_, _28321_, _03714_);
  or _78910_ (_28358_, _28357_, _28356_);
  and _78911_ (_28359_, _28358_, _06840_);
  nor _78912_ (_28361_, _28340_, _06840_);
  or _78913_ (_28362_, _28361_, _28359_);
  and _78914_ (_28363_, _28362_, _03710_);
  nor _78915_ (_28364_, _12052_, _10839_);
  nor _78916_ (_28365_, _28364_, _28344_);
  nor _78917_ (_28366_, _28365_, _03710_);
  or _78918_ (_28367_, _28366_, _07390_);
  nor _78919_ (_28368_, _28367_, _28363_);
  nor _78920_ (_28369_, _28368_, _28331_);
  nor _78921_ (_28370_, _28369_, _04481_);
  and _78922_ (_28372_, _06546_, _05258_);
  nor _78923_ (_28373_, _28321_, _07400_);
  not _78924_ (_28374_, _28373_);
  nor _78925_ (_28375_, _28374_, _28372_);
  or _78926_ (_28376_, _28375_, _03222_);
  nor _78927_ (_28377_, _28376_, _28370_);
  nor _78928_ (_28378_, _12109_, _10802_);
  nor _78929_ (_28379_, _28378_, _28321_);
  nor _78930_ (_28380_, _28379_, _03589_);
  or _78931_ (_28381_, _28380_, _03601_);
  nor _78932_ (_28383_, _28381_, _28377_);
  nor _78933_ (_28384_, _28383_, _28328_);
  or _78934_ (_28385_, _28384_, _03600_);
  and _78935_ (_28386_, _12124_, _05258_);
  or _78936_ (_28387_, _28386_, _28321_);
  or _78937_ (_28388_, _28387_, _07766_);
  and _78938_ (_28389_, _28388_, _07778_);
  and _78939_ (_28390_, _28389_, _28385_);
  nor _78940_ (_28391_, _28390_, _28324_);
  nor _78941_ (_28392_, _28391_, _03622_);
  or _78942_ (_28394_, _28326_, _07777_);
  nor _78943_ (_28395_, _28394_, _28339_);
  nor _78944_ (_28396_, _28395_, _28392_);
  nor _78945_ (_28397_, _28396_, _03790_);
  and _78946_ (_28398_, _12005_, _05258_);
  or _78947_ (_28399_, _28398_, _28321_);
  and _78948_ (_28400_, _28399_, _03790_);
  or _78949_ (_28401_, _28400_, _28397_);
  and _78950_ (_28402_, _28401_, _07795_);
  nor _78951_ (_28403_, _12122_, _10802_);
  nor _78952_ (_28405_, _28403_, _28321_);
  nor _78953_ (_28406_, _28405_, _07795_);
  or _78954_ (_28407_, _28406_, _28402_);
  and _78955_ (_28408_, _28407_, _07793_);
  nor _78956_ (_28409_, _12003_, _10802_);
  nor _78957_ (_28410_, _28409_, _28321_);
  nor _78958_ (_28411_, _28410_, _07793_);
  or _78959_ (_28412_, _28411_, _28408_);
  and _78960_ (_28413_, _28412_, _04246_);
  nor _78961_ (_28414_, _28340_, _04246_);
  or _78962_ (_28416_, _28414_, _28413_);
  and _78963_ (_28417_, _28416_, _03823_);
  and _78964_ (_28418_, _28321_, _03453_);
  nor _78965_ (_28419_, _28418_, _03447_);
  not _78966_ (_28420_, _28419_);
  nor _78967_ (_28421_, _28420_, _28417_);
  and _78968_ (_28422_, _28340_, _03447_);
  or _78969_ (_28423_, _28422_, _28421_);
  nand _78970_ (_28424_, _28423_, _43000_);
  or _78971_ (_28425_, _43000_, \oc8051_golden_model_1.TCON [0]);
  and _78972_ (_28426_, _28425_, _41806_);
  and _78973_ (_43613_, _28426_, _28424_);
  or _78974_ (_28427_, _05258_, \oc8051_golden_model_1.TCON [1]);
  and _78975_ (_28428_, _12213_, _05258_);
  not _78976_ (_28429_, _28428_);
  and _78977_ (_28430_, _28429_, _28427_);
  or _78978_ (_28431_, _28430_, _04081_);
  nand _78979_ (_28432_, _05258_, _03274_);
  and _78980_ (_28433_, _28432_, _28427_);
  and _78981_ (_28434_, _28433_, _04409_);
  not _78982_ (_28437_, \oc8051_golden_model_1.TCON [1]);
  nor _78983_ (_28438_, _04409_, _28437_);
  or _78984_ (_28439_, _28438_, _03610_);
  or _78985_ (_28440_, _28439_, _28434_);
  and _78986_ (_28441_, _28440_, _04055_);
  and _78987_ (_28442_, _28441_, _28431_);
  and _78988_ (_28443_, _12224_, _05927_);
  nor _78989_ (_28444_, _05927_, _28437_);
  or _78990_ (_28445_, _28444_, _03723_);
  or _78991_ (_28446_, _28445_, _28443_);
  and _78992_ (_28448_, _28446_, _14265_);
  or _78993_ (_28449_, _28448_, _28442_);
  nor _78994_ (_28450_, _05258_, _28437_);
  and _78995_ (_28451_, _05258_, _06764_);
  or _78996_ (_28452_, _28451_, _28450_);
  or _78997_ (_28453_, _28452_, _03996_);
  and _78998_ (_28454_, _28453_, _28449_);
  or _78999_ (_28455_, _28454_, _03729_);
  or _79000_ (_28456_, _28433_, _03737_);
  and _79001_ (_28457_, _28456_, _03736_);
  and _79002_ (_28459_, _28457_, _28455_);
  and _79003_ (_28460_, _12211_, _05927_);
  or _79004_ (_28461_, _28460_, _28444_);
  and _79005_ (_28462_, _28461_, _03714_);
  or _79006_ (_28463_, _28462_, _03719_);
  or _79007_ (_28464_, _28463_, _28459_);
  and _79008_ (_28465_, _28443_, _12239_);
  or _79009_ (_28466_, _28444_, _06840_);
  or _79010_ (_28467_, _28466_, _28465_);
  and _79011_ (_28468_, _28467_, _28464_);
  and _79012_ (_28470_, _28468_, _03710_);
  nor _79013_ (_28471_, _12256_, _10839_);
  or _79014_ (_28472_, _28444_, _28471_);
  and _79015_ (_28473_, _28472_, _03505_);
  or _79016_ (_28474_, _28473_, _07390_);
  or _79017_ (_28475_, _28474_, _28470_);
  or _79018_ (_28476_, _28452_, _06838_);
  and _79019_ (_28477_, _28476_, _28475_);
  or _79020_ (_28478_, _28477_, _04481_);
  and _79021_ (_28479_, _06501_, _05258_);
  or _79022_ (_28481_, _28450_, _07400_);
  or _79023_ (_28482_, _28481_, _28479_);
  and _79024_ (_28483_, _28482_, _03589_);
  and _79025_ (_28484_, _28483_, _28478_);
  nor _79026_ (_28485_, _12313_, _10802_);
  or _79027_ (_28486_, _28485_, _28450_);
  and _79028_ (_28487_, _28486_, _03222_);
  or _79029_ (_28488_, _28487_, _28484_);
  and _79030_ (_28489_, _28488_, _03602_);
  or _79031_ (_28490_, _12327_, _10802_);
  and _79032_ (_28492_, _28490_, _03600_);
  nand _79033_ (_28493_, _05258_, _04303_);
  and _79034_ (_28494_, _28493_, _03601_);
  or _79035_ (_28495_, _28494_, _28492_);
  and _79036_ (_28496_, _28495_, _28427_);
  or _79037_ (_28497_, _28496_, _28489_);
  and _79038_ (_28498_, _28497_, _07778_);
  or _79039_ (_28499_, _12333_, _10802_);
  and _79040_ (_28500_, _28427_, _03780_);
  and _79041_ (_28501_, _28500_, _28499_);
  or _79042_ (_28503_, _28501_, _28498_);
  and _79043_ (_28504_, _28503_, _07777_);
  or _79044_ (_28505_, _12207_, _10802_);
  and _79045_ (_28506_, _28427_, _03622_);
  and _79046_ (_28507_, _28506_, _28505_);
  or _79047_ (_28508_, _28507_, _28504_);
  and _79048_ (_28509_, _28508_, _06828_);
  or _79049_ (_28510_, _28450_, _05618_);
  and _79050_ (_28511_, _28433_, _03790_);
  and _79051_ (_28512_, _28511_, _28510_);
  or _79052_ (_28514_, _28512_, _28509_);
  and _79053_ (_28515_, _28514_, _03786_);
  or _79054_ (_28516_, _28493_, _05618_);
  and _79055_ (_28517_, _28427_, _03624_);
  and _79056_ (_28518_, _28517_, _28516_);
  or _79057_ (_28519_, _28432_, _05618_);
  and _79058_ (_28520_, _28427_, _03785_);
  and _79059_ (_28521_, _28520_, _28519_);
  or _79060_ (_28522_, _28521_, _03815_);
  or _79061_ (_28523_, _28522_, _28518_);
  or _79062_ (_28525_, _28523_, _28515_);
  or _79063_ (_28526_, _28430_, _04246_);
  and _79064_ (_28527_, _28526_, _03823_);
  and _79065_ (_28528_, _28527_, _28525_);
  and _79066_ (_28529_, _28461_, _03453_);
  or _79067_ (_28530_, _28529_, _03447_);
  or _79068_ (_28531_, _28530_, _28528_);
  or _79069_ (_28532_, _28450_, _03514_);
  or _79070_ (_28533_, _28532_, _28428_);
  and _79071_ (_28534_, _28533_, _28531_);
  and _79072_ (_28536_, _28534_, _43000_);
  nor _79073_ (_28537_, \oc8051_golden_model_1.TCON [1], rst);
  nor _79074_ (_28538_, _28537_, _00000_);
  or _79075_ (_43614_, _28538_, _28536_);
  not _79076_ (_28539_, \oc8051_golden_model_1.TCON [2]);
  nor _79077_ (_28540_, _05258_, _28539_);
  and _79078_ (_28541_, _05258_, _06332_);
  nor _79079_ (_28542_, _28541_, _28540_);
  and _79080_ (_28543_, _28542_, _03601_);
  nor _79081_ (_28544_, _10802_, _04875_);
  nor _79082_ (_28546_, _28544_, _28540_);
  and _79083_ (_28547_, _28546_, _07390_);
  and _79084_ (_28548_, _05258_, \oc8051_golden_model_1.ACC [2]);
  nor _79085_ (_28549_, _28548_, _28540_);
  nor _79086_ (_28550_, _28549_, _09029_);
  nor _79087_ (_28551_, _04409_, _28539_);
  or _79088_ (_28552_, _28551_, _28550_);
  and _79089_ (_28553_, _28552_, _04081_);
  nor _79090_ (_28554_, _12416_, _10802_);
  nor _79091_ (_28555_, _28554_, _28540_);
  nor _79092_ (_28557_, _28555_, _04081_);
  or _79093_ (_28558_, _28557_, _28553_);
  and _79094_ (_28559_, _28558_, _04055_);
  nor _79095_ (_28560_, _05927_, _28539_);
  and _79096_ (_28561_, _12411_, _05927_);
  nor _79097_ (_28562_, _28561_, _28560_);
  nor _79098_ (_28563_, _28562_, _04055_);
  or _79099_ (_28564_, _28563_, _28559_);
  and _79100_ (_28565_, _28564_, _03996_);
  nor _79101_ (_28566_, _28546_, _03996_);
  or _79102_ (_28568_, _28566_, _28565_);
  and _79103_ (_28569_, _28568_, _03737_);
  nor _79104_ (_28570_, _28549_, _03737_);
  or _79105_ (_28571_, _28570_, _28569_);
  and _79106_ (_28572_, _28571_, _03736_);
  and _79107_ (_28573_, _12409_, _05927_);
  nor _79108_ (_28574_, _28573_, _28560_);
  nor _79109_ (_28575_, _28574_, _03736_);
  or _79110_ (_28576_, _28575_, _03719_);
  or _79111_ (_28577_, _28576_, _28572_);
  and _79112_ (_28579_, _28561_, _12443_);
  or _79113_ (_28580_, _28560_, _06840_);
  or _79114_ (_28581_, _28580_, _28579_);
  and _79115_ (_28582_, _28581_, _03710_);
  and _79116_ (_28583_, _28582_, _28577_);
  nor _79117_ (_28584_, _12461_, _10839_);
  nor _79118_ (_28585_, _28584_, _28560_);
  nor _79119_ (_28586_, _28585_, _03710_);
  nor _79120_ (_28587_, _28586_, _07390_);
  not _79121_ (_28588_, _28587_);
  nor _79122_ (_28590_, _28588_, _28583_);
  nor _79123_ (_28591_, _28590_, _28547_);
  nor _79124_ (_28592_, _28591_, _04481_);
  and _79125_ (_28593_, _06637_, _05258_);
  nor _79126_ (_28594_, _28540_, _07400_);
  not _79127_ (_28595_, _28594_);
  nor _79128_ (_28596_, _28595_, _28593_);
  or _79129_ (_28597_, _28596_, _03222_);
  nor _79130_ (_28598_, _28597_, _28592_);
  nor _79131_ (_28599_, _12519_, _10802_);
  nor _79132_ (_28601_, _28540_, _28599_);
  nor _79133_ (_28602_, _28601_, _03589_);
  or _79134_ (_28603_, _28602_, _03601_);
  nor _79135_ (_28604_, _28603_, _28598_);
  nor _79136_ (_28605_, _28604_, _28543_);
  or _79137_ (_28606_, _28605_, _03600_);
  and _79138_ (_28607_, _12533_, _05258_);
  or _79139_ (_28608_, _28607_, _28540_);
  or _79140_ (_28609_, _28608_, _07766_);
  and _79141_ (_28610_, _28609_, _07778_);
  and _79142_ (_28612_, _28610_, _28606_);
  and _79143_ (_28613_, _12539_, _05258_);
  nor _79144_ (_28614_, _28613_, _28540_);
  nor _79145_ (_28615_, _28614_, _07778_);
  nor _79146_ (_28616_, _28615_, _28612_);
  nor _79147_ (_28617_, _28616_, _03622_);
  nor _79148_ (_28618_, _28540_, _05718_);
  not _79149_ (_28619_, _28618_);
  nor _79150_ (_28620_, _28542_, _07777_);
  and _79151_ (_28621_, _28620_, _28619_);
  nor _79152_ (_28623_, _28621_, _28617_);
  nor _79153_ (_28624_, _28623_, _03790_);
  nor _79154_ (_28625_, _28549_, _06828_);
  and _79155_ (_28626_, _28625_, _28619_);
  or _79156_ (_28627_, _28626_, _28624_);
  and _79157_ (_28628_, _28627_, _07795_);
  nor _79158_ (_28629_, _12532_, _10802_);
  nor _79159_ (_28630_, _28629_, _28540_);
  nor _79160_ (_28631_, _28630_, _07795_);
  or _79161_ (_28632_, _28631_, _28628_);
  and _79162_ (_28634_, _28632_, _07793_);
  nor _79163_ (_28635_, _12538_, _10802_);
  nor _79164_ (_28636_, _28635_, _28540_);
  nor _79165_ (_28637_, _28636_, _07793_);
  or _79166_ (_28638_, _28637_, _28634_);
  and _79167_ (_28639_, _28638_, _04246_);
  nor _79168_ (_28640_, _28555_, _04246_);
  or _79169_ (_28641_, _28640_, _28639_);
  and _79170_ (_28642_, _28641_, _03823_);
  nor _79171_ (_28643_, _28574_, _03823_);
  or _79172_ (_28645_, _28643_, _28642_);
  and _79173_ (_28646_, _28645_, _03514_);
  and _79174_ (_28647_, _12592_, _05258_);
  nor _79175_ (_28648_, _28647_, _28540_);
  nor _79176_ (_28649_, _28648_, _03514_);
  or _79177_ (_28650_, _28649_, _28646_);
  or _79178_ (_28651_, _28650_, _43004_);
  or _79179_ (_28652_, _43000_, \oc8051_golden_model_1.TCON [2]);
  and _79180_ (_28653_, _28652_, _41806_);
  and _79181_ (_43615_, _28653_, _28651_);
  not _79182_ (_28655_, \oc8051_golden_model_1.TCON [3]);
  nor _79183_ (_28656_, _05258_, _28655_);
  and _79184_ (_28657_, _05258_, _06276_);
  nor _79185_ (_28658_, _28657_, _28656_);
  and _79186_ (_28659_, _28658_, _03601_);
  nor _79187_ (_28660_, _10802_, _05005_);
  nor _79188_ (_28661_, _28660_, _28656_);
  and _79189_ (_28662_, _28661_, _07390_);
  and _79190_ (_28663_, _05258_, \oc8051_golden_model_1.ACC [3]);
  nor _79191_ (_28664_, _28663_, _28656_);
  nor _79192_ (_28666_, _28664_, _09029_);
  nor _79193_ (_28667_, _04409_, _28655_);
  or _79194_ (_28668_, _28667_, _28666_);
  and _79195_ (_28669_, _28668_, _04081_);
  nor _79196_ (_28670_, _12627_, _10802_);
  nor _79197_ (_28671_, _28670_, _28656_);
  nor _79198_ (_28672_, _28671_, _04081_);
  or _79199_ (_28673_, _28672_, _28669_);
  and _79200_ (_28674_, _28673_, _04055_);
  nor _79201_ (_28675_, _05927_, _28655_);
  and _79202_ (_28677_, _12631_, _05927_);
  nor _79203_ (_28678_, _28677_, _28675_);
  nor _79204_ (_28679_, _28678_, _04055_);
  or _79205_ (_28680_, _28679_, _03723_);
  or _79206_ (_28681_, _28680_, _28674_);
  nand _79207_ (_28682_, _28661_, _03723_);
  and _79208_ (_28683_, _28682_, _28681_);
  and _79209_ (_28684_, _28683_, _03737_);
  nor _79210_ (_28685_, _28664_, _03737_);
  or _79211_ (_28686_, _28685_, _28684_);
  and _79212_ (_28688_, _28686_, _03736_);
  and _79213_ (_28689_, _12641_, _05927_);
  nor _79214_ (_28690_, _28689_, _28675_);
  nor _79215_ (_28691_, _28690_, _03736_);
  or _79216_ (_28692_, _28691_, _28688_);
  and _79217_ (_28693_, _28692_, _06840_);
  nor _79218_ (_28694_, _28675_, _12648_);
  nor _79219_ (_28695_, _28694_, _28678_);
  and _79220_ (_28696_, _28695_, _03719_);
  or _79221_ (_28697_, _28696_, _28693_);
  and _79222_ (_28699_, _28697_, _03710_);
  nor _79223_ (_28700_, _12612_, _10839_);
  nor _79224_ (_28701_, _28700_, _28675_);
  nor _79225_ (_28702_, _28701_, _03710_);
  nor _79226_ (_28703_, _28702_, _07390_);
  not _79227_ (_28704_, _28703_);
  nor _79228_ (_28705_, _28704_, _28699_);
  nor _79229_ (_28706_, _28705_, _28662_);
  nor _79230_ (_28707_, _28706_, _04481_);
  and _79231_ (_28708_, _06592_, _05258_);
  nor _79232_ (_28710_, _28656_, _07400_);
  not _79233_ (_28711_, _28710_);
  nor _79234_ (_28712_, _28711_, _28708_);
  or _79235_ (_28713_, _28712_, _03222_);
  nor _79236_ (_28714_, _28713_, _28707_);
  nor _79237_ (_28715_, _12718_, _10802_);
  nor _79238_ (_28716_, _28656_, _28715_);
  nor _79239_ (_28717_, _28716_, _03589_);
  or _79240_ (_28718_, _28717_, _03601_);
  nor _79241_ (_28719_, _28718_, _28714_);
  nor _79242_ (_28721_, _28719_, _28659_);
  or _79243_ (_28722_, _28721_, _03600_);
  and _79244_ (_28723_, _12733_, _05258_);
  or _79245_ (_28724_, _28723_, _28656_);
  or _79246_ (_28725_, _28724_, _07766_);
  and _79247_ (_28726_, _28725_, _07778_);
  and _79248_ (_28727_, _28726_, _28722_);
  and _79249_ (_28728_, _12739_, _05258_);
  nor _79250_ (_28729_, _28728_, _28656_);
  nor _79251_ (_28730_, _28729_, _07778_);
  nor _79252_ (_28732_, _28730_, _28727_);
  nor _79253_ (_28733_, _28732_, _03622_);
  nor _79254_ (_28734_, _28656_, _05567_);
  not _79255_ (_28735_, _28734_);
  nor _79256_ (_28736_, _28658_, _07777_);
  and _79257_ (_28737_, _28736_, _28735_);
  nor _79258_ (_28738_, _28737_, _28733_);
  nor _79259_ (_28739_, _28738_, _03790_);
  nor _79260_ (_28740_, _28664_, _06828_);
  and _79261_ (_28741_, _28740_, _28735_);
  or _79262_ (_28743_, _28741_, _28739_);
  and _79263_ (_28744_, _28743_, _07795_);
  nor _79264_ (_28745_, _12732_, _10802_);
  nor _79265_ (_28746_, _28745_, _28656_);
  nor _79266_ (_28747_, _28746_, _07795_);
  or _79267_ (_28748_, _28747_, _28744_);
  and _79268_ (_28749_, _28748_, _07793_);
  nor _79269_ (_28750_, _12738_, _10802_);
  nor _79270_ (_28751_, _28750_, _28656_);
  nor _79271_ (_28752_, _28751_, _07793_);
  or _79272_ (_28754_, _28752_, _28749_);
  and _79273_ (_28755_, _28754_, _04246_);
  nor _79274_ (_28756_, _28671_, _04246_);
  or _79275_ (_28757_, _28756_, _28755_);
  and _79276_ (_28758_, _28757_, _03823_);
  nor _79277_ (_28759_, _28690_, _03823_);
  nor _79278_ (_28760_, _28759_, _03447_);
  not _79279_ (_28761_, _28760_);
  nor _79280_ (_28762_, _28761_, _28758_);
  and _79281_ (_28763_, _12794_, _05258_);
  or _79282_ (_28765_, _28656_, _03514_);
  nor _79283_ (_28766_, _28765_, _28763_);
  nor _79284_ (_28767_, _28766_, _28762_);
  or _79285_ (_28768_, _28767_, _43004_);
  or _79286_ (_28769_, _43000_, \oc8051_golden_model_1.TCON [3]);
  and _79287_ (_28770_, _28769_, _41806_);
  and _79288_ (_43618_, _28770_, _28768_);
  not _79289_ (_28771_, \oc8051_golden_model_1.TCON [4]);
  nor _79290_ (_28772_, _05258_, _28771_);
  nor _79291_ (_28773_, _05777_, _10802_);
  nor _79292_ (_28775_, _28773_, _28772_);
  and _79293_ (_28776_, _28775_, _07390_);
  nor _79294_ (_28777_, _05927_, _28771_);
  and _79295_ (_28778_, _12827_, _05927_);
  nor _79296_ (_28779_, _28778_, _28777_);
  nor _79297_ (_28780_, _28779_, _03736_);
  and _79298_ (_28781_, _05258_, \oc8051_golden_model_1.ACC [4]);
  nor _79299_ (_28782_, _28781_, _28772_);
  nor _79300_ (_28783_, _28782_, _09029_);
  nor _79301_ (_28784_, _04409_, _28771_);
  or _79302_ (_28786_, _28784_, _28783_);
  and _79303_ (_28787_, _28786_, _04081_);
  nor _79304_ (_28788_, _12841_, _10802_);
  nor _79305_ (_28789_, _28788_, _28772_);
  nor _79306_ (_28790_, _28789_, _04081_);
  or _79307_ (_28791_, _28790_, _28787_);
  and _79308_ (_28792_, _28791_, _04055_);
  and _79309_ (_28793_, _12845_, _05927_);
  nor _79310_ (_28794_, _28793_, _28777_);
  nor _79311_ (_28795_, _28794_, _04055_);
  or _79312_ (_28797_, _28795_, _03723_);
  or _79313_ (_28798_, _28797_, _28792_);
  nand _79314_ (_28799_, _28775_, _03723_);
  and _79315_ (_28800_, _28799_, _28798_);
  and _79316_ (_28801_, _28800_, _03737_);
  nor _79317_ (_28802_, _28782_, _03737_);
  or _79318_ (_28803_, _28802_, _28801_);
  and _79319_ (_28804_, _28803_, _03736_);
  nor _79320_ (_28805_, _28804_, _28780_);
  nor _79321_ (_28806_, _28805_, _03719_);
  nor _79322_ (_28807_, _28777_, _12860_);
  or _79323_ (_28808_, _28794_, _06840_);
  nor _79324_ (_28809_, _28808_, _28807_);
  nor _79325_ (_28810_, _28809_, _28806_);
  nor _79326_ (_28811_, _28810_, _03505_);
  nor _79327_ (_28812_, _12825_, _10839_);
  nor _79328_ (_28813_, _28812_, _28777_);
  nor _79329_ (_28814_, _28813_, _03710_);
  nor _79330_ (_28815_, _28814_, _07390_);
  not _79331_ (_28816_, _28815_);
  nor _79332_ (_28818_, _28816_, _28811_);
  nor _79333_ (_28819_, _28818_, _28776_);
  nor _79334_ (_28820_, _28819_, _04481_);
  and _79335_ (_28821_, _06730_, _05258_);
  nor _79336_ (_28822_, _28772_, _07400_);
  not _79337_ (_28823_, _28822_);
  nor _79338_ (_28824_, _28823_, _28821_);
  nor _79339_ (_28825_, _28824_, _03222_);
  not _79340_ (_28826_, _28825_);
  nor _79341_ (_28827_, _28826_, _28820_);
  nor _79342_ (_28829_, _12933_, _10802_);
  nor _79343_ (_28830_, _28829_, _28772_);
  nor _79344_ (_28831_, _28830_, _03589_);
  or _79345_ (_28832_, _28831_, _08828_);
  or _79346_ (_28833_, _28832_, _28827_);
  and _79347_ (_28834_, _12821_, _05258_);
  or _79348_ (_28835_, _28772_, _07766_);
  or _79349_ (_28836_, _28835_, _28834_);
  and _79350_ (_28837_, _06298_, _05258_);
  nor _79351_ (_28838_, _28837_, _28772_);
  and _79352_ (_28840_, _28838_, _03601_);
  nor _79353_ (_28841_, _28840_, _03780_);
  and _79354_ (_28842_, _28841_, _28836_);
  and _79355_ (_28843_, _28842_, _28833_);
  and _79356_ (_28844_, _12817_, _05258_);
  nor _79357_ (_28845_, _28844_, _28772_);
  nor _79358_ (_28846_, _28845_, _07778_);
  nor _79359_ (_28847_, _28846_, _28843_);
  nor _79360_ (_28848_, _28847_, _03622_);
  nor _79361_ (_28849_, _28772_, _05825_);
  not _79362_ (_28851_, _28849_);
  nor _79363_ (_28852_, _28838_, _07777_);
  and _79364_ (_28853_, _28852_, _28851_);
  nor _79365_ (_28854_, _28853_, _28848_);
  nor _79366_ (_28855_, _28854_, _03790_);
  nor _79367_ (_28856_, _28782_, _06828_);
  and _79368_ (_28857_, _28856_, _28851_);
  or _79369_ (_28858_, _28857_, _28855_);
  and _79370_ (_28859_, _28858_, _07795_);
  nor _79371_ (_28860_, _12819_, _10802_);
  nor _79372_ (_28862_, _28860_, _28772_);
  nor _79373_ (_28863_, _28862_, _07795_);
  or _79374_ (_28864_, _28863_, _28859_);
  and _79375_ (_28865_, _28864_, _07793_);
  nor _79376_ (_28866_, _12816_, _10802_);
  nor _79377_ (_28867_, _28866_, _28772_);
  nor _79378_ (_28868_, _28867_, _07793_);
  or _79379_ (_28869_, _28868_, _28865_);
  and _79380_ (_28870_, _28869_, _04246_);
  nor _79381_ (_28871_, _28789_, _04246_);
  or _79382_ (_28873_, _28871_, _28870_);
  and _79383_ (_28874_, _28873_, _03823_);
  nor _79384_ (_28875_, _28779_, _03823_);
  nor _79385_ (_28876_, _28875_, _03447_);
  not _79386_ (_28877_, _28876_);
  nor _79387_ (_28878_, _28877_, _28874_);
  and _79388_ (_28879_, _13003_, _05258_);
  or _79389_ (_28880_, _28772_, _03514_);
  nor _79390_ (_28881_, _28880_, _28879_);
  nor _79391_ (_28882_, _28881_, _28878_);
  or _79392_ (_28884_, _28882_, _43004_);
  or _79393_ (_28885_, _43000_, \oc8051_golden_model_1.TCON [4]);
  and _79394_ (_28886_, _28885_, _41806_);
  and _79395_ (_43619_, _28886_, _28884_);
  not _79396_ (_28887_, \oc8051_golden_model_1.TCON [5]);
  nor _79397_ (_28888_, _05258_, _28887_);
  and _79398_ (_28889_, _06684_, _05258_);
  or _79399_ (_28890_, _28889_, _28888_);
  and _79400_ (_28891_, _28890_, _04481_);
  and _79401_ (_28892_, _05258_, \oc8051_golden_model_1.ACC [5]);
  nor _79402_ (_28894_, _28892_, _28888_);
  nor _79403_ (_28895_, _28894_, _09029_);
  nor _79404_ (_28896_, _04409_, _28887_);
  or _79405_ (_28897_, _28896_, _28895_);
  and _79406_ (_28898_, _28897_, _04081_);
  nor _79407_ (_28899_, _13014_, _10802_);
  nor _79408_ (_28900_, _28899_, _28888_);
  nor _79409_ (_28901_, _28900_, _04081_);
  or _79410_ (_28902_, _28901_, _28898_);
  and _79411_ (_28903_, _28902_, _04055_);
  nor _79412_ (_28905_, _05927_, _28887_);
  and _79413_ (_28906_, _13037_, _05927_);
  nor _79414_ (_28907_, _28906_, _28905_);
  nor _79415_ (_28908_, _28907_, _04055_);
  or _79416_ (_28909_, _28908_, _03723_);
  or _79417_ (_28910_, _28909_, _28903_);
  nor _79418_ (_28911_, _05469_, _10802_);
  nor _79419_ (_28912_, _28911_, _28888_);
  nand _79420_ (_28913_, _28912_, _03723_);
  and _79421_ (_28914_, _28913_, _28910_);
  and _79422_ (_28916_, _28914_, _03737_);
  nor _79423_ (_28917_, _28894_, _03737_);
  or _79424_ (_28918_, _28917_, _28916_);
  and _79425_ (_28919_, _28918_, _03736_);
  and _79426_ (_28920_, _13047_, _05927_);
  nor _79427_ (_28921_, _28920_, _28905_);
  nor _79428_ (_28922_, _28921_, _03736_);
  or _79429_ (_28923_, _28922_, _03719_);
  or _79430_ (_28924_, _28923_, _28919_);
  nor _79431_ (_28925_, _28905_, _13054_);
  nor _79432_ (_28927_, _28925_, _28907_);
  or _79433_ (_28928_, _28927_, _06840_);
  and _79434_ (_28929_, _28928_, _03710_);
  and _79435_ (_28930_, _28929_, _28924_);
  nor _79436_ (_28931_, _13020_, _10839_);
  nor _79437_ (_28932_, _28931_, _28905_);
  nor _79438_ (_28933_, _28932_, _03710_);
  nor _79439_ (_28934_, _28933_, _07390_);
  not _79440_ (_28935_, _28934_);
  nor _79441_ (_28936_, _28935_, _28930_);
  and _79442_ (_28938_, _28912_, _07390_);
  or _79443_ (_28939_, _28938_, _04481_);
  nor _79444_ (_28940_, _28939_, _28936_);
  or _79445_ (_28941_, _28940_, _28891_);
  and _79446_ (_28942_, _28941_, _03589_);
  nor _79447_ (_28943_, _13127_, _10802_);
  nor _79448_ (_28944_, _28943_, _28888_);
  nor _79449_ (_28945_, _28944_, _03589_);
  or _79450_ (_28946_, _28945_, _08828_);
  or _79451_ (_28947_, _28946_, _28942_);
  and _79452_ (_28949_, _13141_, _05258_);
  or _79453_ (_28950_, _28888_, _07766_);
  or _79454_ (_28951_, _28950_, _28949_);
  and _79455_ (_28952_, _06306_, _05258_);
  nor _79456_ (_28953_, _28952_, _28888_);
  and _79457_ (_28954_, _28953_, _03601_);
  nor _79458_ (_28955_, _28954_, _03780_);
  and _79459_ (_28956_, _28955_, _28951_);
  and _79460_ (_28957_, _28956_, _28947_);
  and _79461_ (_28958_, _13147_, _05258_);
  nor _79462_ (_28959_, _28958_, _28888_);
  nor _79463_ (_28960_, _28959_, _07778_);
  nor _79464_ (_28961_, _28960_, _28957_);
  nor _79465_ (_28962_, _28961_, _03622_);
  nor _79466_ (_28963_, _28888_, _05518_);
  not _79467_ (_28964_, _28963_);
  nor _79468_ (_28965_, _28953_, _07777_);
  and _79469_ (_28966_, _28965_, _28964_);
  nor _79470_ (_28967_, _28966_, _28962_);
  nor _79471_ (_28968_, _28967_, _03790_);
  nor _79472_ (_28971_, _28894_, _06828_);
  and _79473_ (_28972_, _28971_, _28964_);
  nor _79474_ (_28973_, _28972_, _03624_);
  not _79475_ (_28974_, _28973_);
  nor _79476_ (_28975_, _28974_, _28968_);
  nor _79477_ (_28976_, _13140_, _10802_);
  or _79478_ (_28977_, _28888_, _07795_);
  nor _79479_ (_28978_, _28977_, _28976_);
  or _79480_ (_28979_, _28978_, _03785_);
  nor _79481_ (_28980_, _28979_, _28975_);
  nor _79482_ (_28982_, _13146_, _10802_);
  nor _79483_ (_28983_, _28982_, _28888_);
  nor _79484_ (_28984_, _28983_, _07793_);
  or _79485_ (_28985_, _28984_, _28980_);
  and _79486_ (_28986_, _28985_, _04246_);
  nor _79487_ (_28987_, _28900_, _04246_);
  or _79488_ (_28988_, _28987_, _28986_);
  and _79489_ (_28989_, _28988_, _03823_);
  nor _79490_ (_28990_, _28921_, _03823_);
  or _79491_ (_28991_, _28990_, _28989_);
  and _79492_ (_28993_, _28991_, _03514_);
  and _79493_ (_28994_, _13199_, _05258_);
  nor _79494_ (_28995_, _28994_, _28888_);
  nor _79495_ (_28996_, _28995_, _03514_);
  or _79496_ (_28997_, _28996_, _28993_);
  or _79497_ (_28998_, _28997_, _43004_);
  or _79498_ (_28999_, _43000_, \oc8051_golden_model_1.TCON [5]);
  and _79499_ (_29000_, _28999_, _41806_);
  and _79500_ (_43620_, _29000_, _28998_);
  not _79501_ (_29001_, \oc8051_golden_model_1.TCON [6]);
  nor _79502_ (_29003_, _05258_, _29001_);
  and _79503_ (_29004_, _06455_, _05258_);
  or _79504_ (_29005_, _29004_, _29003_);
  and _79505_ (_29006_, _29005_, _04481_);
  and _79506_ (_29007_, _05258_, \oc8051_golden_model_1.ACC [6]);
  nor _79507_ (_29008_, _29007_, _29003_);
  nor _79508_ (_29009_, _29008_, _09029_);
  nor _79509_ (_29010_, _04409_, _29001_);
  or _79510_ (_29011_, _29010_, _29009_);
  and _79511_ (_29012_, _29011_, _04081_);
  nor _79512_ (_29014_, _13242_, _10802_);
  nor _79513_ (_29015_, _29014_, _29003_);
  nor _79514_ (_29016_, _29015_, _04081_);
  or _79515_ (_29017_, _29016_, _29012_);
  and _79516_ (_29018_, _29017_, _04055_);
  nor _79517_ (_29019_, _05927_, _29001_);
  and _79518_ (_29020_, _13229_, _05927_);
  nor _79519_ (_29021_, _29020_, _29019_);
  nor _79520_ (_29022_, _29021_, _04055_);
  or _79521_ (_29023_, _29022_, _03723_);
  or _79522_ (_29025_, _29023_, _29018_);
  nor _79523_ (_29026_, _05363_, _10802_);
  nor _79524_ (_29027_, _29026_, _29003_);
  nand _79525_ (_29028_, _29027_, _03723_);
  and _79526_ (_29029_, _29028_, _29025_);
  and _79527_ (_29030_, _29029_, _03737_);
  nor _79528_ (_29031_, _29008_, _03737_);
  or _79529_ (_29032_, _29031_, _29030_);
  and _79530_ (_29033_, _29032_, _03736_);
  and _79531_ (_29034_, _13253_, _05927_);
  nor _79532_ (_29036_, _29034_, _29019_);
  nor _79533_ (_29037_, _29036_, _03736_);
  or _79534_ (_29038_, _29037_, _29033_);
  and _79535_ (_29039_, _29038_, _06840_);
  nor _79536_ (_29040_, _29019_, _13260_);
  nor _79537_ (_29041_, _29040_, _29021_);
  and _79538_ (_29042_, _29041_, _03719_);
  or _79539_ (_29043_, _29042_, _29039_);
  and _79540_ (_29044_, _29043_, _03710_);
  nor _79541_ (_29045_, _13226_, _10839_);
  nor _79542_ (_29047_, _29045_, _29019_);
  nor _79543_ (_29048_, _29047_, _03710_);
  nor _79544_ (_29049_, _29048_, _07390_);
  not _79545_ (_29050_, _29049_);
  nor _79546_ (_29051_, _29050_, _29044_);
  and _79547_ (_29052_, _29027_, _07390_);
  or _79548_ (_29053_, _29052_, _04481_);
  nor _79549_ (_29054_, _29053_, _29051_);
  or _79550_ (_29055_, _29054_, _29006_);
  and _79551_ (_29056_, _29055_, _03589_);
  nor _79552_ (_29058_, _13332_, _10802_);
  nor _79553_ (_29059_, _29058_, _29003_);
  nor _79554_ (_29060_, _29059_, _03589_);
  or _79555_ (_29061_, _29060_, _08828_);
  or _79556_ (_29062_, _29061_, _29056_);
  and _79557_ (_29063_, _13347_, _05258_);
  or _79558_ (_29064_, _29003_, _07766_);
  or _79559_ (_29065_, _29064_, _29063_);
  and _79560_ (_29066_, _13339_, _05258_);
  nor _79561_ (_29067_, _29066_, _29003_);
  and _79562_ (_29069_, _29067_, _03601_);
  nor _79563_ (_29070_, _29069_, _03780_);
  and _79564_ (_29071_, _29070_, _29065_);
  and _79565_ (_29072_, _29071_, _29062_);
  and _79566_ (_29073_, _13353_, _05258_);
  nor _79567_ (_29074_, _29073_, _29003_);
  nor _79568_ (_29075_, _29074_, _07778_);
  nor _79569_ (_29076_, _29075_, _29072_);
  nor _79570_ (_29077_, _29076_, _03622_);
  nor _79571_ (_29078_, _29003_, _05412_);
  not _79572_ (_29080_, _29078_);
  nor _79573_ (_29081_, _29067_, _07777_);
  and _79574_ (_29082_, _29081_, _29080_);
  nor _79575_ (_29083_, _29082_, _29077_);
  nor _79576_ (_29084_, _29083_, _03790_);
  nor _79577_ (_29085_, _29008_, _06828_);
  and _79578_ (_29086_, _29085_, _29080_);
  nor _79579_ (_29087_, _29086_, _03624_);
  not _79580_ (_29088_, _29087_);
  nor _79581_ (_29089_, _29088_, _29084_);
  nor _79582_ (_29091_, _13346_, _10802_);
  or _79583_ (_29092_, _29003_, _07795_);
  nor _79584_ (_29093_, _29092_, _29091_);
  or _79585_ (_29094_, _29093_, _03785_);
  nor _79586_ (_29095_, _29094_, _29089_);
  nor _79587_ (_29096_, _13352_, _10802_);
  nor _79588_ (_29097_, _29096_, _29003_);
  nor _79589_ (_29098_, _29097_, _07793_);
  or _79590_ (_29099_, _29098_, _29095_);
  and _79591_ (_29100_, _29099_, _04246_);
  nor _79592_ (_29102_, _29015_, _04246_);
  or _79593_ (_29103_, _29102_, _29100_);
  and _79594_ (_29104_, _29103_, _03823_);
  nor _79595_ (_29105_, _29036_, _03823_);
  or _79596_ (_29106_, _29105_, _29104_);
  and _79597_ (_29107_, _29106_, _03514_);
  and _79598_ (_29108_, _13402_, _05258_);
  nor _79599_ (_29109_, _29108_, _29003_);
  nor _79600_ (_29110_, _29109_, _03514_);
  or _79601_ (_29111_, _29110_, _29107_);
  or _79602_ (_29113_, _29111_, _43004_);
  or _79603_ (_29114_, _43000_, \oc8051_golden_model_1.TCON [6]);
  and _79604_ (_29115_, _29114_, _41806_);
  and _79605_ (_43621_, _29115_, _29113_);
  not _79606_ (_29116_, \oc8051_golden_model_1.TH0 [0]);
  nor _79607_ (_29117_, _05263_, _29116_);
  nor _79608_ (_29118_, _05666_, _10909_);
  nor _79609_ (_29119_, _29118_, _29117_);
  and _79610_ (_29120_, _29119_, _17166_);
  and _79611_ (_29121_, _05263_, \oc8051_golden_model_1.ACC [0]);
  nor _79612_ (_29123_, _29121_, _29117_);
  nor _79613_ (_29124_, _29123_, _03737_);
  nor _79614_ (_29125_, _29124_, _07390_);
  nor _79615_ (_29126_, _29119_, _04081_);
  nor _79616_ (_29127_, _04409_, _29116_);
  nor _79617_ (_29128_, _29123_, _09029_);
  nor _79618_ (_29129_, _29128_, _29127_);
  nor _79619_ (_29130_, _29129_, _03610_);
  or _79620_ (_29131_, _29130_, _03723_);
  nor _79621_ (_29132_, _29131_, _29126_);
  or _79622_ (_29134_, _29132_, _03729_);
  and _79623_ (_29135_, _29134_, _29125_);
  and _79624_ (_29136_, _05263_, _04620_);
  or _79625_ (_29137_, _29117_, _25480_);
  nor _79626_ (_29138_, _29137_, _29136_);
  nor _79627_ (_29139_, _29138_, _29135_);
  nor _79628_ (_29140_, _29139_, _04481_);
  and _79629_ (_29141_, _06546_, _05263_);
  nor _79630_ (_29142_, _29117_, _07400_);
  not _79631_ (_29143_, _29142_);
  nor _79632_ (_29145_, _29143_, _29141_);
  nor _79633_ (_29146_, _29145_, _29140_);
  nor _79634_ (_29147_, _29146_, _03222_);
  nor _79635_ (_29148_, _12109_, _10909_);
  or _79636_ (_29149_, _29117_, _03589_);
  nor _79637_ (_29150_, _29149_, _29148_);
  or _79638_ (_29151_, _29150_, _03601_);
  nor _79639_ (_29152_, _29151_, _29147_);
  and _79640_ (_29153_, _05263_, _06274_);
  nor _79641_ (_29154_, _29153_, _29117_);
  nand _79642_ (_29156_, _29154_, _07766_);
  and _79643_ (_29157_, _29156_, _08828_);
  nor _79644_ (_29158_, _29157_, _29152_);
  and _79645_ (_29159_, _12124_, _05263_);
  nor _79646_ (_29160_, _29159_, _29117_);
  and _79647_ (_29161_, _29160_, _03600_);
  nor _79648_ (_29162_, _29161_, _29158_);
  nor _79649_ (_29163_, _29162_, _03780_);
  and _79650_ (_29164_, _12128_, _05263_);
  or _79651_ (_29165_, _29117_, _07778_);
  nor _79652_ (_29167_, _29165_, _29164_);
  or _79653_ (_29168_, _29167_, _03622_);
  nor _79654_ (_29169_, _29168_, _29163_);
  or _79655_ (_29170_, _29154_, _07777_);
  nor _79656_ (_29171_, _29170_, _29118_);
  nor _79657_ (_29172_, _29171_, _29169_);
  nor _79658_ (_29173_, _29172_, _03790_);
  and _79659_ (_29174_, _12005_, _05263_);
  or _79660_ (_29175_, _29174_, _29117_);
  and _79661_ (_29176_, _29175_, _03790_);
  or _79662_ (_29178_, _29176_, _29173_);
  and _79663_ (_29179_, _29178_, _07795_);
  nor _79664_ (_29180_, _12122_, _10909_);
  nor _79665_ (_29181_, _29180_, _29117_);
  nor _79666_ (_29182_, _29181_, _07795_);
  or _79667_ (_29183_, _29182_, _29179_);
  and _79668_ (_29184_, _29183_, _07793_);
  nor _79669_ (_29185_, _12003_, _10909_);
  nor _79670_ (_29186_, _29185_, _29117_);
  nor _79671_ (_29187_, _29186_, _07793_);
  nor _79672_ (_29189_, _29187_, _17166_);
  not _79673_ (_29190_, _29189_);
  nor _79674_ (_29191_, _29190_, _29184_);
  nor _79675_ (_29192_, _29191_, _29120_);
  or _79676_ (_29193_, _29192_, _43004_);
  or _79677_ (_29194_, _43000_, \oc8051_golden_model_1.TH0 [0]);
  and _79678_ (_29195_, _29194_, _41806_);
  and _79679_ (_43624_, _29195_, _29193_);
  and _79680_ (_29196_, _06501_, _05263_);
  not _79681_ (_29197_, \oc8051_golden_model_1.TH0 [1]);
  nor _79682_ (_29199_, _05263_, _29197_);
  nor _79683_ (_29200_, _29199_, _07400_);
  not _79684_ (_29201_, _29200_);
  nor _79685_ (_29202_, _29201_, _29196_);
  not _79686_ (_29203_, _29202_);
  nor _79687_ (_29204_, _05263_, \oc8051_golden_model_1.TH0 [1]);
  and _79688_ (_29205_, _05263_, _03274_);
  nor _79689_ (_29206_, _29205_, _29204_);
  and _79690_ (_29207_, _29206_, _03729_);
  and _79691_ (_29208_, _29206_, _04409_);
  nor _79692_ (_29210_, _04409_, _29197_);
  or _79693_ (_29211_, _29210_, _29208_);
  and _79694_ (_29212_, _29211_, _04081_);
  and _79695_ (_29213_, _12213_, _05263_);
  nor _79696_ (_29214_, _29213_, _29204_);
  and _79697_ (_29215_, _29214_, _03610_);
  or _79698_ (_29216_, _29215_, _29212_);
  and _79699_ (_29217_, _29216_, _03996_);
  and _79700_ (_29218_, _05263_, _06764_);
  nor _79701_ (_29219_, _29218_, _29199_);
  nor _79702_ (_29221_, _29219_, _03996_);
  nor _79703_ (_29222_, _29221_, _29217_);
  nor _79704_ (_29223_, _29222_, _03729_);
  or _79705_ (_29224_, _29223_, _07390_);
  nor _79706_ (_29225_, _29224_, _29207_);
  and _79707_ (_29226_, _29219_, _07390_);
  nor _79708_ (_29227_, _29226_, _29225_);
  nor _79709_ (_29228_, _29227_, _04481_);
  nor _79710_ (_29229_, _29228_, _03222_);
  and _79711_ (_29230_, _29229_, _29203_);
  not _79712_ (_29232_, _29204_);
  and _79713_ (_29233_, _12313_, _05263_);
  nor _79714_ (_29234_, _29233_, _03589_);
  and _79715_ (_29235_, _29234_, _29232_);
  nor _79716_ (_29236_, _29235_, _29230_);
  nor _79717_ (_29237_, _29236_, _08828_);
  nor _79718_ (_29238_, _12327_, _10909_);
  nor _79719_ (_29239_, _29238_, _07766_);
  and _79720_ (_29240_, _05263_, _04303_);
  nor _79721_ (_29241_, _29240_, _05886_);
  nor _79722_ (_29243_, _29241_, _29239_);
  nor _79723_ (_29244_, _29243_, _29204_);
  nor _79724_ (_29245_, _29244_, _29237_);
  nor _79725_ (_29246_, _29245_, _03780_);
  nor _79726_ (_29247_, _12333_, _10909_);
  nor _79727_ (_29248_, _29247_, _07778_);
  and _79728_ (_29249_, _29248_, _29232_);
  nor _79729_ (_29250_, _29249_, _29246_);
  nor _79730_ (_29251_, _29250_, _03622_);
  nor _79731_ (_29252_, _12207_, _10909_);
  nor _79732_ (_29254_, _29252_, _07777_);
  and _79733_ (_29255_, _29254_, _29232_);
  nor _79734_ (_29256_, _29255_, _29251_);
  nor _79735_ (_29257_, _29256_, _03790_);
  nor _79736_ (_29258_, _29199_, _05618_);
  nor _79737_ (_29259_, _29258_, _06828_);
  and _79738_ (_29260_, _29259_, _29206_);
  nor _79739_ (_29261_, _29260_, _29257_);
  or _79740_ (_29262_, _29261_, _18499_);
  and _79741_ (_29263_, _29240_, _05617_);
  nor _79742_ (_29265_, _29263_, _07795_);
  and _79743_ (_29266_, _29265_, _29232_);
  nand _79744_ (_29267_, _29205_, _05617_);
  nor _79745_ (_29268_, _29204_, _07793_);
  and _79746_ (_29269_, _29268_, _29267_);
  or _79747_ (_29270_, _29269_, _03815_);
  nor _79748_ (_29271_, _29270_, _29266_);
  and _79749_ (_29272_, _29271_, _29262_);
  nor _79750_ (_29273_, _29214_, _04246_);
  nor _79751_ (_29274_, _29273_, _29272_);
  and _79752_ (_29276_, _29274_, _03514_);
  nor _79753_ (_29277_, _29213_, _29199_);
  nor _79754_ (_29278_, _29277_, _03514_);
  or _79755_ (_29279_, _29278_, _29276_);
  or _79756_ (_29280_, _29279_, _43004_);
  or _79757_ (_29281_, _43000_, \oc8051_golden_model_1.TH0 [1]);
  and _79758_ (_29282_, _29281_, _41806_);
  and _79759_ (_43625_, _29282_, _29280_);
  not _79760_ (_29283_, \oc8051_golden_model_1.TH0 [2]);
  nor _79761_ (_29284_, _05263_, _29283_);
  nor _79762_ (_29286_, _12538_, _10909_);
  nor _79763_ (_29287_, _29286_, _29284_);
  nor _79764_ (_29288_, _29287_, _07793_);
  nor _79765_ (_29289_, _10909_, _04875_);
  nor _79766_ (_29290_, _29289_, _29284_);
  and _79767_ (_29291_, _29290_, _07390_);
  nor _79768_ (_29292_, _12416_, _10909_);
  nor _79769_ (_29293_, _29292_, _29284_);
  nor _79770_ (_29294_, _29293_, _04081_);
  nor _79771_ (_29295_, _04409_, _29283_);
  and _79772_ (_29297_, _05263_, \oc8051_golden_model_1.ACC [2]);
  nor _79773_ (_29298_, _29297_, _29284_);
  nor _79774_ (_29299_, _29298_, _09029_);
  nor _79775_ (_29300_, _29299_, _29295_);
  nor _79776_ (_29301_, _29300_, _03610_);
  or _79777_ (_29302_, _29301_, _29294_);
  and _79778_ (_29303_, _29302_, _03996_);
  nor _79779_ (_29304_, _29290_, _03996_);
  or _79780_ (_29305_, _29304_, _29303_);
  and _79781_ (_29306_, _29305_, _03737_);
  nor _79782_ (_29308_, _29298_, _03737_);
  nor _79783_ (_29309_, _29308_, _07390_);
  not _79784_ (_29310_, _29309_);
  nor _79785_ (_29311_, _29310_, _29306_);
  nor _79786_ (_29312_, _29311_, _29291_);
  nor _79787_ (_29313_, _29312_, _04481_);
  and _79788_ (_29314_, _06637_, _05263_);
  nor _79789_ (_29315_, _29284_, _07400_);
  not _79790_ (_29316_, _29315_);
  nor _79791_ (_29317_, _29316_, _29314_);
  nor _79792_ (_29319_, _29317_, _29313_);
  nor _79793_ (_29320_, _29319_, _03222_);
  nor _79794_ (_29321_, _12519_, _10909_);
  or _79795_ (_29322_, _29284_, _03589_);
  nor _79796_ (_29323_, _29322_, _29321_);
  or _79797_ (_29324_, _29323_, _03601_);
  nor _79798_ (_29325_, _29324_, _29320_);
  and _79799_ (_29326_, _05263_, _06332_);
  nor _79800_ (_29327_, _29326_, _29284_);
  nand _79801_ (_29328_, _29327_, _07766_);
  and _79802_ (_29330_, _29328_, _08828_);
  nor _79803_ (_29331_, _29330_, _29325_);
  and _79804_ (_29332_, _12533_, _05263_);
  nor _79805_ (_29333_, _29332_, _29284_);
  and _79806_ (_29334_, _29333_, _03600_);
  nor _79807_ (_29335_, _29334_, _29331_);
  nor _79808_ (_29336_, _29335_, _03780_);
  and _79809_ (_29337_, _12539_, _05263_);
  or _79810_ (_29338_, _29284_, _07778_);
  nor _79811_ (_29339_, _29338_, _29337_);
  or _79812_ (_29341_, _29339_, _03622_);
  nor _79813_ (_29342_, _29341_, _29336_);
  nor _79814_ (_29343_, _29284_, _05718_);
  not _79815_ (_29344_, _29343_);
  nor _79816_ (_29345_, _29327_, _07777_);
  and _79817_ (_29346_, _29345_, _29344_);
  nor _79818_ (_29347_, _29346_, _29342_);
  nor _79819_ (_29348_, _29347_, _03790_);
  nor _79820_ (_29349_, _29298_, _06828_);
  and _79821_ (_29350_, _29349_, _29344_);
  or _79822_ (_29352_, _29350_, _29348_);
  and _79823_ (_29353_, _29352_, _07795_);
  nor _79824_ (_29354_, _12532_, _10909_);
  nor _79825_ (_29355_, _29354_, _29284_);
  nor _79826_ (_29356_, _29355_, _07795_);
  or _79827_ (_29357_, _29356_, _29353_);
  and _79828_ (_29358_, _29357_, _07793_);
  nor _79829_ (_29359_, _29358_, _29288_);
  nor _79830_ (_29360_, _29359_, _03815_);
  nor _79831_ (_29361_, _29293_, _04246_);
  or _79832_ (_29363_, _29361_, _03447_);
  nor _79833_ (_29364_, _29363_, _29360_);
  and _79834_ (_29365_, _12592_, _05263_);
  or _79835_ (_29366_, _29284_, _03514_);
  nor _79836_ (_29367_, _29366_, _29365_);
  nor _79837_ (_29368_, _29367_, _29364_);
  or _79838_ (_29369_, _29368_, _43004_);
  or _79839_ (_29370_, _43000_, \oc8051_golden_model_1.TH0 [2]);
  and _79840_ (_29371_, _29370_, _41806_);
  and _79841_ (_43626_, _29371_, _29369_);
  not _79842_ (_29373_, \oc8051_golden_model_1.TH0 [3]);
  nor _79843_ (_29374_, _05263_, _29373_);
  nor _79844_ (_29375_, _12738_, _10909_);
  nor _79845_ (_29376_, _29375_, _29374_);
  nor _79846_ (_29377_, _29376_, _07793_);
  and _79847_ (_29378_, _12739_, _05263_);
  nor _79848_ (_29379_, _29378_, _29374_);
  nor _79849_ (_29380_, _29379_, _07778_);
  and _79850_ (_29381_, _06592_, _05263_);
  or _79851_ (_29382_, _29381_, _29374_);
  and _79852_ (_29383_, _29382_, _04481_);
  and _79853_ (_29384_, _05263_, \oc8051_golden_model_1.ACC [3]);
  nor _79854_ (_29385_, _29384_, _29374_);
  nor _79855_ (_29386_, _29385_, _03737_);
  nor _79856_ (_29387_, _29385_, _09029_);
  nor _79857_ (_29388_, _04409_, _29373_);
  or _79858_ (_29389_, _29388_, _29387_);
  and _79859_ (_29390_, _29389_, _04081_);
  nor _79860_ (_29391_, _12627_, _10909_);
  nor _79861_ (_29392_, _29391_, _29374_);
  nor _79862_ (_29394_, _29392_, _04081_);
  or _79863_ (_29395_, _29394_, _29390_);
  and _79864_ (_29396_, _29395_, _03996_);
  nor _79865_ (_29397_, _10909_, _05005_);
  nor _79866_ (_29398_, _29397_, _29374_);
  nor _79867_ (_29399_, _29398_, _03996_);
  nor _79868_ (_29400_, _29399_, _29396_);
  nor _79869_ (_29401_, _29400_, _03729_);
  or _79870_ (_29402_, _29401_, _07390_);
  nor _79871_ (_29403_, _29402_, _29386_);
  and _79872_ (_29405_, _29398_, _07390_);
  or _79873_ (_29406_, _29405_, _04481_);
  nor _79874_ (_29407_, _29406_, _29403_);
  or _79875_ (_29408_, _29407_, _29383_);
  and _79876_ (_29409_, _29408_, _03589_);
  nor _79877_ (_29410_, _12718_, _10909_);
  nor _79878_ (_29411_, _29410_, _29374_);
  nor _79879_ (_29412_, _29411_, _03589_);
  or _79880_ (_29413_, _29412_, _08828_);
  or _79881_ (_29414_, _29413_, _29409_);
  and _79882_ (_29416_, _12733_, _05263_);
  or _79883_ (_29417_, _29374_, _07766_);
  or _79884_ (_29418_, _29417_, _29416_);
  and _79885_ (_29419_, _05263_, _06276_);
  nor _79886_ (_29420_, _29419_, _29374_);
  and _79887_ (_29421_, _29420_, _03601_);
  nor _79888_ (_29422_, _29421_, _03780_);
  and _79889_ (_29423_, _29422_, _29418_);
  and _79890_ (_29424_, _29423_, _29414_);
  nor _79891_ (_29425_, _29424_, _29380_);
  nor _79892_ (_29427_, _29425_, _03622_);
  nor _79893_ (_29428_, _29374_, _05567_);
  not _79894_ (_29429_, _29428_);
  nor _79895_ (_29430_, _29420_, _07777_);
  and _79896_ (_29431_, _29430_, _29429_);
  nor _79897_ (_29432_, _29431_, _29427_);
  nor _79898_ (_29433_, _29432_, _03790_);
  nor _79899_ (_29434_, _29385_, _06828_);
  and _79900_ (_29435_, _29434_, _29429_);
  nor _79901_ (_29436_, _29435_, _03624_);
  not _79902_ (_29438_, _29436_);
  nor _79903_ (_29439_, _29438_, _29433_);
  nor _79904_ (_29440_, _12732_, _10909_);
  or _79905_ (_29441_, _29374_, _07795_);
  nor _79906_ (_29442_, _29441_, _29440_);
  or _79907_ (_29443_, _29442_, _03785_);
  nor _79908_ (_29444_, _29443_, _29439_);
  nor _79909_ (_29445_, _29444_, _29377_);
  nor _79910_ (_29446_, _29445_, _03815_);
  nor _79911_ (_29447_, _29392_, _04246_);
  or _79912_ (_29449_, _29447_, _03447_);
  nor _79913_ (_29450_, _29449_, _29446_);
  and _79914_ (_29451_, _12794_, _05263_);
  or _79915_ (_29452_, _29374_, _03514_);
  nor _79916_ (_29453_, _29452_, _29451_);
  nor _79917_ (_29454_, _29453_, _29450_);
  or _79918_ (_29455_, _29454_, _43004_);
  or _79919_ (_29456_, _43000_, \oc8051_golden_model_1.TH0 [3]);
  and _79920_ (_29457_, _29456_, _41806_);
  and _79921_ (_43627_, _29457_, _29455_);
  not _79922_ (_29459_, \oc8051_golden_model_1.TH0 [4]);
  nor _79923_ (_29460_, _05263_, _29459_);
  nor _79924_ (_29461_, _12816_, _10909_);
  nor _79925_ (_29462_, _29461_, _29460_);
  nor _79926_ (_29463_, _29462_, _07793_);
  and _79927_ (_29464_, _12817_, _05263_);
  nor _79928_ (_29465_, _29464_, _29460_);
  nor _79929_ (_29466_, _29465_, _07778_);
  and _79930_ (_29467_, _06298_, _05263_);
  nor _79931_ (_29468_, _29467_, _29460_);
  and _79932_ (_29470_, _29468_, _03601_);
  and _79933_ (_29471_, _05263_, \oc8051_golden_model_1.ACC [4]);
  nor _79934_ (_29472_, _29471_, _29460_);
  nor _79935_ (_29473_, _29472_, _03737_);
  nor _79936_ (_29474_, _29472_, _09029_);
  nor _79937_ (_29475_, _04409_, _29459_);
  or _79938_ (_29476_, _29475_, _29474_);
  and _79939_ (_29477_, _29476_, _04081_);
  nor _79940_ (_29478_, _12841_, _10909_);
  nor _79941_ (_29479_, _29478_, _29460_);
  nor _79942_ (_29481_, _29479_, _04081_);
  or _79943_ (_29482_, _29481_, _29477_);
  and _79944_ (_29483_, _29482_, _03996_);
  nor _79945_ (_29484_, _05777_, _10909_);
  nor _79946_ (_29485_, _29484_, _29460_);
  nor _79947_ (_29486_, _29485_, _03996_);
  nor _79948_ (_29487_, _29486_, _29483_);
  nor _79949_ (_29488_, _29487_, _03729_);
  or _79950_ (_29489_, _29488_, _07390_);
  nor _79951_ (_29490_, _29489_, _29473_);
  and _79952_ (_29492_, _29485_, _07390_);
  nor _79953_ (_29493_, _29492_, _29490_);
  nor _79954_ (_29494_, _29493_, _04481_);
  and _79955_ (_29495_, _06730_, _05263_);
  nor _79956_ (_29496_, _29460_, _07400_);
  not _79957_ (_29497_, _29496_);
  nor _79958_ (_29498_, _29497_, _29495_);
  or _79959_ (_29499_, _29498_, _03222_);
  nor _79960_ (_29500_, _29499_, _29494_);
  nor _79961_ (_29501_, _12933_, _10909_);
  nor _79962_ (_29502_, _29501_, _29460_);
  nor _79963_ (_29503_, _29502_, _03589_);
  or _79964_ (_29504_, _29503_, _03601_);
  nor _79965_ (_29505_, _29504_, _29500_);
  nor _79966_ (_29506_, _29505_, _29470_);
  or _79967_ (_29507_, _29506_, _03600_);
  and _79968_ (_29508_, _12821_, _05263_);
  or _79969_ (_29509_, _29508_, _29460_);
  or _79970_ (_29510_, _29509_, _07766_);
  and _79971_ (_29511_, _29510_, _07778_);
  and _79972_ (_29514_, _29511_, _29507_);
  nor _79973_ (_29515_, _29514_, _29466_);
  nor _79974_ (_29516_, _29515_, _03622_);
  nor _79975_ (_29517_, _29460_, _05825_);
  not _79976_ (_29518_, _29517_);
  nor _79977_ (_29519_, _29468_, _07777_);
  and _79978_ (_29520_, _29519_, _29518_);
  nor _79979_ (_29521_, _29520_, _29516_);
  nor _79980_ (_29522_, _29521_, _03790_);
  nor _79981_ (_29523_, _29472_, _06828_);
  and _79982_ (_29525_, _29523_, _29518_);
  nor _79983_ (_29526_, _29525_, _03624_);
  not _79984_ (_29527_, _29526_);
  nor _79985_ (_29528_, _29527_, _29522_);
  nor _79986_ (_29529_, _12819_, _10909_);
  or _79987_ (_29530_, _29460_, _07795_);
  nor _79988_ (_29531_, _29530_, _29529_);
  or _79989_ (_29532_, _29531_, _03785_);
  nor _79990_ (_29533_, _29532_, _29528_);
  nor _79991_ (_29534_, _29533_, _29463_);
  nor _79992_ (_29536_, _29534_, _03815_);
  nor _79993_ (_29537_, _29479_, _04246_);
  or _79994_ (_29538_, _29537_, _03447_);
  nor _79995_ (_29539_, _29538_, _29536_);
  and _79996_ (_29540_, _13003_, _05263_);
  or _79997_ (_29541_, _29460_, _03514_);
  nor _79998_ (_29542_, _29541_, _29540_);
  nor _79999_ (_29543_, _29542_, _29539_);
  or _80000_ (_29544_, _29543_, _43004_);
  or _80001_ (_29545_, _43000_, \oc8051_golden_model_1.TH0 [4]);
  and _80002_ (_29547_, _29545_, _41806_);
  and _80003_ (_43628_, _29547_, _29544_);
  not _80004_ (_29548_, \oc8051_golden_model_1.TH0 [5]);
  nor _80005_ (_29549_, _05263_, _29548_);
  nor _80006_ (_29550_, _13146_, _10909_);
  nor _80007_ (_29551_, _29550_, _29549_);
  nor _80008_ (_29552_, _29551_, _07793_);
  and _80009_ (_29553_, _13147_, _05263_);
  nor _80010_ (_29554_, _29553_, _29549_);
  nor _80011_ (_29555_, _29554_, _07778_);
  and _80012_ (_29557_, _06684_, _05263_);
  or _80013_ (_29558_, _29557_, _29549_);
  and _80014_ (_29559_, _29558_, _04481_);
  and _80015_ (_29560_, _05263_, \oc8051_golden_model_1.ACC [5]);
  nor _80016_ (_29561_, _29560_, _29549_);
  nor _80017_ (_29562_, _29561_, _03737_);
  nor _80018_ (_29563_, _29561_, _09029_);
  nor _80019_ (_29564_, _04409_, _29548_);
  or _80020_ (_29565_, _29564_, _29563_);
  and _80021_ (_29566_, _29565_, _04081_);
  nor _80022_ (_29568_, _13014_, _10909_);
  nor _80023_ (_29569_, _29568_, _29549_);
  nor _80024_ (_29570_, _29569_, _04081_);
  or _80025_ (_29571_, _29570_, _29566_);
  and _80026_ (_29572_, _29571_, _03996_);
  nor _80027_ (_29573_, _05469_, _10909_);
  nor _80028_ (_29574_, _29573_, _29549_);
  nor _80029_ (_29575_, _29574_, _03996_);
  nor _80030_ (_29576_, _29575_, _29572_);
  nor _80031_ (_29577_, _29576_, _03729_);
  or _80032_ (_29579_, _29577_, _07390_);
  nor _80033_ (_29580_, _29579_, _29562_);
  and _80034_ (_29581_, _29574_, _07390_);
  or _80035_ (_29582_, _29581_, _04481_);
  nor _80036_ (_29583_, _29582_, _29580_);
  or _80037_ (_29584_, _29583_, _29559_);
  and _80038_ (_29585_, _29584_, _03589_);
  nor _80039_ (_29586_, _13127_, _10909_);
  nor _80040_ (_29587_, _29586_, _29549_);
  nor _80041_ (_29588_, _29587_, _03589_);
  or _80042_ (_29590_, _29588_, _08828_);
  or _80043_ (_29591_, _29590_, _29585_);
  and _80044_ (_29592_, _13141_, _05263_);
  or _80045_ (_29593_, _29549_, _07766_);
  or _80046_ (_29594_, _29593_, _29592_);
  and _80047_ (_29595_, _06306_, _05263_);
  nor _80048_ (_29596_, _29595_, _29549_);
  and _80049_ (_29597_, _29596_, _03601_);
  nor _80050_ (_29598_, _29597_, _03780_);
  and _80051_ (_29599_, _29598_, _29594_);
  and _80052_ (_29601_, _29599_, _29591_);
  nor _80053_ (_29602_, _29601_, _29555_);
  nor _80054_ (_29603_, _29602_, _03622_);
  nor _80055_ (_29604_, _29549_, _05518_);
  not _80056_ (_29605_, _29604_);
  nor _80057_ (_29606_, _29596_, _07777_);
  and _80058_ (_29607_, _29606_, _29605_);
  nor _80059_ (_29608_, _29607_, _29603_);
  nor _80060_ (_29609_, _29608_, _03790_);
  nor _80061_ (_29610_, _29561_, _06828_);
  and _80062_ (_29612_, _29610_, _29605_);
  or _80063_ (_29613_, _29612_, _29609_);
  and _80064_ (_29614_, _29613_, _07795_);
  nor _80065_ (_29615_, _13140_, _10909_);
  nor _80066_ (_29616_, _29615_, _29549_);
  nor _80067_ (_29617_, _29616_, _07795_);
  or _80068_ (_29618_, _29617_, _29614_);
  and _80069_ (_29619_, _29618_, _07793_);
  nor _80070_ (_29620_, _29619_, _29552_);
  nor _80071_ (_29621_, _29620_, _03815_);
  nor _80072_ (_29623_, _29569_, _04246_);
  or _80073_ (_29624_, _29623_, _03447_);
  nor _80074_ (_29625_, _29624_, _29621_);
  and _80075_ (_29626_, _13199_, _05263_);
  or _80076_ (_29627_, _29549_, _03514_);
  nor _80077_ (_29628_, _29627_, _29626_);
  nor _80078_ (_29629_, _29628_, _29625_);
  or _80079_ (_29630_, _29629_, _43004_);
  or _80080_ (_29631_, _43000_, \oc8051_golden_model_1.TH0 [5]);
  and _80081_ (_29632_, _29631_, _41806_);
  and _80082_ (_43629_, _29632_, _29630_);
  not _80083_ (_29634_, \oc8051_golden_model_1.TH0 [6]);
  nor _80084_ (_29635_, _05263_, _29634_);
  nor _80085_ (_29636_, _13352_, _10909_);
  nor _80086_ (_29637_, _29636_, _29635_);
  nor _80087_ (_29638_, _29637_, _07793_);
  and _80088_ (_29639_, _13353_, _05263_);
  nor _80089_ (_29640_, _29639_, _29635_);
  nor _80090_ (_29641_, _29640_, _07778_);
  and _80091_ (_29642_, _06455_, _05263_);
  or _80092_ (_29644_, _29642_, _29635_);
  and _80093_ (_29645_, _29644_, _04481_);
  and _80094_ (_29646_, _05263_, \oc8051_golden_model_1.ACC [6]);
  nor _80095_ (_29647_, _29646_, _29635_);
  nor _80096_ (_29648_, _29647_, _03737_);
  nor _80097_ (_29649_, _29647_, _09029_);
  nor _80098_ (_29650_, _04409_, _29634_);
  or _80099_ (_29651_, _29650_, _29649_);
  and _80100_ (_29652_, _29651_, _04081_);
  nor _80101_ (_29653_, _13242_, _10909_);
  nor _80102_ (_29655_, _29653_, _29635_);
  nor _80103_ (_29656_, _29655_, _04081_);
  or _80104_ (_29657_, _29656_, _29652_);
  and _80105_ (_29658_, _29657_, _03996_);
  nor _80106_ (_29659_, _05363_, _10909_);
  nor _80107_ (_29660_, _29659_, _29635_);
  nor _80108_ (_29661_, _29660_, _03996_);
  nor _80109_ (_29662_, _29661_, _29658_);
  nor _80110_ (_29663_, _29662_, _03729_);
  or _80111_ (_29664_, _29663_, _07390_);
  nor _80112_ (_29666_, _29664_, _29648_);
  and _80113_ (_29667_, _29660_, _07390_);
  or _80114_ (_29668_, _29667_, _04481_);
  nor _80115_ (_29669_, _29668_, _29666_);
  or _80116_ (_29670_, _29669_, _29645_);
  and _80117_ (_29671_, _29670_, _03589_);
  nor _80118_ (_29672_, _13332_, _10909_);
  nor _80119_ (_29673_, _29672_, _29635_);
  nor _80120_ (_29674_, _29673_, _03589_);
  or _80121_ (_29675_, _29674_, _08828_);
  or _80122_ (_29677_, _29675_, _29671_);
  and _80123_ (_29678_, _13347_, _05263_);
  or _80124_ (_29679_, _29635_, _07766_);
  or _80125_ (_29680_, _29679_, _29678_);
  and _80126_ (_29681_, _13339_, _05263_);
  nor _80127_ (_29682_, _29681_, _29635_);
  and _80128_ (_29683_, _29682_, _03601_);
  nor _80129_ (_29684_, _29683_, _03780_);
  and _80130_ (_29685_, _29684_, _29680_);
  and _80131_ (_29686_, _29685_, _29677_);
  nor _80132_ (_29688_, _29686_, _29641_);
  nor _80133_ (_29689_, _29688_, _03622_);
  nor _80134_ (_29690_, _29635_, _05412_);
  not _80135_ (_29691_, _29690_);
  nor _80136_ (_29692_, _29682_, _07777_);
  and _80137_ (_29693_, _29692_, _29691_);
  nor _80138_ (_29694_, _29693_, _29689_);
  nor _80139_ (_29695_, _29694_, _03790_);
  nor _80140_ (_29696_, _29647_, _06828_);
  and _80141_ (_29697_, _29696_, _29691_);
  nor _80142_ (_29699_, _29697_, _03624_);
  not _80143_ (_29700_, _29699_);
  nor _80144_ (_29701_, _29700_, _29695_);
  nor _80145_ (_29702_, _13346_, _10909_);
  or _80146_ (_29703_, _29635_, _07795_);
  nor _80147_ (_29704_, _29703_, _29702_);
  or _80148_ (_29705_, _29704_, _03785_);
  nor _80149_ (_29706_, _29705_, _29701_);
  nor _80150_ (_29707_, _29706_, _29638_);
  nor _80151_ (_29708_, _29707_, _03815_);
  nor _80152_ (_29710_, _29655_, _04246_);
  or _80153_ (_29711_, _29710_, _03447_);
  nor _80154_ (_29712_, _29711_, _29708_);
  and _80155_ (_29713_, _13402_, _05263_);
  or _80156_ (_29714_, _29635_, _03514_);
  nor _80157_ (_29715_, _29714_, _29713_);
  nor _80158_ (_29716_, _29715_, _29712_);
  or _80159_ (_29717_, _29716_, _43004_);
  or _80160_ (_29718_, _43000_, \oc8051_golden_model_1.TH0 [6]);
  and _80161_ (_29719_, _29718_, _41806_);
  and _80162_ (_43630_, _29719_, _29717_);
  not _80163_ (_29721_, \oc8051_golden_model_1.TH1 [0]);
  nor _80164_ (_29722_, _05278_, _29721_);
  nor _80165_ (_29723_, _05666_, _10991_);
  nor _80166_ (_29724_, _29723_, _29722_);
  and _80167_ (_29725_, _29724_, _17166_);
  and _80168_ (_29726_, _05278_, \oc8051_golden_model_1.ACC [0]);
  nor _80169_ (_29727_, _29726_, _29722_);
  nor _80170_ (_29728_, _29727_, _03737_);
  nor _80171_ (_29729_, _29727_, _09029_);
  nor _80172_ (_29731_, _04409_, _29721_);
  or _80173_ (_29732_, _29731_, _29729_);
  and _80174_ (_29733_, _29732_, _04081_);
  nor _80175_ (_29734_, _29724_, _04081_);
  or _80176_ (_29735_, _29734_, _29733_);
  and _80177_ (_29736_, _29735_, _03996_);
  and _80178_ (_29737_, _05278_, _04620_);
  nor _80179_ (_29738_, _29737_, _29722_);
  nor _80180_ (_29739_, _29738_, _03996_);
  nor _80181_ (_29740_, _29739_, _29736_);
  nor _80182_ (_29742_, _29740_, _03729_);
  or _80183_ (_29743_, _29742_, _07390_);
  nor _80184_ (_29744_, _29743_, _29728_);
  and _80185_ (_29745_, _29738_, _07390_);
  nor _80186_ (_29746_, _29745_, _29744_);
  nor _80187_ (_29747_, _29746_, _04481_);
  and _80188_ (_29748_, _06546_, _05278_);
  nor _80189_ (_29749_, _29722_, _07400_);
  not _80190_ (_29750_, _29749_);
  nor _80191_ (_29751_, _29750_, _29748_);
  nor _80192_ (_29753_, _29751_, _29747_);
  nor _80193_ (_29754_, _29753_, _03222_);
  nor _80194_ (_29755_, _12109_, _10991_);
  or _80195_ (_29756_, _29722_, _03589_);
  nor _80196_ (_29757_, _29756_, _29755_);
  or _80197_ (_29758_, _29757_, _03601_);
  nor _80198_ (_29759_, _29758_, _29754_);
  and _80199_ (_29760_, _05278_, _06274_);
  nor _80200_ (_29761_, _29760_, _29722_);
  nand _80201_ (_29762_, _29761_, _07766_);
  and _80202_ (_29763_, _29762_, _08828_);
  nor _80203_ (_29764_, _29763_, _29759_);
  and _80204_ (_29765_, _12124_, _05278_);
  nor _80205_ (_29766_, _29765_, _29722_);
  and _80206_ (_29767_, _29766_, _03600_);
  nor _80207_ (_29768_, _29767_, _29764_);
  nor _80208_ (_29769_, _29768_, _03780_);
  and _80209_ (_29770_, _12128_, _05278_);
  or _80210_ (_29771_, _29722_, _07778_);
  nor _80211_ (_29772_, _29771_, _29770_);
  or _80212_ (_29775_, _29772_, _03622_);
  nor _80213_ (_29776_, _29775_, _29769_);
  or _80214_ (_29777_, _29761_, _07777_);
  nor _80215_ (_29778_, _29777_, _29723_);
  nor _80216_ (_29779_, _29778_, _29776_);
  nor _80217_ (_29780_, _29779_, _03790_);
  nor _80218_ (_29781_, _29722_, _05666_);
  or _80219_ (_29782_, _29781_, _06828_);
  nor _80220_ (_29783_, _29782_, _29727_);
  or _80221_ (_29784_, _29783_, _29780_);
  and _80222_ (_29786_, _29784_, _07795_);
  nor _80223_ (_29787_, _12122_, _10991_);
  nor _80224_ (_29788_, _29787_, _29722_);
  nor _80225_ (_29789_, _29788_, _07795_);
  or _80226_ (_29790_, _29789_, _29786_);
  and _80227_ (_29791_, _29790_, _07793_);
  nor _80228_ (_29792_, _12003_, _10991_);
  nor _80229_ (_29793_, _29792_, _29722_);
  nor _80230_ (_29794_, _29793_, _07793_);
  nor _80231_ (_29795_, _29794_, _17166_);
  not _80232_ (_29797_, _29795_);
  nor _80233_ (_29798_, _29797_, _29791_);
  nor _80234_ (_29799_, _29798_, _29725_);
  or _80235_ (_29800_, _29799_, _43004_);
  or _80236_ (_29801_, _43000_, \oc8051_golden_model_1.TH1 [0]);
  and _80237_ (_29802_, _29801_, _41806_);
  and _80238_ (_43631_, _29802_, _29800_);
  and _80239_ (_29803_, _06501_, _05278_);
  not _80240_ (_29804_, \oc8051_golden_model_1.TH1 [1]);
  nor _80241_ (_29805_, _05278_, _29804_);
  nor _80242_ (_29807_, _29805_, _07400_);
  not _80243_ (_29808_, _29807_);
  nor _80244_ (_29809_, _29808_, _29803_);
  not _80245_ (_29810_, _29809_);
  and _80246_ (_29811_, _05278_, _06764_);
  or _80247_ (_29812_, _29805_, _25480_);
  nor _80248_ (_29813_, _29812_, _29811_);
  nor _80249_ (_29814_, _05278_, \oc8051_golden_model_1.TH1 [1]);
  and _80250_ (_29815_, _05278_, _03274_);
  nor _80251_ (_29816_, _29815_, _29814_);
  and _80252_ (_29818_, _29816_, _03729_);
  nor _80253_ (_29819_, _29818_, _07390_);
  and _80254_ (_29820_, _12213_, _05278_);
  nor _80255_ (_29821_, _29820_, _29814_);
  and _80256_ (_29822_, _29821_, _03610_);
  and _80257_ (_29823_, _29816_, _04409_);
  nor _80258_ (_29824_, _04409_, _29804_);
  nor _80259_ (_29825_, _29824_, _29823_);
  nor _80260_ (_29826_, _29825_, _03610_);
  or _80261_ (_29827_, _29826_, _03723_);
  nor _80262_ (_29829_, _29827_, _29822_);
  or _80263_ (_29830_, _29829_, _03729_);
  and _80264_ (_29831_, _29830_, _29819_);
  nor _80265_ (_29832_, _29831_, _29813_);
  nor _80266_ (_29833_, _29832_, _04481_);
  nor _80267_ (_29834_, _29833_, _03222_);
  and _80268_ (_29835_, _29834_, _29810_);
  not _80269_ (_29836_, _29814_);
  and _80270_ (_29837_, _12313_, _05278_);
  nor _80271_ (_29838_, _29837_, _03589_);
  and _80272_ (_29840_, _29838_, _29836_);
  nor _80273_ (_29841_, _29840_, _29835_);
  nor _80274_ (_29842_, _29841_, _08828_);
  nor _80275_ (_29843_, _12327_, _10991_);
  nor _80276_ (_29844_, _29843_, _07766_);
  and _80277_ (_29845_, _05278_, _04303_);
  nor _80278_ (_29846_, _29845_, _05886_);
  nor _80279_ (_29847_, _29846_, _29844_);
  nor _80280_ (_29848_, _29847_, _29814_);
  nor _80281_ (_29849_, _29848_, _29842_);
  nor _80282_ (_29851_, _29849_, _03780_);
  nor _80283_ (_29852_, _12333_, _10991_);
  nor _80284_ (_29853_, _29852_, _07778_);
  and _80285_ (_29854_, _29853_, _29836_);
  nor _80286_ (_29855_, _29854_, _29851_);
  nor _80287_ (_29856_, _29855_, _03622_);
  nor _80288_ (_29857_, _12207_, _10991_);
  nor _80289_ (_29858_, _29857_, _07777_);
  and _80290_ (_29859_, _29858_, _29836_);
  nor _80291_ (_29860_, _29859_, _29856_);
  nor _80292_ (_29862_, _29860_, _03790_);
  nor _80293_ (_29863_, _29805_, _05618_);
  nor _80294_ (_29864_, _29863_, _06828_);
  and _80295_ (_29865_, _29864_, _29816_);
  nor _80296_ (_29866_, _29865_, _29862_);
  or _80297_ (_29867_, _29866_, _18499_);
  nand _80298_ (_29868_, _29815_, _05617_);
  nor _80299_ (_29869_, _29814_, _07793_);
  and _80300_ (_29870_, _29869_, _29868_);
  nor _80301_ (_29871_, _29870_, _03815_);
  and _80302_ (_29873_, _29845_, _05617_);
  or _80303_ (_29874_, _29814_, _07795_);
  or _80304_ (_29875_, _29874_, _29873_);
  and _80305_ (_29876_, _29875_, _29871_);
  and _80306_ (_29877_, _29876_, _29867_);
  nor _80307_ (_29878_, _29821_, _04246_);
  nor _80308_ (_29879_, _29878_, _29877_);
  and _80309_ (_29880_, _29879_, _03514_);
  nor _80310_ (_29881_, _29820_, _29805_);
  nor _80311_ (_29882_, _29881_, _03514_);
  or _80312_ (_29884_, _29882_, _29880_);
  or _80313_ (_29885_, _29884_, _43004_);
  or _80314_ (_29886_, _43000_, \oc8051_golden_model_1.TH1 [1]);
  and _80315_ (_29887_, _29886_, _41806_);
  and _80316_ (_43632_, _29887_, _29885_);
  not _80317_ (_29888_, \oc8051_golden_model_1.TH1 [2]);
  nor _80318_ (_29889_, _05278_, _29888_);
  nor _80319_ (_29890_, _12538_, _10991_);
  nor _80320_ (_29891_, _29890_, _29889_);
  nor _80321_ (_29892_, _29891_, _07793_);
  and _80322_ (_29894_, _12539_, _05278_);
  nor _80323_ (_29895_, _29894_, _29889_);
  nor _80324_ (_29896_, _29895_, _07778_);
  and _80325_ (_29897_, _05278_, \oc8051_golden_model_1.ACC [2]);
  nor _80326_ (_29898_, _29897_, _29889_);
  nor _80327_ (_29899_, _29898_, _03737_);
  nor _80328_ (_29900_, _29898_, _09029_);
  nor _80329_ (_29901_, _04409_, _29888_);
  or _80330_ (_29902_, _29901_, _29900_);
  and _80331_ (_29903_, _29902_, _04081_);
  nor _80332_ (_29905_, _12416_, _10991_);
  nor _80333_ (_29906_, _29905_, _29889_);
  nor _80334_ (_29907_, _29906_, _04081_);
  or _80335_ (_29908_, _29907_, _29903_);
  and _80336_ (_29909_, _29908_, _03996_);
  nor _80337_ (_29910_, _10991_, _04875_);
  nor _80338_ (_29911_, _29910_, _29889_);
  nor _80339_ (_29912_, _29911_, _03996_);
  nor _80340_ (_29913_, _29912_, _29909_);
  nor _80341_ (_29914_, _29913_, _03729_);
  or _80342_ (_29916_, _29914_, _07390_);
  nor _80343_ (_29917_, _29916_, _29899_);
  and _80344_ (_29918_, _29911_, _07390_);
  nor _80345_ (_29919_, _29918_, _29917_);
  nor _80346_ (_29920_, _29919_, _04481_);
  and _80347_ (_29921_, _06637_, _05278_);
  nor _80348_ (_29922_, _29889_, _07400_);
  not _80349_ (_29923_, _29922_);
  nor _80350_ (_29924_, _29923_, _29921_);
  nor _80351_ (_29925_, _29924_, _03222_);
  not _80352_ (_29927_, _29925_);
  nor _80353_ (_29928_, _29927_, _29920_);
  nor _80354_ (_29929_, _12519_, _10991_);
  nor _80355_ (_29930_, _29929_, _29889_);
  nor _80356_ (_29931_, _29930_, _03589_);
  or _80357_ (_29932_, _29931_, _08828_);
  or _80358_ (_29933_, _29932_, _29928_);
  and _80359_ (_29934_, _12533_, _05278_);
  or _80360_ (_29935_, _29889_, _07766_);
  or _80361_ (_29936_, _29935_, _29934_);
  and _80362_ (_29938_, _05278_, _06332_);
  nor _80363_ (_29939_, _29938_, _29889_);
  and _80364_ (_29940_, _29939_, _03601_);
  nor _80365_ (_29941_, _29940_, _03780_);
  and _80366_ (_29942_, _29941_, _29936_);
  and _80367_ (_29943_, _29942_, _29933_);
  nor _80368_ (_29944_, _29943_, _29896_);
  nor _80369_ (_29945_, _29944_, _03622_);
  nor _80370_ (_29946_, _29889_, _05718_);
  not _80371_ (_29947_, _29946_);
  nor _80372_ (_29949_, _29939_, _07777_);
  and _80373_ (_29950_, _29949_, _29947_);
  nor _80374_ (_29951_, _29950_, _29945_);
  nor _80375_ (_29952_, _29951_, _03790_);
  nor _80376_ (_29953_, _29898_, _06828_);
  and _80377_ (_29954_, _29953_, _29947_);
  or _80378_ (_29955_, _29954_, _29952_);
  and _80379_ (_29956_, _29955_, _07795_);
  nor _80380_ (_29957_, _12532_, _10991_);
  nor _80381_ (_29958_, _29957_, _29889_);
  nor _80382_ (_29960_, _29958_, _07795_);
  or _80383_ (_29961_, _29960_, _29956_);
  and _80384_ (_29962_, _29961_, _07793_);
  nor _80385_ (_29963_, _29962_, _29892_);
  nor _80386_ (_29964_, _29963_, _03815_);
  nor _80387_ (_29965_, _29906_, _04246_);
  or _80388_ (_29966_, _29965_, _03447_);
  nor _80389_ (_29967_, _29966_, _29964_);
  and _80390_ (_29968_, _12592_, _05278_);
  or _80391_ (_29969_, _29889_, _03514_);
  nor _80392_ (_29971_, _29969_, _29968_);
  nor _80393_ (_29972_, _29971_, _29967_);
  or _80394_ (_29973_, _29972_, _43004_);
  or _80395_ (_29974_, _43000_, \oc8051_golden_model_1.TH1 [2]);
  and _80396_ (_29975_, _29974_, _41806_);
  and _80397_ (_43633_, _29975_, _29973_);
  not _80398_ (_29976_, \oc8051_golden_model_1.TH1 [3]);
  nor _80399_ (_29977_, _05278_, _29976_);
  nor _80400_ (_29978_, _12738_, _10991_);
  nor _80401_ (_29979_, _29978_, _29977_);
  nor _80402_ (_29981_, _29979_, _07793_);
  and _80403_ (_29982_, _12739_, _05278_);
  nor _80404_ (_29983_, _29982_, _29977_);
  nor _80405_ (_29984_, _29983_, _07778_);
  and _80406_ (_29985_, _06592_, _05278_);
  or _80407_ (_29986_, _29985_, _29977_);
  and _80408_ (_29987_, _29986_, _04481_);
  and _80409_ (_29988_, _05278_, \oc8051_golden_model_1.ACC [3]);
  nor _80410_ (_29989_, _29988_, _29977_);
  nor _80411_ (_29990_, _29989_, _03737_);
  nor _80412_ (_29992_, _29989_, _09029_);
  nor _80413_ (_29993_, _04409_, _29976_);
  or _80414_ (_29994_, _29993_, _29992_);
  and _80415_ (_29995_, _29994_, _04081_);
  nor _80416_ (_29996_, _12627_, _10991_);
  nor _80417_ (_29997_, _29996_, _29977_);
  nor _80418_ (_29998_, _29997_, _04081_);
  or _80419_ (_29999_, _29998_, _29995_);
  and _80420_ (_30000_, _29999_, _03996_);
  nor _80421_ (_30001_, _10991_, _05005_);
  nor _80422_ (_30003_, _30001_, _29977_);
  nor _80423_ (_30004_, _30003_, _03996_);
  nor _80424_ (_30005_, _30004_, _30000_);
  nor _80425_ (_30006_, _30005_, _03729_);
  or _80426_ (_30007_, _30006_, _07390_);
  nor _80427_ (_30008_, _30007_, _29990_);
  and _80428_ (_30009_, _30003_, _07390_);
  or _80429_ (_30010_, _30009_, _04481_);
  nor _80430_ (_30011_, _30010_, _30008_);
  or _80431_ (_30012_, _30011_, _29987_);
  and _80432_ (_30014_, _30012_, _03589_);
  nor _80433_ (_30015_, _12718_, _10991_);
  nor _80434_ (_30016_, _30015_, _29977_);
  nor _80435_ (_30017_, _30016_, _03589_);
  or _80436_ (_30018_, _30017_, _08828_);
  or _80437_ (_30019_, _30018_, _30014_);
  and _80438_ (_30020_, _12733_, _05278_);
  or _80439_ (_30021_, _29977_, _07766_);
  or _80440_ (_30022_, _30021_, _30020_);
  and _80441_ (_30023_, _05278_, _06276_);
  nor _80442_ (_30025_, _30023_, _29977_);
  and _80443_ (_30026_, _30025_, _03601_);
  nor _80444_ (_30027_, _30026_, _03780_);
  and _80445_ (_30028_, _30027_, _30022_);
  and _80446_ (_30029_, _30028_, _30019_);
  nor _80447_ (_30030_, _30029_, _29984_);
  nor _80448_ (_30031_, _30030_, _03622_);
  nor _80449_ (_30032_, _29977_, _05567_);
  not _80450_ (_30033_, _30032_);
  nor _80451_ (_30034_, _30025_, _07777_);
  and _80452_ (_30036_, _30034_, _30033_);
  nor _80453_ (_30037_, _30036_, _30031_);
  nor _80454_ (_30038_, _30037_, _03790_);
  nor _80455_ (_30039_, _29989_, _06828_);
  and _80456_ (_30040_, _30039_, _30033_);
  or _80457_ (_30041_, _30040_, _30038_);
  and _80458_ (_30042_, _30041_, _07795_);
  nor _80459_ (_30043_, _12732_, _10991_);
  nor _80460_ (_30044_, _30043_, _29977_);
  nor _80461_ (_30045_, _30044_, _07795_);
  or _80462_ (_30047_, _30045_, _30042_);
  and _80463_ (_30048_, _30047_, _07793_);
  nor _80464_ (_30049_, _30048_, _29981_);
  nor _80465_ (_30050_, _30049_, _03815_);
  nor _80466_ (_30051_, _29997_, _04246_);
  or _80467_ (_30052_, _30051_, _03447_);
  nor _80468_ (_30053_, _30052_, _30050_);
  and _80469_ (_30054_, _12794_, _05278_);
  or _80470_ (_30055_, _29977_, _03514_);
  nor _80471_ (_30056_, _30055_, _30054_);
  nor _80472_ (_30058_, _30056_, _30053_);
  or _80473_ (_30059_, _30058_, _43004_);
  or _80474_ (_30060_, _43000_, \oc8051_golden_model_1.TH1 [3]);
  and _80475_ (_30061_, _30060_, _41806_);
  and _80476_ (_43634_, _30061_, _30059_);
  not _80477_ (_30062_, \oc8051_golden_model_1.TH1 [4]);
  nor _80478_ (_30063_, _05278_, _30062_);
  nor _80479_ (_30064_, _12816_, _10991_);
  nor _80480_ (_30065_, _30064_, _30063_);
  nor _80481_ (_30066_, _30065_, _07793_);
  and _80482_ (_30067_, _12817_, _05278_);
  nor _80483_ (_30068_, _30067_, _30063_);
  nor _80484_ (_30069_, _30068_, _07778_);
  and _80485_ (_30070_, _06298_, _05278_);
  nor _80486_ (_30071_, _30070_, _30063_);
  and _80487_ (_30072_, _30071_, _03601_);
  nor _80488_ (_30073_, _05777_, _10991_);
  nor _80489_ (_30074_, _30073_, _30063_);
  and _80490_ (_30075_, _30074_, _07390_);
  and _80491_ (_30076_, _05278_, \oc8051_golden_model_1.ACC [4]);
  nor _80492_ (_30079_, _30076_, _30063_);
  nor _80493_ (_30080_, _30079_, _03737_);
  nor _80494_ (_30081_, _30079_, _09029_);
  nor _80495_ (_30082_, _04409_, _30062_);
  or _80496_ (_30083_, _30082_, _30081_);
  and _80497_ (_30084_, _30083_, _04081_);
  nor _80498_ (_30085_, _12841_, _10991_);
  nor _80499_ (_30086_, _30085_, _30063_);
  nor _80500_ (_30087_, _30086_, _04081_);
  or _80501_ (_30088_, _30087_, _30084_);
  and _80502_ (_30089_, _30088_, _03996_);
  nor _80503_ (_30090_, _30074_, _03996_);
  nor _80504_ (_30091_, _30090_, _30089_);
  nor _80505_ (_30092_, _30091_, _03729_);
  or _80506_ (_30093_, _30092_, _07390_);
  nor _80507_ (_30094_, _30093_, _30080_);
  nor _80508_ (_30095_, _30094_, _30075_);
  nor _80509_ (_30096_, _30095_, _04481_);
  and _80510_ (_30097_, _06730_, _05278_);
  nor _80511_ (_30098_, _30063_, _07400_);
  not _80512_ (_30100_, _30098_);
  nor _80513_ (_30101_, _30100_, _30097_);
  or _80514_ (_30102_, _30101_, _03222_);
  nor _80515_ (_30103_, _30102_, _30096_);
  nor _80516_ (_30104_, _12933_, _10991_);
  nor _80517_ (_30105_, _30104_, _30063_);
  nor _80518_ (_30106_, _30105_, _03589_);
  or _80519_ (_30107_, _30106_, _03601_);
  nor _80520_ (_30108_, _30107_, _30103_);
  nor _80521_ (_30109_, _30108_, _30072_);
  or _80522_ (_30111_, _30109_, _03600_);
  and _80523_ (_30112_, _12821_, _05278_);
  or _80524_ (_30113_, _30112_, _30063_);
  or _80525_ (_30114_, _30113_, _07766_);
  and _80526_ (_30115_, _30114_, _07778_);
  and _80527_ (_30116_, _30115_, _30111_);
  nor _80528_ (_30117_, _30116_, _30069_);
  nor _80529_ (_30118_, _30117_, _03622_);
  nor _80530_ (_30119_, _30063_, _05825_);
  not _80531_ (_30120_, _30119_);
  nor _80532_ (_30122_, _30071_, _07777_);
  and _80533_ (_30123_, _30122_, _30120_);
  nor _80534_ (_30124_, _30123_, _30118_);
  nor _80535_ (_30125_, _30124_, _03790_);
  nor _80536_ (_30126_, _30079_, _06828_);
  and _80537_ (_30127_, _30126_, _30120_);
  nor _80538_ (_30128_, _30127_, _03624_);
  not _80539_ (_30129_, _30128_);
  nor _80540_ (_30130_, _30129_, _30125_);
  nor _80541_ (_30131_, _12819_, _10991_);
  or _80542_ (_30133_, _30063_, _07795_);
  nor _80543_ (_30134_, _30133_, _30131_);
  or _80544_ (_30135_, _30134_, _03785_);
  nor _80545_ (_30136_, _30135_, _30130_);
  nor _80546_ (_30137_, _30136_, _30066_);
  nor _80547_ (_30138_, _30137_, _03815_);
  nor _80548_ (_30139_, _30086_, _04246_);
  or _80549_ (_30140_, _30139_, _03447_);
  nor _80550_ (_30141_, _30140_, _30138_);
  and _80551_ (_30142_, _13003_, _05278_);
  or _80552_ (_30144_, _30063_, _03514_);
  nor _80553_ (_30145_, _30144_, _30142_);
  nor _80554_ (_30146_, _30145_, _30141_);
  or _80555_ (_30147_, _30146_, _43004_);
  or _80556_ (_30148_, _43000_, \oc8051_golden_model_1.TH1 [4]);
  and _80557_ (_30149_, _30148_, _41806_);
  and _80558_ (_43635_, _30149_, _30147_);
  not _80559_ (_30150_, \oc8051_golden_model_1.TH1 [5]);
  nor _80560_ (_30151_, _05278_, _30150_);
  nor _80561_ (_30152_, _13146_, _10991_);
  nor _80562_ (_30154_, _30152_, _30151_);
  nor _80563_ (_30155_, _30154_, _07793_);
  and _80564_ (_30156_, _13147_, _05278_);
  nor _80565_ (_30157_, _30156_, _30151_);
  nor _80566_ (_30158_, _30157_, _07778_);
  and _80567_ (_30159_, _06684_, _05278_);
  or _80568_ (_30160_, _30159_, _30151_);
  and _80569_ (_30161_, _30160_, _04481_);
  and _80570_ (_30162_, _05278_, \oc8051_golden_model_1.ACC [5]);
  nor _80571_ (_30163_, _30162_, _30151_);
  nor _80572_ (_30165_, _30163_, _03737_);
  nor _80573_ (_30166_, _30163_, _09029_);
  nor _80574_ (_30167_, _04409_, _30150_);
  or _80575_ (_30168_, _30167_, _30166_);
  and _80576_ (_30169_, _30168_, _04081_);
  nor _80577_ (_30170_, _13014_, _10991_);
  nor _80578_ (_30171_, _30170_, _30151_);
  nor _80579_ (_30172_, _30171_, _04081_);
  or _80580_ (_30173_, _30172_, _30169_);
  and _80581_ (_30174_, _30173_, _03996_);
  nor _80582_ (_30176_, _05469_, _10991_);
  nor _80583_ (_30177_, _30176_, _30151_);
  nor _80584_ (_30178_, _30177_, _03996_);
  nor _80585_ (_30179_, _30178_, _30174_);
  nor _80586_ (_30180_, _30179_, _03729_);
  or _80587_ (_30181_, _30180_, _07390_);
  nor _80588_ (_30182_, _30181_, _30165_);
  and _80589_ (_30183_, _30177_, _07390_);
  or _80590_ (_30184_, _30183_, _04481_);
  nor _80591_ (_30185_, _30184_, _30182_);
  or _80592_ (_30187_, _30185_, _30161_);
  and _80593_ (_30188_, _30187_, _03589_);
  nor _80594_ (_30189_, _13127_, _10991_);
  nor _80595_ (_30190_, _30189_, _30151_);
  nor _80596_ (_30191_, _30190_, _03589_);
  or _80597_ (_30192_, _30191_, _08828_);
  or _80598_ (_30193_, _30192_, _30188_);
  and _80599_ (_30194_, _13141_, _05278_);
  or _80600_ (_30195_, _30151_, _07766_);
  or _80601_ (_30196_, _30195_, _30194_);
  and _80602_ (_30198_, _06306_, _05278_);
  nor _80603_ (_30199_, _30198_, _30151_);
  and _80604_ (_30200_, _30199_, _03601_);
  nor _80605_ (_30201_, _30200_, _03780_);
  and _80606_ (_30202_, _30201_, _30196_);
  and _80607_ (_30203_, _30202_, _30193_);
  nor _80608_ (_30204_, _30203_, _30158_);
  nor _80609_ (_30205_, _30204_, _03622_);
  nor _80610_ (_30206_, _30151_, _05518_);
  not _80611_ (_30207_, _30206_);
  nor _80612_ (_30209_, _30199_, _07777_);
  and _80613_ (_30210_, _30209_, _30207_);
  nor _80614_ (_30211_, _30210_, _30205_);
  nor _80615_ (_30212_, _30211_, _03790_);
  nor _80616_ (_30213_, _30163_, _06828_);
  and _80617_ (_30214_, _30213_, _30207_);
  nor _80618_ (_30215_, _30214_, _03624_);
  not _80619_ (_30216_, _30215_);
  nor _80620_ (_30217_, _30216_, _30212_);
  nor _80621_ (_30218_, _13140_, _10991_);
  or _80622_ (_30220_, _30151_, _07795_);
  nor _80623_ (_30221_, _30220_, _30218_);
  or _80624_ (_30222_, _30221_, _03785_);
  nor _80625_ (_30223_, _30222_, _30217_);
  nor _80626_ (_30224_, _30223_, _30155_);
  nor _80627_ (_30225_, _30224_, _03815_);
  nor _80628_ (_30226_, _30171_, _04246_);
  or _80629_ (_30227_, _30226_, _03447_);
  nor _80630_ (_30228_, _30227_, _30225_);
  and _80631_ (_30229_, _13199_, _05278_);
  or _80632_ (_30231_, _30151_, _03514_);
  nor _80633_ (_30232_, _30231_, _30229_);
  nor _80634_ (_30233_, _30232_, _30228_);
  or _80635_ (_30234_, _30233_, _43004_);
  or _80636_ (_30235_, _43000_, \oc8051_golden_model_1.TH1 [5]);
  and _80637_ (_30236_, _30235_, _41806_);
  and _80638_ (_43638_, _30236_, _30234_);
  not _80639_ (_30237_, \oc8051_golden_model_1.TH1 [6]);
  nor _80640_ (_30238_, _05278_, _30237_);
  nor _80641_ (_30239_, _13352_, _10991_);
  nor _80642_ (_30241_, _30239_, _30238_);
  nor _80643_ (_30242_, _30241_, _07793_);
  and _80644_ (_30243_, _13353_, _05278_);
  nor _80645_ (_30244_, _30243_, _30238_);
  nor _80646_ (_30245_, _30244_, _07778_);
  and _80647_ (_30246_, _06455_, _05278_);
  or _80648_ (_30247_, _30246_, _30238_);
  and _80649_ (_30248_, _30247_, _04481_);
  and _80650_ (_30249_, _05278_, \oc8051_golden_model_1.ACC [6]);
  nor _80651_ (_30250_, _30249_, _30238_);
  nor _80652_ (_30252_, _30250_, _03737_);
  nor _80653_ (_30253_, _30250_, _09029_);
  nor _80654_ (_30254_, _04409_, _30237_);
  or _80655_ (_30255_, _30254_, _30253_);
  and _80656_ (_30256_, _30255_, _04081_);
  nor _80657_ (_30257_, _13242_, _10991_);
  nor _80658_ (_30258_, _30257_, _30238_);
  nor _80659_ (_30259_, _30258_, _04081_);
  or _80660_ (_30260_, _30259_, _30256_);
  and _80661_ (_30261_, _30260_, _03996_);
  nor _80662_ (_30263_, _05363_, _10991_);
  nor _80663_ (_30264_, _30263_, _30238_);
  nor _80664_ (_30265_, _30264_, _03996_);
  nor _80665_ (_30266_, _30265_, _30261_);
  nor _80666_ (_30267_, _30266_, _03729_);
  or _80667_ (_30268_, _30267_, _07390_);
  nor _80668_ (_30269_, _30268_, _30252_);
  and _80669_ (_30270_, _30264_, _07390_);
  or _80670_ (_30271_, _30270_, _04481_);
  nor _80671_ (_30272_, _30271_, _30269_);
  or _80672_ (_30274_, _30272_, _30248_);
  and _80673_ (_30275_, _30274_, _03589_);
  nor _80674_ (_30276_, _13332_, _10991_);
  nor _80675_ (_30277_, _30276_, _30238_);
  nor _80676_ (_30278_, _30277_, _03589_);
  or _80677_ (_30279_, _30278_, _08828_);
  or _80678_ (_30280_, _30279_, _30275_);
  and _80679_ (_30281_, _13347_, _05278_);
  or _80680_ (_30282_, _30238_, _07766_);
  or _80681_ (_30283_, _30282_, _30281_);
  and _80682_ (_30285_, _13339_, _05278_);
  nor _80683_ (_30286_, _30285_, _30238_);
  and _80684_ (_30287_, _30286_, _03601_);
  nor _80685_ (_30288_, _30287_, _03780_);
  and _80686_ (_30289_, _30288_, _30283_);
  and _80687_ (_30290_, _30289_, _30280_);
  nor _80688_ (_30291_, _30290_, _30245_);
  nor _80689_ (_30292_, _30291_, _03622_);
  nor _80690_ (_30293_, _30238_, _05412_);
  not _80691_ (_30294_, _30293_);
  nor _80692_ (_30296_, _30286_, _07777_);
  and _80693_ (_30297_, _30296_, _30294_);
  nor _80694_ (_30298_, _30297_, _30292_);
  nor _80695_ (_30299_, _30298_, _03790_);
  nor _80696_ (_30300_, _30250_, _06828_);
  and _80697_ (_30301_, _30300_, _30294_);
  or _80698_ (_30302_, _30301_, _30299_);
  and _80699_ (_30303_, _30302_, _07795_);
  nor _80700_ (_30304_, _13346_, _10991_);
  nor _80701_ (_30305_, _30304_, _30238_);
  nor _80702_ (_30307_, _30305_, _07795_);
  or _80703_ (_30308_, _30307_, _30303_);
  and _80704_ (_30309_, _30308_, _07793_);
  nor _80705_ (_30310_, _30309_, _30242_);
  nor _80706_ (_30311_, _30310_, _03815_);
  nor _80707_ (_30312_, _30258_, _04246_);
  or _80708_ (_30313_, _30312_, _03447_);
  nor _80709_ (_30314_, _30313_, _30311_);
  and _80710_ (_30315_, _13402_, _05278_);
  or _80711_ (_30316_, _30238_, _03514_);
  nor _80712_ (_30318_, _30316_, _30315_);
  nor _80713_ (_30319_, _30318_, _30314_);
  or _80714_ (_30320_, _30319_, _43004_);
  or _80715_ (_30321_, _43000_, \oc8051_golden_model_1.TH1 [6]);
  and _80716_ (_30322_, _30321_, _41806_);
  and _80717_ (_43639_, _30322_, _30320_);
  not _80718_ (_30323_, \oc8051_golden_model_1.TL0 [0]);
  nor _80719_ (_30324_, _05284_, _30323_);
  nor _80720_ (_30325_, _05666_, _11072_);
  nor _80721_ (_30326_, _30325_, _30324_);
  and _80722_ (_30328_, _30326_, _17166_);
  and _80723_ (_30329_, _05284_, \oc8051_golden_model_1.ACC [0]);
  nor _80724_ (_30330_, _30329_, _30324_);
  nor _80725_ (_30331_, _30330_, _03737_);
  nor _80726_ (_30332_, _30331_, _07390_);
  nor _80727_ (_30333_, _30326_, _04081_);
  nor _80728_ (_30334_, _04409_, _30323_);
  nor _80729_ (_30335_, _30330_, _09029_);
  nor _80730_ (_30336_, _30335_, _30334_);
  nor _80731_ (_30337_, _30336_, _03610_);
  or _80732_ (_30339_, _30337_, _03723_);
  nor _80733_ (_30340_, _30339_, _30333_);
  or _80734_ (_30341_, _30340_, _03729_);
  and _80735_ (_30342_, _30341_, _30332_);
  and _80736_ (_30343_, _05284_, _04620_);
  or _80737_ (_30344_, _30324_, _25480_);
  nor _80738_ (_30345_, _30344_, _30343_);
  nor _80739_ (_30346_, _30345_, _30342_);
  nor _80740_ (_30347_, _30346_, _04481_);
  and _80741_ (_30348_, _06546_, _05284_);
  nor _80742_ (_30350_, _30324_, _07400_);
  not _80743_ (_30351_, _30350_);
  nor _80744_ (_30352_, _30351_, _30348_);
  nor _80745_ (_30353_, _30352_, _30347_);
  nor _80746_ (_30354_, _30353_, _03222_);
  nor _80747_ (_30355_, _12109_, _11072_);
  or _80748_ (_30356_, _30324_, _03589_);
  nor _80749_ (_30357_, _30356_, _30355_);
  or _80750_ (_30358_, _30357_, _03601_);
  nor _80751_ (_30359_, _30358_, _30354_);
  and _80752_ (_30361_, _05284_, _06274_);
  nor _80753_ (_30362_, _30361_, _30324_);
  nor _80754_ (_30363_, _30362_, _05886_);
  or _80755_ (_30364_, _30363_, _30359_);
  and _80756_ (_30365_, _30364_, _07766_);
  and _80757_ (_30366_, _12124_, _05284_);
  nor _80758_ (_30367_, _30366_, _30324_);
  nor _80759_ (_30368_, _30367_, _07766_);
  or _80760_ (_30369_, _30368_, _30365_);
  nor _80761_ (_30370_, _30369_, _03780_);
  and _80762_ (_30372_, _12128_, _05284_);
  or _80763_ (_30373_, _30324_, _07778_);
  nor _80764_ (_30374_, _30373_, _30372_);
  or _80765_ (_30375_, _30374_, _03622_);
  nor _80766_ (_30376_, _30375_, _30370_);
  or _80767_ (_30377_, _30362_, _07777_);
  nor _80768_ (_30378_, _30377_, _30325_);
  nor _80769_ (_30379_, _30378_, _30376_);
  nor _80770_ (_30380_, _30379_, _03790_);
  nor _80771_ (_30381_, _30324_, _05666_);
  or _80772_ (_30383_, _30381_, _06828_);
  nor _80773_ (_30384_, _30383_, _30330_);
  or _80774_ (_30385_, _30384_, _30380_);
  and _80775_ (_30386_, _30385_, _07795_);
  nor _80776_ (_30387_, _12122_, _11072_);
  nor _80777_ (_30388_, _30387_, _30324_);
  nor _80778_ (_30389_, _30388_, _07795_);
  or _80779_ (_30390_, _30389_, _30386_);
  and _80780_ (_30391_, _30390_, _07793_);
  nor _80781_ (_30392_, _12003_, _11072_);
  nor _80782_ (_30393_, _30392_, _30324_);
  nor _80783_ (_30394_, _30393_, _07793_);
  nor _80784_ (_30395_, _30394_, _17166_);
  not _80785_ (_30396_, _30395_);
  nor _80786_ (_30397_, _30396_, _30391_);
  nor _80787_ (_30398_, _30397_, _30328_);
  or _80788_ (_30399_, _30398_, _43004_);
  or _80789_ (_30400_, _43000_, \oc8051_golden_model_1.TL0 [0]);
  and _80790_ (_30401_, _30400_, _41806_);
  and _80791_ (_43640_, _30401_, _30399_);
  and _80792_ (_30404_, _06501_, _05284_);
  not _80793_ (_30405_, \oc8051_golden_model_1.TL0 [1]);
  nor _80794_ (_30406_, _05284_, _30405_);
  nor _80795_ (_30407_, _30406_, _07400_);
  not _80796_ (_30408_, _30407_);
  nor _80797_ (_30409_, _30408_, _30404_);
  not _80798_ (_30410_, _30409_);
  and _80799_ (_30411_, _05284_, _06764_);
  nor _80800_ (_30412_, _30411_, _30406_);
  and _80801_ (_30413_, _30412_, _07390_);
  nor _80802_ (_30415_, _05284_, \oc8051_golden_model_1.TL0 [1]);
  and _80803_ (_30416_, _05284_, _03274_);
  nor _80804_ (_30417_, _30416_, _30415_);
  and _80805_ (_30418_, _30417_, _03729_);
  and _80806_ (_30419_, _30417_, _04409_);
  nor _80807_ (_30420_, _04409_, _30405_);
  or _80808_ (_30421_, _30420_, _30419_);
  and _80809_ (_30422_, _30421_, _04081_);
  and _80810_ (_30423_, _12213_, _05284_);
  nor _80811_ (_30424_, _30423_, _30415_);
  and _80812_ (_30426_, _30424_, _03610_);
  or _80813_ (_30427_, _30426_, _30422_);
  and _80814_ (_30428_, _30427_, _03996_);
  nor _80815_ (_30429_, _30412_, _03996_);
  nor _80816_ (_30430_, _30429_, _30428_);
  nor _80817_ (_30431_, _30430_, _03729_);
  or _80818_ (_30432_, _30431_, _07390_);
  nor _80819_ (_30433_, _30432_, _30418_);
  nor _80820_ (_30434_, _30433_, _30413_);
  nor _80821_ (_30435_, _30434_, _04481_);
  nor _80822_ (_30437_, _30435_, _03222_);
  and _80823_ (_30438_, _30437_, _30410_);
  not _80824_ (_30439_, _30415_);
  and _80825_ (_30440_, _12313_, _05284_);
  nor _80826_ (_30441_, _30440_, _03589_);
  and _80827_ (_30442_, _30441_, _30439_);
  nor _80828_ (_30443_, _30442_, _30438_);
  nor _80829_ (_30444_, _30443_, _08828_);
  nor _80830_ (_30445_, _12327_, _11072_);
  nor _80831_ (_30446_, _30445_, _07766_);
  and _80832_ (_30448_, _05284_, _04303_);
  nor _80833_ (_30449_, _30448_, _05886_);
  nor _80834_ (_30450_, _30449_, _30446_);
  nor _80835_ (_30451_, _30450_, _30415_);
  nor _80836_ (_30452_, _30451_, _30444_);
  nor _80837_ (_30453_, _30452_, _03780_);
  nor _80838_ (_30454_, _12333_, _11072_);
  nor _80839_ (_30455_, _30454_, _07778_);
  and _80840_ (_30456_, _30455_, _30439_);
  nor _80841_ (_30457_, _30456_, _30453_);
  nor _80842_ (_30459_, _30457_, _03622_);
  nor _80843_ (_30460_, _12207_, _11072_);
  nor _80844_ (_30461_, _30460_, _07777_);
  and _80845_ (_30462_, _30461_, _30439_);
  nor _80846_ (_30463_, _30462_, _30459_);
  nor _80847_ (_30464_, _30463_, _03790_);
  nor _80848_ (_30465_, _30406_, _05618_);
  nor _80849_ (_30466_, _30465_, _06828_);
  and _80850_ (_30467_, _30466_, _30417_);
  nor _80851_ (_30469_, _30467_, _30464_);
  or _80852_ (_30472_, _30469_, _18499_);
  and _80853_ (_30474_, _30416_, _05617_);
  nor _80854_ (_30476_, _30474_, _07793_);
  and _80855_ (_30478_, _30476_, _30439_);
  nor _80856_ (_30480_, _30478_, _03815_);
  and _80857_ (_30482_, _30448_, _05617_);
  or _80858_ (_30484_, _30415_, _07795_);
  or _80859_ (_30486_, _30484_, _30482_);
  and _80860_ (_30488_, _30486_, _30480_);
  and _80861_ (_30490_, _30488_, _30472_);
  nor _80862_ (_30492_, _30424_, _04246_);
  nor _80863_ (_30493_, _30492_, _30490_);
  and _80864_ (_30494_, _30493_, _03514_);
  nor _80865_ (_30495_, _30423_, _30406_);
  nor _80866_ (_30496_, _30495_, _03514_);
  or _80867_ (_30497_, _30496_, _30494_);
  or _80868_ (_30498_, _30497_, _43004_);
  or _80869_ (_30499_, _43000_, \oc8051_golden_model_1.TL0 [1]);
  and _80870_ (_30500_, _30499_, _41806_);
  and _80871_ (_43643_, _30500_, _30498_);
  not _80872_ (_30502_, \oc8051_golden_model_1.TL0 [2]);
  nor _80873_ (_30503_, _05284_, _30502_);
  nor _80874_ (_30504_, _12538_, _11072_);
  nor _80875_ (_30505_, _30504_, _30503_);
  nor _80876_ (_30506_, _30505_, _07793_);
  nor _80877_ (_30507_, _11072_, _04875_);
  nor _80878_ (_30508_, _30507_, _30503_);
  and _80879_ (_30509_, _30508_, _07390_);
  nor _80880_ (_30510_, _12416_, _11072_);
  nor _80881_ (_30511_, _30510_, _30503_);
  nor _80882_ (_30513_, _30511_, _04081_);
  nor _80883_ (_30514_, _04409_, _30502_);
  and _80884_ (_30515_, _05284_, \oc8051_golden_model_1.ACC [2]);
  nor _80885_ (_30516_, _30515_, _30503_);
  nor _80886_ (_30517_, _30516_, _09029_);
  nor _80887_ (_30518_, _30517_, _30514_);
  nor _80888_ (_30519_, _30518_, _03610_);
  or _80889_ (_30520_, _30519_, _30513_);
  and _80890_ (_30521_, _30520_, _03996_);
  nor _80891_ (_30522_, _30508_, _03996_);
  or _80892_ (_30524_, _30522_, _30521_);
  and _80893_ (_30525_, _30524_, _03737_);
  nor _80894_ (_30526_, _30516_, _03737_);
  nor _80895_ (_30527_, _30526_, _07390_);
  not _80896_ (_30528_, _30527_);
  nor _80897_ (_30529_, _30528_, _30525_);
  nor _80898_ (_30530_, _30529_, _30509_);
  nor _80899_ (_30531_, _30530_, _04481_);
  and _80900_ (_30532_, _06637_, _05284_);
  nor _80901_ (_30533_, _30503_, _07400_);
  not _80902_ (_30535_, _30533_);
  nor _80903_ (_30536_, _30535_, _30532_);
  nor _80904_ (_30537_, _30536_, _30531_);
  nor _80905_ (_30538_, _30537_, _03222_);
  nor _80906_ (_30539_, _12519_, _11072_);
  or _80907_ (_30540_, _30503_, _03589_);
  nor _80908_ (_30541_, _30540_, _30539_);
  or _80909_ (_30542_, _30541_, _03601_);
  nor _80910_ (_30543_, _30542_, _30538_);
  and _80911_ (_30544_, _05284_, _06332_);
  nor _80912_ (_30546_, _30544_, _30503_);
  nor _80913_ (_30547_, _30546_, _05886_);
  or _80914_ (_30548_, _30547_, _30543_);
  and _80915_ (_30549_, _30548_, _07766_);
  and _80916_ (_30550_, _12533_, _05284_);
  nor _80917_ (_30551_, _30550_, _30503_);
  nor _80918_ (_30552_, _30551_, _07766_);
  or _80919_ (_30553_, _30552_, _30549_);
  nor _80920_ (_30554_, _30553_, _03780_);
  and _80921_ (_30555_, _12539_, _05284_);
  or _80922_ (_30557_, _30503_, _07778_);
  nor _80923_ (_30558_, _30557_, _30555_);
  or _80924_ (_30559_, _30558_, _03622_);
  nor _80925_ (_30560_, _30559_, _30554_);
  nor _80926_ (_30561_, _30503_, _05718_);
  or _80927_ (_30562_, _30546_, _07777_);
  nor _80928_ (_30563_, _30562_, _30561_);
  nor _80929_ (_30564_, _30563_, _30560_);
  nor _80930_ (_30565_, _30564_, _03790_);
  or _80931_ (_30566_, _30561_, _06828_);
  or _80932_ (_30568_, _30566_, _30516_);
  and _80933_ (_30569_, _30568_, _07795_);
  not _80934_ (_30570_, _30569_);
  nor _80935_ (_30571_, _30570_, _30565_);
  nor _80936_ (_30572_, _12532_, _11072_);
  or _80937_ (_30573_, _30503_, _07795_);
  nor _80938_ (_30574_, _30573_, _30572_);
  or _80939_ (_30575_, _30574_, _03785_);
  nor _80940_ (_30576_, _30575_, _30571_);
  nor _80941_ (_30577_, _30576_, _30506_);
  nor _80942_ (_30579_, _30577_, _03815_);
  nor _80943_ (_30580_, _30511_, _04246_);
  or _80944_ (_30581_, _30580_, _03447_);
  nor _80945_ (_30582_, _30581_, _30579_);
  and _80946_ (_30583_, _12592_, _05284_);
  or _80947_ (_30584_, _30503_, _03514_);
  nor _80948_ (_30585_, _30584_, _30583_);
  nor _80949_ (_30586_, _30585_, _30582_);
  or _80950_ (_30587_, _30586_, _43004_);
  or _80951_ (_30588_, _43000_, \oc8051_golden_model_1.TL0 [2]);
  and _80952_ (_30590_, _30588_, _41806_);
  and _80953_ (_43644_, _30590_, _30587_);
  not _80954_ (_30591_, \oc8051_golden_model_1.TL0 [3]);
  nor _80955_ (_30592_, _05284_, _30591_);
  nor _80956_ (_30593_, _12738_, _11072_);
  nor _80957_ (_30594_, _30593_, _30592_);
  nor _80958_ (_30595_, _30594_, _07793_);
  and _80959_ (_30596_, _12739_, _05284_);
  nor _80960_ (_30597_, _30596_, _30592_);
  nor _80961_ (_30598_, _30597_, _07778_);
  and _80962_ (_30600_, _06592_, _05284_);
  or _80963_ (_30601_, _30600_, _30592_);
  and _80964_ (_30602_, _30601_, _04481_);
  and _80965_ (_30603_, _05284_, \oc8051_golden_model_1.ACC [3]);
  nor _80966_ (_30604_, _30603_, _30592_);
  nor _80967_ (_30605_, _30604_, _03737_);
  nor _80968_ (_30606_, _30604_, _09029_);
  nor _80969_ (_30607_, _04409_, _30591_);
  or _80970_ (_30608_, _30607_, _30606_);
  and _80971_ (_30609_, _30608_, _04081_);
  nor _80972_ (_30611_, _12627_, _11072_);
  nor _80973_ (_30612_, _30611_, _30592_);
  nor _80974_ (_30613_, _30612_, _04081_);
  or _80975_ (_30614_, _30613_, _30609_);
  and _80976_ (_30615_, _30614_, _03996_);
  nor _80977_ (_30616_, _11072_, _05005_);
  nor _80978_ (_30617_, _30616_, _30592_);
  nor _80979_ (_30618_, _30617_, _03996_);
  nor _80980_ (_30619_, _30618_, _30615_);
  nor _80981_ (_30620_, _30619_, _03729_);
  or _80982_ (_30622_, _30620_, _07390_);
  nor _80983_ (_30623_, _30622_, _30605_);
  and _80984_ (_30624_, _30617_, _07390_);
  or _80985_ (_30625_, _30624_, _04481_);
  nor _80986_ (_30626_, _30625_, _30623_);
  or _80987_ (_30627_, _30626_, _30602_);
  and _80988_ (_30628_, _30627_, _03589_);
  nor _80989_ (_30629_, _12718_, _11072_);
  nor _80990_ (_30630_, _30629_, _30592_);
  nor _80991_ (_30631_, _30630_, _03589_);
  or _80992_ (_30633_, _30631_, _08828_);
  or _80993_ (_30634_, _30633_, _30628_);
  and _80994_ (_30635_, _12733_, _05284_);
  or _80995_ (_30636_, _30592_, _07766_);
  or _80996_ (_30637_, _30636_, _30635_);
  and _80997_ (_30638_, _05284_, _06276_);
  nor _80998_ (_30639_, _30638_, _30592_);
  and _80999_ (_30640_, _30639_, _03601_);
  nor _81000_ (_30641_, _30640_, _03780_);
  and _81001_ (_30642_, _30641_, _30637_);
  and _81002_ (_30644_, _30642_, _30634_);
  nor _81003_ (_30645_, _30644_, _30598_);
  nor _81004_ (_30646_, _30645_, _03622_);
  nor _81005_ (_30647_, _30592_, _05567_);
  not _81006_ (_30648_, _30647_);
  nor _81007_ (_30649_, _30639_, _07777_);
  and _81008_ (_30650_, _30649_, _30648_);
  nor _81009_ (_30651_, _30650_, _30646_);
  nor _81010_ (_30652_, _30651_, _03790_);
  nor _81011_ (_30653_, _30604_, _06828_);
  and _81012_ (_30655_, _30653_, _30648_);
  or _81013_ (_30656_, _30655_, _30652_);
  and _81014_ (_30657_, _30656_, _07795_);
  nor _81015_ (_30658_, _12732_, _11072_);
  nor _81016_ (_30659_, _30658_, _30592_);
  nor _81017_ (_30660_, _30659_, _07795_);
  or _81018_ (_30661_, _30660_, _30657_);
  and _81019_ (_30662_, _30661_, _07793_);
  nor _81020_ (_30663_, _30662_, _30595_);
  nor _81021_ (_30664_, _30663_, _03815_);
  nor _81022_ (_30666_, _30612_, _04246_);
  or _81023_ (_30667_, _30666_, _03447_);
  nor _81024_ (_30668_, _30667_, _30664_);
  and _81025_ (_30669_, _12794_, _05284_);
  or _81026_ (_30670_, _30592_, _03514_);
  nor _81027_ (_30671_, _30670_, _30669_);
  nor _81028_ (_30672_, _30671_, _30668_);
  or _81029_ (_30673_, _30672_, _43004_);
  or _81030_ (_30674_, _43000_, \oc8051_golden_model_1.TL0 [3]);
  and _81031_ (_30675_, _30674_, _41806_);
  and _81032_ (_43645_, _30675_, _30673_);
  not _81033_ (_30677_, \oc8051_golden_model_1.TL0 [4]);
  nor _81034_ (_30678_, _05284_, _30677_);
  nor _81035_ (_30679_, _12816_, _11072_);
  nor _81036_ (_30680_, _30679_, _30678_);
  nor _81037_ (_30681_, _30680_, _07793_);
  and _81038_ (_30682_, _12817_, _05284_);
  nor _81039_ (_30683_, _30682_, _30678_);
  nor _81040_ (_30684_, _30683_, _07778_);
  and _81041_ (_30685_, _06298_, _05284_);
  nor _81042_ (_30687_, _30685_, _30678_);
  and _81043_ (_30688_, _30687_, _03601_);
  nor _81044_ (_30689_, _05777_, _11072_);
  nor _81045_ (_30690_, _30689_, _30678_);
  and _81046_ (_30691_, _30690_, _07390_);
  and _81047_ (_30692_, _05284_, \oc8051_golden_model_1.ACC [4]);
  nor _81048_ (_30693_, _30692_, _30678_);
  nor _81049_ (_30694_, _30693_, _03737_);
  nor _81050_ (_30695_, _30693_, _09029_);
  nor _81051_ (_30696_, _04409_, _30677_);
  or _81052_ (_30698_, _30696_, _30695_);
  and _81053_ (_30699_, _30698_, _04081_);
  nor _81054_ (_30700_, _12841_, _11072_);
  nor _81055_ (_30701_, _30700_, _30678_);
  nor _81056_ (_30702_, _30701_, _04081_);
  or _81057_ (_30703_, _30702_, _30699_);
  and _81058_ (_30704_, _30703_, _03996_);
  nor _81059_ (_30705_, _30690_, _03996_);
  nor _81060_ (_30706_, _30705_, _30704_);
  nor _81061_ (_30707_, _30706_, _03729_);
  or _81062_ (_30709_, _30707_, _07390_);
  nor _81063_ (_30710_, _30709_, _30694_);
  nor _81064_ (_30711_, _30710_, _30691_);
  nor _81065_ (_30712_, _30711_, _04481_);
  and _81066_ (_30713_, _06730_, _05284_);
  nor _81067_ (_30714_, _30678_, _07400_);
  not _81068_ (_30715_, _30714_);
  nor _81069_ (_30716_, _30715_, _30713_);
  or _81070_ (_30717_, _30716_, _03222_);
  nor _81071_ (_30718_, _30717_, _30712_);
  nor _81072_ (_30720_, _12933_, _11072_);
  nor _81073_ (_30721_, _30720_, _30678_);
  nor _81074_ (_30722_, _30721_, _03589_);
  or _81075_ (_30723_, _30722_, _03601_);
  nor _81076_ (_30724_, _30723_, _30718_);
  nor _81077_ (_30725_, _30724_, _30688_);
  or _81078_ (_30726_, _30725_, _03600_);
  and _81079_ (_30727_, _12821_, _05284_);
  or _81080_ (_30728_, _30727_, _30678_);
  or _81081_ (_30729_, _30728_, _07766_);
  and _81082_ (_30731_, _30729_, _07778_);
  and _81083_ (_30732_, _30731_, _30726_);
  nor _81084_ (_30733_, _30732_, _30684_);
  nor _81085_ (_30734_, _30733_, _03622_);
  nor _81086_ (_30735_, _30678_, _05825_);
  not _81087_ (_30736_, _30735_);
  nor _81088_ (_30737_, _30687_, _07777_);
  and _81089_ (_30738_, _30737_, _30736_);
  nor _81090_ (_30739_, _30738_, _30734_);
  nor _81091_ (_30740_, _30739_, _03790_);
  nor _81092_ (_30742_, _30693_, _06828_);
  and _81093_ (_30743_, _30742_, _30736_);
  or _81094_ (_30744_, _30743_, _30740_);
  and _81095_ (_30745_, _30744_, _07795_);
  nor _81096_ (_30746_, _12819_, _11072_);
  nor _81097_ (_30747_, _30746_, _30678_);
  nor _81098_ (_30748_, _30747_, _07795_);
  or _81099_ (_30749_, _30748_, _30745_);
  and _81100_ (_30750_, _30749_, _07793_);
  nor _81101_ (_30751_, _30750_, _30681_);
  nor _81102_ (_30753_, _30751_, _03815_);
  nor _81103_ (_30754_, _30701_, _04246_);
  or _81104_ (_30755_, _30754_, _03447_);
  nor _81105_ (_30756_, _30755_, _30753_);
  and _81106_ (_30757_, _13003_, _05284_);
  or _81107_ (_30758_, _30678_, _03514_);
  nor _81108_ (_30759_, _30758_, _30757_);
  nor _81109_ (_30760_, _30759_, _30756_);
  or _81110_ (_30761_, _30760_, _43004_);
  or _81111_ (_30762_, _43000_, \oc8051_golden_model_1.TL0 [4]);
  and _81112_ (_30764_, _30762_, _41806_);
  and _81113_ (_43646_, _30764_, _30761_);
  not _81114_ (_30765_, \oc8051_golden_model_1.TL0 [5]);
  nor _81115_ (_30766_, _05284_, _30765_);
  nor _81116_ (_30767_, _13146_, _11072_);
  nor _81117_ (_30768_, _30767_, _30766_);
  nor _81118_ (_30769_, _30768_, _07793_);
  and _81119_ (_30770_, _13147_, _05284_);
  nor _81120_ (_30771_, _30770_, _30766_);
  nor _81121_ (_30772_, _30771_, _07778_);
  and _81122_ (_30774_, _06684_, _05284_);
  or _81123_ (_30775_, _30774_, _30766_);
  and _81124_ (_30776_, _30775_, _04481_);
  and _81125_ (_30777_, _05284_, \oc8051_golden_model_1.ACC [5]);
  nor _81126_ (_30778_, _30777_, _30766_);
  nor _81127_ (_30779_, _30778_, _03737_);
  nor _81128_ (_30780_, _30778_, _09029_);
  nor _81129_ (_30781_, _04409_, _30765_);
  or _81130_ (_30782_, _30781_, _30780_);
  and _81131_ (_30783_, _30782_, _04081_);
  nor _81132_ (_30785_, _13014_, _11072_);
  nor _81133_ (_30786_, _30785_, _30766_);
  nor _81134_ (_30787_, _30786_, _04081_);
  or _81135_ (_30788_, _30787_, _30783_);
  and _81136_ (_30789_, _30788_, _03996_);
  nor _81137_ (_30790_, _05469_, _11072_);
  nor _81138_ (_30791_, _30790_, _30766_);
  nor _81139_ (_30792_, _30791_, _03996_);
  nor _81140_ (_30793_, _30792_, _30789_);
  nor _81141_ (_30794_, _30793_, _03729_);
  or _81142_ (_30796_, _30794_, _07390_);
  nor _81143_ (_30797_, _30796_, _30779_);
  and _81144_ (_30798_, _30791_, _07390_);
  or _81145_ (_30799_, _30798_, _04481_);
  nor _81146_ (_30800_, _30799_, _30797_);
  or _81147_ (_30801_, _30800_, _30776_);
  and _81148_ (_30802_, _30801_, _03589_);
  nor _81149_ (_30803_, _13127_, _11072_);
  nor _81150_ (_30804_, _30803_, _30766_);
  nor _81151_ (_30805_, _30804_, _03589_);
  or _81152_ (_30807_, _30805_, _08828_);
  or _81153_ (_30808_, _30807_, _30802_);
  and _81154_ (_30809_, _13141_, _05284_);
  or _81155_ (_30810_, _30766_, _07766_);
  or _81156_ (_30811_, _30810_, _30809_);
  and _81157_ (_30812_, _06306_, _05284_);
  nor _81158_ (_30813_, _30812_, _30766_);
  and _81159_ (_30814_, _30813_, _03601_);
  nor _81160_ (_30815_, _30814_, _03780_);
  and _81161_ (_30816_, _30815_, _30811_);
  and _81162_ (_30817_, _30816_, _30808_);
  nor _81163_ (_30818_, _30817_, _30772_);
  nor _81164_ (_30819_, _30818_, _03622_);
  nor _81165_ (_30820_, _30766_, _05518_);
  not _81166_ (_30821_, _30820_);
  nor _81167_ (_30822_, _30813_, _07777_);
  and _81168_ (_30823_, _30822_, _30821_);
  nor _81169_ (_30824_, _30823_, _30819_);
  nor _81170_ (_30825_, _30824_, _03790_);
  nor _81171_ (_30826_, _30778_, _06828_);
  and _81172_ (_30828_, _30826_, _30821_);
  nor _81173_ (_30829_, _30828_, _03624_);
  not _81174_ (_30830_, _30829_);
  nor _81175_ (_30831_, _30830_, _30825_);
  nor _81176_ (_30832_, _13140_, _11072_);
  or _81177_ (_30833_, _30766_, _07795_);
  nor _81178_ (_30834_, _30833_, _30832_);
  or _81179_ (_30835_, _30834_, _03785_);
  nor _81180_ (_30836_, _30835_, _30831_);
  nor _81181_ (_30837_, _30836_, _30769_);
  nor _81182_ (_30839_, _30837_, _03815_);
  nor _81183_ (_30840_, _30786_, _04246_);
  or _81184_ (_30841_, _30840_, _03447_);
  nor _81185_ (_30842_, _30841_, _30839_);
  and _81186_ (_30843_, _13199_, _05284_);
  or _81187_ (_30844_, _30766_, _03514_);
  nor _81188_ (_30845_, _30844_, _30843_);
  nor _81189_ (_30846_, _30845_, _30842_);
  or _81190_ (_30847_, _30846_, _43004_);
  or _81191_ (_30848_, _43000_, \oc8051_golden_model_1.TL0 [5]);
  and _81192_ (_30850_, _30848_, _41806_);
  and _81193_ (_43647_, _30850_, _30847_);
  not _81194_ (_30851_, \oc8051_golden_model_1.TL0 [6]);
  nor _81195_ (_30852_, _05284_, _30851_);
  nor _81196_ (_30853_, _13352_, _11072_);
  nor _81197_ (_30854_, _30853_, _30852_);
  nor _81198_ (_30855_, _30854_, _07793_);
  and _81199_ (_30856_, _13353_, _05284_);
  nor _81200_ (_30857_, _30856_, _30852_);
  nor _81201_ (_30858_, _30857_, _07778_);
  and _81202_ (_30860_, _06455_, _05284_);
  or _81203_ (_30861_, _30860_, _30852_);
  and _81204_ (_30862_, _30861_, _04481_);
  and _81205_ (_30863_, _05284_, \oc8051_golden_model_1.ACC [6]);
  nor _81206_ (_30864_, _30863_, _30852_);
  nor _81207_ (_30865_, _30864_, _03737_);
  nor _81208_ (_30866_, _30864_, _09029_);
  nor _81209_ (_30867_, _04409_, _30851_);
  or _81210_ (_30868_, _30867_, _30866_);
  and _81211_ (_30869_, _30868_, _04081_);
  nor _81212_ (_30871_, _13242_, _11072_);
  nor _81213_ (_30872_, _30871_, _30852_);
  nor _81214_ (_30873_, _30872_, _04081_);
  or _81215_ (_30874_, _30873_, _30869_);
  and _81216_ (_30875_, _30874_, _03996_);
  nor _81217_ (_30876_, _05363_, _11072_);
  nor _81218_ (_30877_, _30876_, _30852_);
  nor _81219_ (_30878_, _30877_, _03996_);
  nor _81220_ (_30879_, _30878_, _30875_);
  nor _81221_ (_30880_, _30879_, _03729_);
  or _81222_ (_30881_, _30880_, _07390_);
  nor _81223_ (_30882_, _30881_, _30865_);
  and _81224_ (_30883_, _30877_, _07390_);
  or _81225_ (_30884_, _30883_, _04481_);
  nor _81226_ (_30885_, _30884_, _30882_);
  or _81227_ (_30886_, _30885_, _30862_);
  and _81228_ (_30887_, _30886_, _03589_);
  nor _81229_ (_30888_, _13332_, _11072_);
  nor _81230_ (_30889_, _30888_, _30852_);
  nor _81231_ (_30890_, _30889_, _03589_);
  or _81232_ (_30893_, _30890_, _08828_);
  or _81233_ (_30894_, _30893_, _30887_);
  and _81234_ (_30895_, _13347_, _05284_);
  or _81235_ (_30896_, _30852_, _07766_);
  or _81236_ (_30897_, _30896_, _30895_);
  and _81237_ (_30898_, _13339_, _05284_);
  nor _81238_ (_30899_, _30898_, _30852_);
  and _81239_ (_30900_, _30899_, _03601_);
  nor _81240_ (_30901_, _30900_, _03780_);
  and _81241_ (_30902_, _30901_, _30897_);
  and _81242_ (_30904_, _30902_, _30894_);
  nor _81243_ (_30905_, _30904_, _30858_);
  nor _81244_ (_30906_, _30905_, _03622_);
  nor _81245_ (_30907_, _30852_, _05412_);
  not _81246_ (_30908_, _30907_);
  nor _81247_ (_30909_, _30899_, _07777_);
  and _81248_ (_30910_, _30909_, _30908_);
  nor _81249_ (_30911_, _30910_, _30906_);
  nor _81250_ (_30912_, _30911_, _03790_);
  nor _81251_ (_30913_, _30864_, _06828_);
  and _81252_ (_30915_, _30913_, _30908_);
  nor _81253_ (_30916_, _30915_, _03624_);
  not _81254_ (_30917_, _30916_);
  nor _81255_ (_30918_, _30917_, _30912_);
  nor _81256_ (_30919_, _13346_, _11072_);
  or _81257_ (_30920_, _30852_, _07795_);
  nor _81258_ (_30921_, _30920_, _30919_);
  or _81259_ (_30922_, _30921_, _03785_);
  nor _81260_ (_30923_, _30922_, _30918_);
  nor _81261_ (_30924_, _30923_, _30855_);
  nor _81262_ (_30926_, _30924_, _03815_);
  nor _81263_ (_30927_, _30872_, _04246_);
  or _81264_ (_30928_, _30927_, _03447_);
  nor _81265_ (_30929_, _30928_, _30926_);
  and _81266_ (_30930_, _13402_, _05284_);
  or _81267_ (_30931_, _30852_, _03514_);
  nor _81268_ (_30932_, _30931_, _30930_);
  nor _81269_ (_30933_, _30932_, _30929_);
  or _81270_ (_30934_, _30933_, _43004_);
  or _81271_ (_30935_, _43000_, \oc8051_golden_model_1.TL0 [6]);
  and _81272_ (_30937_, _30935_, _41806_);
  and _81273_ (_43648_, _30937_, _30934_);
  not _81274_ (_30938_, \oc8051_golden_model_1.TL1 [0]);
  nor _81275_ (_30939_, _05271_, _30938_);
  nor _81276_ (_30940_, _05666_, _11154_);
  nor _81277_ (_30941_, _30940_, _30939_);
  and _81278_ (_30942_, _30941_, _17166_);
  and _81279_ (_30943_, _05271_, \oc8051_golden_model_1.ACC [0]);
  nor _81280_ (_30944_, _30943_, _30939_);
  nor _81281_ (_30945_, _30944_, _03737_);
  nor _81282_ (_30947_, _30944_, _09029_);
  nor _81283_ (_30948_, _04409_, _30938_);
  or _81284_ (_30949_, _30948_, _30947_);
  and _81285_ (_30950_, _30949_, _04081_);
  nor _81286_ (_30951_, _30941_, _04081_);
  or _81287_ (_30952_, _30951_, _30950_);
  and _81288_ (_30953_, _30952_, _03996_);
  and _81289_ (_30954_, _05271_, _04620_);
  nor _81290_ (_30955_, _30954_, _30939_);
  nor _81291_ (_30956_, _30955_, _03996_);
  nor _81292_ (_30958_, _30956_, _30953_);
  nor _81293_ (_30959_, _30958_, _03729_);
  or _81294_ (_30960_, _30959_, _07390_);
  nor _81295_ (_30961_, _30960_, _30945_);
  and _81296_ (_30962_, _30955_, _07390_);
  nor _81297_ (_30963_, _30962_, _30961_);
  nor _81298_ (_30964_, _30963_, _04481_);
  and _81299_ (_30965_, _06546_, _05271_);
  nor _81300_ (_30966_, _30939_, _07400_);
  not _81301_ (_30967_, _30966_);
  nor _81302_ (_30969_, _30967_, _30965_);
  nor _81303_ (_30970_, _30969_, _30964_);
  nor _81304_ (_30971_, _30970_, _03222_);
  nor _81305_ (_30972_, _12109_, _11154_);
  or _81306_ (_30973_, _30939_, _03589_);
  nor _81307_ (_30974_, _30973_, _30972_);
  or _81308_ (_30975_, _30974_, _03601_);
  nor _81309_ (_30976_, _30975_, _30971_);
  and _81310_ (_30977_, _05271_, _06274_);
  nor _81311_ (_30978_, _30977_, _30939_);
  nor _81312_ (_30980_, _30978_, _05886_);
  or _81313_ (_30981_, _30980_, _30976_);
  and _81314_ (_30982_, _30981_, _07766_);
  and _81315_ (_30983_, _12124_, _05271_);
  nor _81316_ (_30984_, _30983_, _30939_);
  nor _81317_ (_30985_, _30984_, _07766_);
  or _81318_ (_30986_, _30985_, _30982_);
  nor _81319_ (_30987_, _30986_, _03780_);
  and _81320_ (_30988_, _12128_, _05271_);
  or _81321_ (_30989_, _30939_, _07778_);
  nor _81322_ (_30991_, _30989_, _30988_);
  or _81323_ (_30992_, _30991_, _03622_);
  nor _81324_ (_30993_, _30992_, _30987_);
  or _81325_ (_30994_, _30978_, _07777_);
  nor _81326_ (_30995_, _30994_, _30940_);
  nor _81327_ (_30996_, _30995_, _30993_);
  nor _81328_ (_30997_, _30996_, _03790_);
  nor _81329_ (_30998_, _30939_, _05666_);
  or _81330_ (_30999_, _30998_, _06828_);
  nor _81331_ (_31000_, _30999_, _30944_);
  or _81332_ (_31002_, _31000_, _30997_);
  and _81333_ (_31003_, _31002_, _07795_);
  nor _81334_ (_31004_, _12122_, _11154_);
  nor _81335_ (_31005_, _31004_, _30939_);
  nor _81336_ (_31006_, _31005_, _07795_);
  or _81337_ (_31007_, _31006_, _31003_);
  and _81338_ (_31008_, _31007_, _07793_);
  nor _81339_ (_31009_, _12003_, _11154_);
  nor _81340_ (_31010_, _31009_, _30939_);
  nor _81341_ (_31011_, _31010_, _07793_);
  nor _81342_ (_31013_, _31011_, _17166_);
  not _81343_ (_31014_, _31013_);
  nor _81344_ (_31015_, _31014_, _31008_);
  nor _81345_ (_31016_, _31015_, _30942_);
  or _81346_ (_31017_, _31016_, _43004_);
  or _81347_ (_31018_, _43000_, \oc8051_golden_model_1.TL1 [0]);
  and _81348_ (_31019_, _31018_, _41806_);
  and _81349_ (_43649_, _31019_, _31017_);
  and _81350_ (_31020_, _06501_, _05271_);
  not _81351_ (_31021_, \oc8051_golden_model_1.TL1 [1]);
  nor _81352_ (_31023_, _05271_, _31021_);
  nor _81353_ (_31024_, _31023_, _07400_);
  not _81354_ (_31025_, _31024_);
  nor _81355_ (_31026_, _31025_, _31020_);
  not _81356_ (_31027_, _31026_);
  nor _81357_ (_31028_, _05271_, \oc8051_golden_model_1.TL1 [1]);
  and _81358_ (_31029_, _05271_, _03274_);
  nor _81359_ (_31030_, _31029_, _31028_);
  and _81360_ (_31031_, _31030_, _03729_);
  and _81361_ (_31032_, _31030_, _04409_);
  nor _81362_ (_31034_, _04409_, _31021_);
  or _81363_ (_31035_, _31034_, _31032_);
  and _81364_ (_31036_, _31035_, _04081_);
  and _81365_ (_31037_, _12213_, _05271_);
  nor _81366_ (_31038_, _31037_, _31028_);
  and _81367_ (_31039_, _31038_, _03610_);
  or _81368_ (_31040_, _31039_, _31036_);
  and _81369_ (_31041_, _31040_, _03996_);
  and _81370_ (_31042_, _05271_, _06764_);
  nor _81371_ (_31043_, _31042_, _31023_);
  nor _81372_ (_31045_, _31043_, _03996_);
  nor _81373_ (_31046_, _31045_, _31041_);
  nor _81374_ (_31047_, _31046_, _03729_);
  or _81375_ (_31048_, _31047_, _07390_);
  nor _81376_ (_31049_, _31048_, _31031_);
  and _81377_ (_31050_, _31043_, _07390_);
  nor _81378_ (_31051_, _31050_, _31049_);
  nor _81379_ (_31052_, _31051_, _04481_);
  nor _81380_ (_31053_, _31052_, _03222_);
  and _81381_ (_31054_, _31053_, _31027_);
  not _81382_ (_31056_, _31028_);
  and _81383_ (_31057_, _12313_, _05271_);
  nor _81384_ (_31058_, _31057_, _03589_);
  and _81385_ (_31059_, _31058_, _31056_);
  nor _81386_ (_31060_, _31059_, _31054_);
  nor _81387_ (_31061_, _31060_, _08828_);
  nor _81388_ (_31062_, _12327_, _11154_);
  nor _81389_ (_31063_, _31062_, _07766_);
  and _81390_ (_31064_, _05271_, _04303_);
  nor _81391_ (_31065_, _31064_, _05886_);
  nor _81392_ (_31067_, _31065_, _31063_);
  nor _81393_ (_31068_, _31067_, _31028_);
  nor _81394_ (_31069_, _31068_, _31061_);
  nor _81395_ (_31070_, _31069_, _03780_);
  nor _81396_ (_31071_, _12333_, _11154_);
  nor _81397_ (_31072_, _31071_, _07778_);
  and _81398_ (_31073_, _31072_, _31056_);
  nor _81399_ (_31074_, _31073_, _31070_);
  nor _81400_ (_31075_, _31074_, _03622_);
  nor _81401_ (_31076_, _12207_, _11154_);
  nor _81402_ (_31078_, _31076_, _07777_);
  and _81403_ (_31079_, _31078_, _31056_);
  nor _81404_ (_31080_, _31079_, _31075_);
  nor _81405_ (_31081_, _31080_, _03790_);
  nor _81406_ (_31082_, _31023_, _05618_);
  nor _81407_ (_31083_, _31082_, _06828_);
  and _81408_ (_31084_, _31083_, _31030_);
  nor _81409_ (_31085_, _31084_, _31081_);
  or _81410_ (_31086_, _31085_, _18499_);
  and _81411_ (_31087_, _31064_, _05617_);
  nor _81412_ (_31089_, _31087_, _07795_);
  and _81413_ (_31090_, _31089_, _31056_);
  not _81414_ (_31091_, _31090_);
  nand _81415_ (_31092_, _31029_, _05617_);
  nor _81416_ (_31093_, _31028_, _07793_);
  and _81417_ (_31094_, _31093_, _31092_);
  nor _81418_ (_31095_, _31094_, _03815_);
  and _81419_ (_31096_, _31095_, _31091_);
  and _81420_ (_31097_, _31096_, _31086_);
  nor _81421_ (_31098_, _31038_, _04246_);
  nor _81422_ (_31100_, _31098_, _31097_);
  and _81423_ (_31101_, _31100_, _03514_);
  nor _81424_ (_31102_, _31037_, _31023_);
  nor _81425_ (_31103_, _31102_, _03514_);
  or _81426_ (_31104_, _31103_, _31101_);
  or _81427_ (_31105_, _31104_, _43004_);
  or _81428_ (_31106_, _43000_, \oc8051_golden_model_1.TL1 [1]);
  and _81429_ (_31107_, _31106_, _41806_);
  and _81430_ (_43650_, _31107_, _31105_);
  not _81431_ (_31108_, \oc8051_golden_model_1.TL1 [2]);
  nor _81432_ (_31109_, _05271_, _31108_);
  nor _81433_ (_31110_, _12538_, _11154_);
  nor _81434_ (_31111_, _31110_, _31109_);
  nor _81435_ (_31112_, _31111_, _07793_);
  and _81436_ (_31113_, _12539_, _05271_);
  nor _81437_ (_31114_, _31113_, _31109_);
  nor _81438_ (_31115_, _31114_, _07778_);
  and _81439_ (_31116_, _05271_, \oc8051_golden_model_1.ACC [2]);
  nor _81440_ (_31117_, _31116_, _31109_);
  nor _81441_ (_31118_, _31117_, _03737_);
  nor _81442_ (_31121_, _31117_, _09029_);
  nor _81443_ (_31122_, _04409_, _31108_);
  or _81444_ (_31123_, _31122_, _31121_);
  and _81445_ (_31124_, _31123_, _04081_);
  nor _81446_ (_31125_, _12416_, _11154_);
  nor _81447_ (_31126_, _31125_, _31109_);
  nor _81448_ (_31127_, _31126_, _04081_);
  or _81449_ (_31128_, _31127_, _31124_);
  and _81450_ (_31129_, _31128_, _03996_);
  nor _81451_ (_31130_, _11154_, _04875_);
  nor _81452_ (_31132_, _31130_, _31109_);
  nor _81453_ (_31133_, _31132_, _03996_);
  nor _81454_ (_31134_, _31133_, _31129_);
  nor _81455_ (_31135_, _31134_, _03729_);
  or _81456_ (_31136_, _31135_, _07390_);
  nor _81457_ (_31137_, _31136_, _31118_);
  and _81458_ (_31138_, _31132_, _07390_);
  nor _81459_ (_31139_, _31138_, _31137_);
  nor _81460_ (_31140_, _31139_, _04481_);
  and _81461_ (_31141_, _06637_, _05271_);
  nor _81462_ (_31143_, _31109_, _07400_);
  not _81463_ (_31144_, _31143_);
  nor _81464_ (_31145_, _31144_, _31141_);
  nor _81465_ (_31146_, _31145_, _03222_);
  not _81466_ (_31147_, _31146_);
  nor _81467_ (_31148_, _31147_, _31140_);
  nor _81468_ (_31149_, _12519_, _11154_);
  nor _81469_ (_31150_, _31149_, _31109_);
  nor _81470_ (_31151_, _31150_, _03589_);
  or _81471_ (_31152_, _31151_, _08828_);
  or _81472_ (_31154_, _31152_, _31148_);
  and _81473_ (_31155_, _12533_, _05271_);
  or _81474_ (_31156_, _31109_, _07766_);
  or _81475_ (_31157_, _31156_, _31155_);
  and _81476_ (_31158_, _05271_, _06332_);
  nor _81477_ (_31159_, _31158_, _31109_);
  and _81478_ (_31160_, _31159_, _03601_);
  nor _81479_ (_31161_, _31160_, _03780_);
  and _81480_ (_31162_, _31161_, _31157_);
  and _81481_ (_31163_, _31162_, _31154_);
  nor _81482_ (_31165_, _31163_, _31115_);
  nor _81483_ (_31166_, _31165_, _03622_);
  nor _81484_ (_31167_, _31109_, _05718_);
  not _81485_ (_31168_, _31167_);
  nor _81486_ (_31169_, _31159_, _07777_);
  and _81487_ (_31170_, _31169_, _31168_);
  nor _81488_ (_31171_, _31170_, _31166_);
  nor _81489_ (_31172_, _31171_, _03790_);
  nor _81490_ (_31173_, _31117_, _06828_);
  and _81491_ (_31174_, _31173_, _31168_);
  nor _81492_ (_31176_, _31174_, _03624_);
  not _81493_ (_31177_, _31176_);
  nor _81494_ (_31178_, _31177_, _31172_);
  nor _81495_ (_31179_, _12532_, _11154_);
  or _81496_ (_31180_, _31109_, _07795_);
  nor _81497_ (_31181_, _31180_, _31179_);
  or _81498_ (_31182_, _31181_, _03785_);
  nor _81499_ (_31183_, _31182_, _31178_);
  nor _81500_ (_31184_, _31183_, _31112_);
  nor _81501_ (_31185_, _31184_, _03815_);
  nor _81502_ (_31187_, _31126_, _04246_);
  or _81503_ (_31188_, _31187_, _03447_);
  nor _81504_ (_31189_, _31188_, _31185_);
  and _81505_ (_31190_, _12592_, _05271_);
  or _81506_ (_31191_, _31109_, _03514_);
  nor _81507_ (_31192_, _31191_, _31190_);
  nor _81508_ (_31193_, _31192_, _31189_);
  or _81509_ (_31194_, _31193_, _43004_);
  or _81510_ (_31195_, _43000_, \oc8051_golden_model_1.TL1 [2]);
  and _81511_ (_31196_, _31195_, _41806_);
  and _81512_ (_43651_, _31196_, _31194_);
  not _81513_ (_31198_, \oc8051_golden_model_1.TL1 [3]);
  nor _81514_ (_31199_, _05271_, _31198_);
  nor _81515_ (_31200_, _12738_, _11154_);
  nor _81516_ (_31201_, _31200_, _31199_);
  nor _81517_ (_31202_, _31201_, _07793_);
  and _81518_ (_31203_, _12739_, _05271_);
  nor _81519_ (_31204_, _31203_, _31199_);
  nor _81520_ (_31205_, _31204_, _07778_);
  and _81521_ (_31206_, _06592_, _05271_);
  or _81522_ (_31208_, _31206_, _31199_);
  and _81523_ (_31209_, _31208_, _04481_);
  and _81524_ (_31210_, _05271_, \oc8051_golden_model_1.ACC [3]);
  nor _81525_ (_31211_, _31210_, _31199_);
  nor _81526_ (_31212_, _31211_, _03737_);
  nor _81527_ (_31213_, _31211_, _09029_);
  nor _81528_ (_31214_, _04409_, _31198_);
  or _81529_ (_31215_, _31214_, _31213_);
  and _81530_ (_31216_, _31215_, _04081_);
  nor _81531_ (_31217_, _12627_, _11154_);
  nor _81532_ (_31219_, _31217_, _31199_);
  nor _81533_ (_31220_, _31219_, _04081_);
  or _81534_ (_31221_, _31220_, _31216_);
  and _81535_ (_31222_, _31221_, _03996_);
  nor _81536_ (_31223_, _11154_, _05005_);
  nor _81537_ (_31224_, _31223_, _31199_);
  nor _81538_ (_31225_, _31224_, _03996_);
  nor _81539_ (_31226_, _31225_, _31222_);
  nor _81540_ (_31227_, _31226_, _03729_);
  or _81541_ (_31228_, _31227_, _07390_);
  nor _81542_ (_31230_, _31228_, _31212_);
  and _81543_ (_31231_, _31224_, _07390_);
  or _81544_ (_31232_, _31231_, _04481_);
  nor _81545_ (_31233_, _31232_, _31230_);
  or _81546_ (_31234_, _31233_, _31209_);
  and _81547_ (_31235_, _31234_, _03589_);
  nor _81548_ (_31236_, _12718_, _11154_);
  nor _81549_ (_31237_, _31236_, _31199_);
  nor _81550_ (_31238_, _31237_, _03589_);
  or _81551_ (_31239_, _31238_, _08828_);
  or _81552_ (_31241_, _31239_, _31235_);
  and _81553_ (_31242_, _12733_, _05271_);
  or _81554_ (_31243_, _31199_, _07766_);
  or _81555_ (_31244_, _31243_, _31242_);
  and _81556_ (_31245_, _05271_, _06276_);
  nor _81557_ (_31246_, _31245_, _31199_);
  and _81558_ (_31247_, _31246_, _03601_);
  nor _81559_ (_31248_, _31247_, _03780_);
  and _81560_ (_31249_, _31248_, _31244_);
  and _81561_ (_31250_, _31249_, _31241_);
  nor _81562_ (_31252_, _31250_, _31205_);
  nor _81563_ (_31253_, _31252_, _03622_);
  nor _81564_ (_31254_, _31199_, _05567_);
  not _81565_ (_31255_, _31254_);
  nor _81566_ (_31256_, _31246_, _07777_);
  and _81567_ (_31257_, _31256_, _31255_);
  nor _81568_ (_31258_, _31257_, _31253_);
  nor _81569_ (_31259_, _31258_, _03790_);
  nor _81570_ (_31260_, _31211_, _06828_);
  and _81571_ (_31261_, _31260_, _31255_);
  nor _81572_ (_31263_, _31261_, _03624_);
  not _81573_ (_31264_, _31263_);
  nor _81574_ (_31265_, _31264_, _31259_);
  nor _81575_ (_31266_, _12732_, _11154_);
  or _81576_ (_31267_, _31199_, _07795_);
  nor _81577_ (_31268_, _31267_, _31266_);
  or _81578_ (_31269_, _31268_, _03785_);
  nor _81579_ (_31270_, _31269_, _31265_);
  nor _81580_ (_31271_, _31270_, _31202_);
  nor _81581_ (_31272_, _31271_, _03815_);
  nor _81582_ (_31274_, _31219_, _04246_);
  or _81583_ (_31275_, _31274_, _03447_);
  nor _81584_ (_31276_, _31275_, _31272_);
  and _81585_ (_31277_, _12794_, _05271_);
  or _81586_ (_31278_, _31199_, _03514_);
  nor _81587_ (_31279_, _31278_, _31277_);
  nor _81588_ (_31280_, _31279_, _31276_);
  or _81589_ (_31281_, _31280_, _43004_);
  or _81590_ (_31282_, _43000_, \oc8051_golden_model_1.TL1 [3]);
  and _81591_ (_31283_, _31282_, _41806_);
  and _81592_ (_43652_, _31283_, _31281_);
  not _81593_ (_31285_, \oc8051_golden_model_1.TL1 [4]);
  nor _81594_ (_31286_, _05271_, _31285_);
  nor _81595_ (_31287_, _12816_, _11154_);
  nor _81596_ (_31288_, _31287_, _31286_);
  nor _81597_ (_31289_, _31288_, _07793_);
  and _81598_ (_31290_, _12817_, _05271_);
  nor _81599_ (_31291_, _31290_, _31286_);
  nor _81600_ (_31292_, _31291_, _07778_);
  and _81601_ (_31293_, _06298_, _05271_);
  nor _81602_ (_31295_, _31293_, _31286_);
  and _81603_ (_31296_, _31295_, _03601_);
  nor _81604_ (_31297_, _05777_, _11154_);
  nor _81605_ (_31298_, _31297_, _31286_);
  and _81606_ (_31299_, _31298_, _07390_);
  and _81607_ (_31300_, _05271_, \oc8051_golden_model_1.ACC [4]);
  nor _81608_ (_31301_, _31300_, _31286_);
  nor _81609_ (_31302_, _31301_, _03737_);
  nor _81610_ (_31303_, _31301_, _09029_);
  nor _81611_ (_31304_, _04409_, _31285_);
  or _81612_ (_31306_, _31304_, _31303_);
  and _81613_ (_31307_, _31306_, _04081_);
  nor _81614_ (_31308_, _12841_, _11154_);
  nor _81615_ (_31309_, _31308_, _31286_);
  nor _81616_ (_31310_, _31309_, _04081_);
  or _81617_ (_31311_, _31310_, _31307_);
  and _81618_ (_31312_, _31311_, _03996_);
  nor _81619_ (_31313_, _31298_, _03996_);
  nor _81620_ (_31314_, _31313_, _31312_);
  nor _81621_ (_31315_, _31314_, _03729_);
  or _81622_ (_31317_, _31315_, _07390_);
  nor _81623_ (_31318_, _31317_, _31302_);
  nor _81624_ (_31319_, _31318_, _31299_);
  nor _81625_ (_31320_, _31319_, _04481_);
  and _81626_ (_31321_, _06730_, _05271_);
  nor _81627_ (_31322_, _31286_, _07400_);
  not _81628_ (_31323_, _31322_);
  nor _81629_ (_31324_, _31323_, _31321_);
  or _81630_ (_31325_, _31324_, _03222_);
  nor _81631_ (_31326_, _31325_, _31320_);
  nor _81632_ (_31328_, _12933_, _11154_);
  nor _81633_ (_31329_, _31328_, _31286_);
  nor _81634_ (_31330_, _31329_, _03589_);
  or _81635_ (_31331_, _31330_, _03601_);
  nor _81636_ (_31332_, _31331_, _31326_);
  nor _81637_ (_31333_, _31332_, _31296_);
  or _81638_ (_31334_, _31333_, _03600_);
  and _81639_ (_31335_, _12821_, _05271_);
  or _81640_ (_31336_, _31335_, _31286_);
  or _81641_ (_31337_, _31336_, _07766_);
  and _81642_ (_31339_, _31337_, _07778_);
  and _81643_ (_31340_, _31339_, _31334_);
  nor _81644_ (_31341_, _31340_, _31292_);
  nor _81645_ (_31342_, _31341_, _03622_);
  nor _81646_ (_31343_, _31286_, _05825_);
  not _81647_ (_31344_, _31343_);
  nor _81648_ (_31345_, _31295_, _07777_);
  and _81649_ (_31346_, _31345_, _31344_);
  nor _81650_ (_31347_, _31346_, _31342_);
  nor _81651_ (_31348_, _31347_, _03790_);
  nor _81652_ (_31350_, _31301_, _06828_);
  and _81653_ (_31351_, _31350_, _31344_);
  nor _81654_ (_31352_, _31351_, _03624_);
  not _81655_ (_31353_, _31352_);
  nor _81656_ (_31354_, _31353_, _31348_);
  nor _81657_ (_31355_, _12819_, _11154_);
  or _81658_ (_31356_, _31286_, _07795_);
  nor _81659_ (_31357_, _31356_, _31355_);
  or _81660_ (_31358_, _31357_, _03785_);
  nor _81661_ (_31359_, _31358_, _31354_);
  nor _81662_ (_31361_, _31359_, _31289_);
  nor _81663_ (_31362_, _31361_, _03815_);
  nor _81664_ (_31363_, _31309_, _04246_);
  or _81665_ (_31364_, _31363_, _03447_);
  nor _81666_ (_31365_, _31364_, _31362_);
  and _81667_ (_31366_, _13003_, _05271_);
  or _81668_ (_31367_, _31286_, _03514_);
  nor _81669_ (_31368_, _31367_, _31366_);
  nor _81670_ (_31369_, _31368_, _31365_);
  or _81671_ (_31370_, _31369_, _43004_);
  or _81672_ (_31372_, _43000_, \oc8051_golden_model_1.TL1 [4]);
  and _81673_ (_31373_, _31372_, _41806_);
  and _81674_ (_43653_, _31373_, _31370_);
  not _81675_ (_31374_, \oc8051_golden_model_1.TL1 [5]);
  nor _81676_ (_31375_, _05271_, _31374_);
  nor _81677_ (_31376_, _13146_, _11154_);
  nor _81678_ (_31377_, _31376_, _31375_);
  nor _81679_ (_31378_, _31377_, _07793_);
  and _81680_ (_31379_, _13147_, _05271_);
  nor _81681_ (_31380_, _31379_, _31375_);
  nor _81682_ (_31382_, _31380_, _07778_);
  and _81683_ (_31383_, _06684_, _05271_);
  or _81684_ (_31384_, _31383_, _31375_);
  and _81685_ (_31385_, _31384_, _04481_);
  and _81686_ (_31386_, _05271_, \oc8051_golden_model_1.ACC [5]);
  nor _81687_ (_31387_, _31386_, _31375_);
  nor _81688_ (_31388_, _31387_, _03737_);
  nor _81689_ (_31389_, _31387_, _09029_);
  nor _81690_ (_31390_, _04409_, _31374_);
  or _81691_ (_31391_, _31390_, _31389_);
  and _81692_ (_31393_, _31391_, _04081_);
  nor _81693_ (_31394_, _13014_, _11154_);
  nor _81694_ (_31395_, _31394_, _31375_);
  nor _81695_ (_31396_, _31395_, _04081_);
  or _81696_ (_31397_, _31396_, _31393_);
  and _81697_ (_31398_, _31397_, _03996_);
  nor _81698_ (_31399_, _05469_, _11154_);
  nor _81699_ (_31400_, _31399_, _31375_);
  nor _81700_ (_31401_, _31400_, _03996_);
  nor _81701_ (_31402_, _31401_, _31398_);
  nor _81702_ (_31404_, _31402_, _03729_);
  or _81703_ (_31405_, _31404_, _07390_);
  nor _81704_ (_31406_, _31405_, _31388_);
  and _81705_ (_31407_, _31400_, _07390_);
  or _81706_ (_31408_, _31407_, _04481_);
  nor _81707_ (_31409_, _31408_, _31406_);
  or _81708_ (_31410_, _31409_, _31385_);
  and _81709_ (_31411_, _31410_, _03589_);
  nor _81710_ (_31412_, _13127_, _11154_);
  nor _81711_ (_31413_, _31412_, _31375_);
  nor _81712_ (_31415_, _31413_, _03589_);
  or _81713_ (_31416_, _31415_, _08828_);
  or _81714_ (_31417_, _31416_, _31411_);
  and _81715_ (_31418_, _13141_, _05271_);
  or _81716_ (_31419_, _31375_, _07766_);
  or _81717_ (_31420_, _31419_, _31418_);
  and _81718_ (_31421_, _06306_, _05271_);
  nor _81719_ (_31422_, _31421_, _31375_);
  and _81720_ (_31423_, _31422_, _03601_);
  nor _81721_ (_31424_, _31423_, _03780_);
  and _81722_ (_31426_, _31424_, _31420_);
  and _81723_ (_31427_, _31426_, _31417_);
  nor _81724_ (_31428_, _31427_, _31382_);
  nor _81725_ (_31429_, _31428_, _03622_);
  nor _81726_ (_31430_, _31375_, _05518_);
  not _81727_ (_31431_, _31430_);
  nor _81728_ (_31432_, _31422_, _07777_);
  and _81729_ (_31433_, _31432_, _31431_);
  nor _81730_ (_31434_, _31433_, _31429_);
  nor _81731_ (_31435_, _31434_, _03790_);
  nor _81732_ (_31437_, _31387_, _06828_);
  and _81733_ (_31438_, _31437_, _31431_);
  nor _81734_ (_31439_, _31438_, _03624_);
  not _81735_ (_31440_, _31439_);
  nor _81736_ (_31441_, _31440_, _31435_);
  nor _81737_ (_31442_, _13140_, _11154_);
  or _81738_ (_31443_, _31375_, _07795_);
  nor _81739_ (_31444_, _31443_, _31442_);
  or _81740_ (_31445_, _31444_, _03785_);
  nor _81741_ (_31446_, _31445_, _31441_);
  nor _81742_ (_31448_, _31446_, _31378_);
  nor _81743_ (_31449_, _31448_, _03815_);
  nor _81744_ (_31450_, _31395_, _04246_);
  or _81745_ (_31451_, _31450_, _03447_);
  nor _81746_ (_31452_, _31451_, _31449_);
  and _81747_ (_31453_, _13199_, _05271_);
  or _81748_ (_31454_, _31375_, _03514_);
  nor _81749_ (_31455_, _31454_, _31453_);
  nor _81750_ (_31456_, _31455_, _31452_);
  or _81751_ (_31457_, _31456_, _43004_);
  or _81752_ (_31459_, _43000_, \oc8051_golden_model_1.TL1 [5]);
  and _81753_ (_31460_, _31459_, _41806_);
  and _81754_ (_43654_, _31460_, _31457_);
  not _81755_ (_31461_, \oc8051_golden_model_1.TL1 [6]);
  nor _81756_ (_31462_, _05271_, _31461_);
  nor _81757_ (_31463_, _13352_, _11154_);
  nor _81758_ (_31464_, _31463_, _31462_);
  nor _81759_ (_31465_, _31464_, _07793_);
  and _81760_ (_31466_, _13353_, _05271_);
  nor _81761_ (_31467_, _31466_, _31462_);
  nor _81762_ (_31469_, _31467_, _07778_);
  and _81763_ (_31470_, _06455_, _05271_);
  or _81764_ (_31471_, _31470_, _31462_);
  and _81765_ (_31472_, _31471_, _04481_);
  and _81766_ (_31473_, _05271_, \oc8051_golden_model_1.ACC [6]);
  nor _81767_ (_31474_, _31473_, _31462_);
  nor _81768_ (_31475_, _31474_, _03737_);
  nor _81769_ (_31476_, _31474_, _09029_);
  nor _81770_ (_31477_, _04409_, _31461_);
  or _81771_ (_31478_, _31477_, _31476_);
  and _81772_ (_31480_, _31478_, _04081_);
  nor _81773_ (_31481_, _13242_, _11154_);
  nor _81774_ (_31482_, _31481_, _31462_);
  nor _81775_ (_31483_, _31482_, _04081_);
  or _81776_ (_31484_, _31483_, _31480_);
  and _81777_ (_31485_, _31484_, _03996_);
  nor _81778_ (_31486_, _05363_, _11154_);
  nor _81779_ (_31487_, _31486_, _31462_);
  nor _81780_ (_31488_, _31487_, _03996_);
  nor _81781_ (_31489_, _31488_, _31485_);
  nor _81782_ (_31491_, _31489_, _03729_);
  or _81783_ (_31492_, _31491_, _07390_);
  nor _81784_ (_31493_, _31492_, _31475_);
  and _81785_ (_31494_, _31487_, _07390_);
  or _81786_ (_31495_, _31494_, _04481_);
  nor _81787_ (_31496_, _31495_, _31493_);
  or _81788_ (_31497_, _31496_, _31472_);
  and _81789_ (_31498_, _31497_, _03589_);
  nor _81790_ (_31499_, _13332_, _11154_);
  nor _81791_ (_31500_, _31499_, _31462_);
  nor _81792_ (_31502_, _31500_, _03589_);
  or _81793_ (_31503_, _31502_, _08828_);
  or _81794_ (_31504_, _31503_, _31498_);
  and _81795_ (_31505_, _13347_, _05271_);
  or _81796_ (_31506_, _31462_, _07766_);
  or _81797_ (_31507_, _31506_, _31505_);
  and _81798_ (_31508_, _13339_, _05271_);
  nor _81799_ (_31509_, _31508_, _31462_);
  and _81800_ (_31510_, _31509_, _03601_);
  nor _81801_ (_31511_, _31510_, _03780_);
  and _81802_ (_31513_, _31511_, _31507_);
  and _81803_ (_31514_, _31513_, _31504_);
  nor _81804_ (_31515_, _31514_, _31469_);
  nor _81805_ (_31516_, _31515_, _03622_);
  nor _81806_ (_31517_, _31462_, _05412_);
  not _81807_ (_31518_, _31517_);
  nor _81808_ (_31519_, _31509_, _07777_);
  and _81809_ (_31520_, _31519_, _31518_);
  nor _81810_ (_31521_, _31520_, _31516_);
  nor _81811_ (_31522_, _31521_, _03790_);
  nor _81812_ (_31524_, _31474_, _06828_);
  and _81813_ (_31525_, _31524_, _31518_);
  or _81814_ (_31526_, _31525_, _31522_);
  and _81815_ (_31527_, _31526_, _07795_);
  nor _81816_ (_31528_, _13346_, _11154_);
  nor _81817_ (_31529_, _31528_, _31462_);
  nor _81818_ (_31530_, _31529_, _07795_);
  or _81819_ (_31531_, _31530_, _31527_);
  and _81820_ (_31532_, _31531_, _07793_);
  nor _81821_ (_31533_, _31532_, _31465_);
  nor _81822_ (_31535_, _31533_, _03815_);
  nor _81823_ (_31536_, _31482_, _04246_);
  or _81824_ (_31537_, _31536_, _03447_);
  nor _81825_ (_31538_, _31537_, _31535_);
  and _81826_ (_31539_, _13402_, _05271_);
  or _81827_ (_31540_, _31462_, _03514_);
  nor _81828_ (_31541_, _31540_, _31539_);
  nor _81829_ (_31542_, _31541_, _31538_);
  or _81830_ (_31543_, _31542_, _43004_);
  or _81831_ (_31544_, _43000_, \oc8051_golden_model_1.TL1 [6]);
  and _81832_ (_31546_, _31544_, _41806_);
  and _81833_ (_43655_, _31546_, _31543_);
  not _81834_ (_31547_, \oc8051_golden_model_1.TMOD [0]);
  nor _81835_ (_31548_, _05286_, _31547_);
  nor _81836_ (_31549_, _05666_, _11236_);
  nor _81837_ (_31550_, _31549_, _31548_);
  and _81838_ (_31551_, _31550_, _17166_);
  and _81839_ (_31552_, _05286_, \oc8051_golden_model_1.ACC [0]);
  nor _81840_ (_31553_, _31552_, _31548_);
  nor _81841_ (_31554_, _31553_, _03737_);
  nor _81842_ (_31555_, _31553_, _09029_);
  nor _81843_ (_31556_, _04409_, _31547_);
  or _81844_ (_31557_, _31556_, _31555_);
  and _81845_ (_31558_, _31557_, _04081_);
  nor _81846_ (_31559_, _31550_, _04081_);
  or _81847_ (_31560_, _31559_, _31558_);
  and _81848_ (_31561_, _31560_, _03996_);
  and _81849_ (_31562_, _05286_, _04620_);
  nor _81850_ (_31563_, _31562_, _31548_);
  nor _81851_ (_31564_, _31563_, _03996_);
  nor _81852_ (_31566_, _31564_, _31561_);
  nor _81853_ (_31567_, _31566_, _03729_);
  or _81854_ (_31568_, _31567_, _07390_);
  nor _81855_ (_31569_, _31568_, _31554_);
  and _81856_ (_31570_, _31563_, _07390_);
  nor _81857_ (_31571_, _31570_, _31569_);
  nor _81858_ (_31572_, _31571_, _04481_);
  and _81859_ (_31573_, _06546_, _05286_);
  nor _81860_ (_31574_, _31548_, _07400_);
  not _81861_ (_31575_, _31574_);
  nor _81862_ (_31577_, _31575_, _31573_);
  nor _81863_ (_31578_, _31577_, _31572_);
  nor _81864_ (_31579_, _31578_, _03222_);
  nor _81865_ (_31580_, _12109_, _11236_);
  or _81866_ (_31581_, _31548_, _03589_);
  nor _81867_ (_31582_, _31581_, _31580_);
  or _81868_ (_31583_, _31582_, _03601_);
  nor _81869_ (_31584_, _31583_, _31579_);
  and _81870_ (_31585_, _05286_, _06274_);
  nor _81871_ (_31586_, _31585_, _31548_);
  nor _81872_ (_31588_, _31586_, _05886_);
  or _81873_ (_31589_, _31588_, _31584_);
  and _81874_ (_31590_, _31589_, _07766_);
  and _81875_ (_31591_, _12124_, _05286_);
  nor _81876_ (_31592_, _31591_, _31548_);
  nor _81877_ (_31593_, _31592_, _07766_);
  or _81878_ (_31594_, _31593_, _31590_);
  nor _81879_ (_31595_, _31594_, _03780_);
  and _81880_ (_31596_, _12128_, _05286_);
  or _81881_ (_31597_, _31548_, _07778_);
  nor _81882_ (_31599_, _31597_, _31596_);
  or _81883_ (_31600_, _31599_, _03622_);
  nor _81884_ (_31601_, _31600_, _31595_);
  or _81885_ (_31602_, _31586_, _07777_);
  nor _81886_ (_31603_, _31602_, _31549_);
  nor _81887_ (_31604_, _31603_, _31601_);
  nor _81888_ (_31605_, _31604_, _03790_);
  and _81889_ (_31606_, _12005_, _05286_);
  or _81890_ (_31607_, _31606_, _31548_);
  and _81891_ (_31608_, _31607_, _03790_);
  or _81892_ (_31610_, _31608_, _31605_);
  and _81893_ (_31611_, _31610_, _07795_);
  nor _81894_ (_31612_, _12122_, _11236_);
  nor _81895_ (_31613_, _31612_, _31548_);
  nor _81896_ (_31614_, _31613_, _07795_);
  or _81897_ (_31615_, _31614_, _31611_);
  and _81898_ (_31616_, _31615_, _07793_);
  nor _81899_ (_31617_, _12003_, _11236_);
  nor _81900_ (_31618_, _31617_, _31548_);
  nor _81901_ (_31619_, _31618_, _07793_);
  nor _81902_ (_31621_, _31619_, _17166_);
  not _81903_ (_31622_, _31621_);
  nor _81904_ (_31623_, _31622_, _31616_);
  nor _81905_ (_31624_, _31623_, _31551_);
  or _81906_ (_31625_, _31624_, _43004_);
  or _81907_ (_31626_, _43000_, \oc8051_golden_model_1.TMOD [0]);
  and _81908_ (_31627_, _31626_, _41806_);
  and _81909_ (_43658_, _31627_, _31625_);
  and _81910_ (_31628_, _06501_, _05286_);
  not _81911_ (_31629_, \oc8051_golden_model_1.TMOD [1]);
  nor _81912_ (_31631_, _05286_, _31629_);
  nor _81913_ (_31632_, _31631_, _07400_);
  not _81914_ (_31633_, _31632_);
  nor _81915_ (_31634_, _31633_, _31628_);
  not _81916_ (_31635_, _31634_);
  and _81917_ (_31636_, _05286_, _06764_);
  nor _81918_ (_31637_, _31636_, _31631_);
  and _81919_ (_31638_, _31637_, _07390_);
  nor _81920_ (_31639_, _05286_, \oc8051_golden_model_1.TMOD [1]);
  and _81921_ (_31640_, _05286_, _03274_);
  nor _81922_ (_31642_, _31640_, _31639_);
  and _81923_ (_31643_, _31642_, _03729_);
  and _81924_ (_31644_, _31642_, _04409_);
  nor _81925_ (_31645_, _04409_, _31629_);
  or _81926_ (_31646_, _31645_, _31644_);
  and _81927_ (_31647_, _31646_, _04081_);
  and _81928_ (_31648_, _12213_, _05286_);
  nor _81929_ (_31649_, _31648_, _31639_);
  and _81930_ (_31650_, _31649_, _03610_);
  or _81931_ (_31651_, _31650_, _31647_);
  and _81932_ (_31653_, _31651_, _03996_);
  nor _81933_ (_31654_, _31637_, _03996_);
  nor _81934_ (_31655_, _31654_, _31653_);
  nor _81935_ (_31656_, _31655_, _03729_);
  or _81936_ (_31657_, _31656_, _07390_);
  nor _81937_ (_31658_, _31657_, _31643_);
  nor _81938_ (_31659_, _31658_, _31638_);
  nor _81939_ (_31660_, _31659_, _04481_);
  nor _81940_ (_31661_, _31660_, _03222_);
  and _81941_ (_31662_, _31661_, _31635_);
  not _81942_ (_31664_, _31639_);
  and _81943_ (_31665_, _12313_, _05286_);
  nor _81944_ (_31666_, _31665_, _03589_);
  and _81945_ (_31667_, _31666_, _31664_);
  nor _81946_ (_31668_, _31667_, _31662_);
  nor _81947_ (_31669_, _31668_, _08828_);
  nor _81948_ (_31670_, _12327_, _11236_);
  nor _81949_ (_31671_, _31670_, _07766_);
  and _81950_ (_31672_, _05286_, _04303_);
  nor _81951_ (_31673_, _31672_, _05886_);
  nor _81952_ (_31675_, _31673_, _31671_);
  nor _81953_ (_31676_, _31675_, _31639_);
  nor _81954_ (_31677_, _31676_, _31669_);
  nor _81955_ (_31678_, _31677_, _03780_);
  nor _81956_ (_31679_, _12333_, _11236_);
  nor _81957_ (_31680_, _31679_, _07778_);
  and _81958_ (_31681_, _31680_, _31664_);
  nor _81959_ (_31682_, _31681_, _31678_);
  nor _81960_ (_31683_, _31682_, _03622_);
  nor _81961_ (_31684_, _12207_, _11236_);
  nor _81962_ (_31685_, _31684_, _07777_);
  and _81963_ (_31686_, _31685_, _31664_);
  nor _81964_ (_31687_, _31686_, _31683_);
  nor _81965_ (_31688_, _31687_, _03790_);
  nor _81966_ (_31689_, _31631_, _05618_);
  nor _81967_ (_31690_, _31689_, _06828_);
  and _81968_ (_31691_, _31690_, _31642_);
  nor _81969_ (_31692_, _31691_, _31688_);
  or _81970_ (_31693_, _31692_, _18499_);
  and _81971_ (_31694_, _31672_, _05617_);
  nor _81972_ (_31697_, _31694_, _07795_);
  and _81973_ (_31698_, _31697_, _31664_);
  nand _81974_ (_31699_, _31640_, _05617_);
  nor _81975_ (_31700_, _31639_, _07793_);
  and _81976_ (_31701_, _31700_, _31699_);
  or _81977_ (_31702_, _31701_, _03815_);
  nor _81978_ (_31703_, _31702_, _31698_);
  and _81979_ (_31704_, _31703_, _31693_);
  nor _81980_ (_31705_, _31649_, _04246_);
  nor _81981_ (_31706_, _31705_, _31704_);
  and _81982_ (_31708_, _31706_, _03514_);
  nor _81983_ (_31709_, _31648_, _31631_);
  nor _81984_ (_31710_, _31709_, _03514_);
  or _81985_ (_31711_, _31710_, _31708_);
  or _81986_ (_31712_, _31711_, _43004_);
  or _81987_ (_31713_, _43000_, \oc8051_golden_model_1.TMOD [1]);
  and _81988_ (_31714_, _31713_, _41806_);
  and _81989_ (_43659_, _31714_, _31712_);
  not _81990_ (_31715_, \oc8051_golden_model_1.TMOD [2]);
  nor _81991_ (_31716_, _05286_, _31715_);
  nor _81992_ (_31718_, _12538_, _11236_);
  nor _81993_ (_31719_, _31718_, _31716_);
  nor _81994_ (_31720_, _31719_, _07793_);
  and _81995_ (_31721_, _12539_, _05286_);
  nor _81996_ (_31722_, _31721_, _31716_);
  nor _81997_ (_31723_, _31722_, _07778_);
  and _81998_ (_31724_, _05286_, \oc8051_golden_model_1.ACC [2]);
  nor _81999_ (_31725_, _31724_, _31716_);
  nor _82000_ (_31726_, _31725_, _03737_);
  nor _82001_ (_31727_, _31725_, _09029_);
  nor _82002_ (_31729_, _04409_, _31715_);
  or _82003_ (_31730_, _31729_, _31727_);
  and _82004_ (_31731_, _31730_, _04081_);
  nor _82005_ (_31732_, _12416_, _11236_);
  nor _82006_ (_31733_, _31732_, _31716_);
  nor _82007_ (_31734_, _31733_, _04081_);
  or _82008_ (_31735_, _31734_, _31731_);
  and _82009_ (_31736_, _31735_, _03996_);
  nor _82010_ (_31737_, _11236_, _04875_);
  nor _82011_ (_31738_, _31737_, _31716_);
  nor _82012_ (_31740_, _31738_, _03996_);
  nor _82013_ (_31741_, _31740_, _31736_);
  nor _82014_ (_31742_, _31741_, _03729_);
  or _82015_ (_31743_, _31742_, _07390_);
  nor _82016_ (_31744_, _31743_, _31726_);
  and _82017_ (_31745_, _31738_, _07390_);
  nor _82018_ (_31746_, _31745_, _31744_);
  nor _82019_ (_31747_, _31746_, _04481_);
  and _82020_ (_31748_, _06637_, _05286_);
  nor _82021_ (_31749_, _31716_, _07400_);
  not _82022_ (_31751_, _31749_);
  nor _82023_ (_31752_, _31751_, _31748_);
  nor _82024_ (_31753_, _31752_, _03222_);
  not _82025_ (_31754_, _31753_);
  nor _82026_ (_31755_, _31754_, _31747_);
  nor _82027_ (_31756_, _12519_, _11236_);
  nor _82028_ (_31757_, _31756_, _31716_);
  nor _82029_ (_31758_, _31757_, _03589_);
  or _82030_ (_31759_, _31758_, _08828_);
  or _82031_ (_31760_, _31759_, _31755_);
  and _82032_ (_31762_, _12533_, _05286_);
  or _82033_ (_31763_, _31716_, _07766_);
  or _82034_ (_31764_, _31763_, _31762_);
  and _82035_ (_31765_, _05286_, _06332_);
  nor _82036_ (_31766_, _31765_, _31716_);
  and _82037_ (_31767_, _31766_, _03601_);
  nor _82038_ (_31768_, _31767_, _03780_);
  and _82039_ (_31769_, _31768_, _31764_);
  and _82040_ (_31770_, _31769_, _31760_);
  nor _82041_ (_31771_, _31770_, _31723_);
  nor _82042_ (_31773_, _31771_, _03622_);
  nor _82043_ (_31774_, _31716_, _05718_);
  not _82044_ (_31775_, _31774_);
  nor _82045_ (_31776_, _31766_, _07777_);
  and _82046_ (_31777_, _31776_, _31775_);
  nor _82047_ (_31778_, _31777_, _31773_);
  nor _82048_ (_31779_, _31778_, _03790_);
  nor _82049_ (_31780_, _31725_, _06828_);
  and _82050_ (_31781_, _31780_, _31775_);
  nor _82051_ (_31782_, _31781_, _03624_);
  not _82052_ (_31784_, _31782_);
  nor _82053_ (_31785_, _31784_, _31779_);
  nor _82054_ (_31786_, _12532_, _11236_);
  or _82055_ (_31787_, _31716_, _07795_);
  nor _82056_ (_31788_, _31787_, _31786_);
  or _82057_ (_31789_, _31788_, _03785_);
  nor _82058_ (_31790_, _31789_, _31785_);
  nor _82059_ (_31791_, _31790_, _31720_);
  nor _82060_ (_31792_, _31791_, _03815_);
  nor _82061_ (_31793_, _31733_, _04246_);
  or _82062_ (_31795_, _31793_, _03447_);
  nor _82063_ (_31796_, _31795_, _31792_);
  and _82064_ (_31797_, _12592_, _05286_);
  or _82065_ (_31798_, _31716_, _03514_);
  nor _82066_ (_31799_, _31798_, _31797_);
  nor _82067_ (_31800_, _31799_, _31796_);
  or _82068_ (_31801_, _31800_, _43004_);
  or _82069_ (_31802_, _43000_, \oc8051_golden_model_1.TMOD [2]);
  and _82070_ (_31803_, _31802_, _41806_);
  and _82071_ (_43660_, _31803_, _31801_);
  not _82072_ (_31805_, \oc8051_golden_model_1.TMOD [3]);
  nor _82073_ (_31806_, _05286_, _31805_);
  nor _82074_ (_31807_, _12738_, _11236_);
  nor _82075_ (_31808_, _31807_, _31806_);
  nor _82076_ (_31809_, _31808_, _07793_);
  and _82077_ (_31810_, _12739_, _05286_);
  nor _82078_ (_31811_, _31810_, _31806_);
  nor _82079_ (_31812_, _31811_, _07778_);
  and _82080_ (_31813_, _06592_, _05286_);
  or _82081_ (_31814_, _31813_, _31806_);
  and _82082_ (_31816_, _31814_, _04481_);
  and _82083_ (_31817_, _05286_, \oc8051_golden_model_1.ACC [3]);
  nor _82084_ (_31818_, _31817_, _31806_);
  nor _82085_ (_31819_, _31818_, _03737_);
  nor _82086_ (_31820_, _31818_, _09029_);
  nor _82087_ (_31821_, _04409_, _31805_);
  or _82088_ (_31822_, _31821_, _31820_);
  and _82089_ (_31823_, _31822_, _04081_);
  nor _82090_ (_31824_, _12627_, _11236_);
  nor _82091_ (_31825_, _31824_, _31806_);
  nor _82092_ (_31827_, _31825_, _04081_);
  or _82093_ (_31828_, _31827_, _31823_);
  and _82094_ (_31829_, _31828_, _03996_);
  nor _82095_ (_31830_, _11236_, _05005_);
  nor _82096_ (_31831_, _31830_, _31806_);
  nor _82097_ (_31832_, _31831_, _03996_);
  nor _82098_ (_31833_, _31832_, _31829_);
  nor _82099_ (_31834_, _31833_, _03729_);
  or _82100_ (_31835_, _31834_, _07390_);
  nor _82101_ (_31836_, _31835_, _31819_);
  and _82102_ (_31838_, _31831_, _07390_);
  or _82103_ (_31839_, _31838_, _04481_);
  nor _82104_ (_31840_, _31839_, _31836_);
  or _82105_ (_31841_, _31840_, _31816_);
  and _82106_ (_31842_, _31841_, _03589_);
  nor _82107_ (_31843_, _12718_, _11236_);
  nor _82108_ (_31844_, _31843_, _31806_);
  nor _82109_ (_31845_, _31844_, _03589_);
  or _82110_ (_31846_, _31845_, _08828_);
  or _82111_ (_31847_, _31846_, _31842_);
  and _82112_ (_31849_, _12733_, _05286_);
  or _82113_ (_31850_, _31806_, _07766_);
  or _82114_ (_31851_, _31850_, _31849_);
  and _82115_ (_31852_, _05286_, _06276_);
  nor _82116_ (_31853_, _31852_, _31806_);
  and _82117_ (_31854_, _31853_, _03601_);
  nor _82118_ (_31855_, _31854_, _03780_);
  and _82119_ (_31856_, _31855_, _31851_);
  and _82120_ (_31857_, _31856_, _31847_);
  nor _82121_ (_31858_, _31857_, _31812_);
  nor _82122_ (_31860_, _31858_, _03622_);
  nor _82123_ (_31861_, _31806_, _05567_);
  not _82124_ (_31862_, _31861_);
  nor _82125_ (_31863_, _31853_, _07777_);
  and _82126_ (_31864_, _31863_, _31862_);
  nor _82127_ (_31865_, _31864_, _31860_);
  nor _82128_ (_31866_, _31865_, _03790_);
  nor _82129_ (_31867_, _31818_, _06828_);
  and _82130_ (_31868_, _31867_, _31862_);
  or _82131_ (_31869_, _31868_, _31866_);
  and _82132_ (_31871_, _31869_, _07795_);
  nor _82133_ (_31872_, _12732_, _11236_);
  nor _82134_ (_31873_, _31872_, _31806_);
  nor _82135_ (_31874_, _31873_, _07795_);
  or _82136_ (_31875_, _31874_, _31871_);
  and _82137_ (_31876_, _31875_, _07793_);
  nor _82138_ (_31877_, _31876_, _31809_);
  nor _82139_ (_31878_, _31877_, _03815_);
  nor _82140_ (_31879_, _31825_, _04246_);
  or _82141_ (_31880_, _31879_, _03447_);
  nor _82142_ (_31882_, _31880_, _31878_);
  and _82143_ (_31883_, _12794_, _05286_);
  or _82144_ (_31884_, _31806_, _03514_);
  nor _82145_ (_31885_, _31884_, _31883_);
  nor _82146_ (_31886_, _31885_, _31882_);
  or _82147_ (_31887_, _31886_, _43004_);
  or _82148_ (_31888_, _43000_, \oc8051_golden_model_1.TMOD [3]);
  and _82149_ (_31889_, _31888_, _41806_);
  and _82150_ (_43663_, _31889_, _31887_);
  not _82151_ (_31890_, \oc8051_golden_model_1.TMOD [4]);
  nor _82152_ (_31892_, _05286_, _31890_);
  nor _82153_ (_31893_, _12816_, _11236_);
  nor _82154_ (_31894_, _31893_, _31892_);
  nor _82155_ (_31895_, _31894_, _07793_);
  and _82156_ (_31896_, _12817_, _05286_);
  nor _82157_ (_31897_, _31896_, _31892_);
  nor _82158_ (_31898_, _31897_, _07778_);
  and _82159_ (_31899_, _06298_, _05286_);
  nor _82160_ (_31900_, _31899_, _31892_);
  and _82161_ (_31901_, _31900_, _03601_);
  and _82162_ (_31903_, _05286_, \oc8051_golden_model_1.ACC [4]);
  nor _82163_ (_31904_, _31903_, _31892_);
  nor _82164_ (_31905_, _31904_, _03737_);
  nor _82165_ (_31906_, _31904_, _09029_);
  nor _82166_ (_31907_, _04409_, _31890_);
  or _82167_ (_31908_, _31907_, _31906_);
  and _82168_ (_31909_, _31908_, _04081_);
  nor _82169_ (_31910_, _12841_, _11236_);
  nor _82170_ (_31911_, _31910_, _31892_);
  nor _82171_ (_31912_, _31911_, _04081_);
  or _82172_ (_31914_, _31912_, _31909_);
  and _82173_ (_31915_, _31914_, _03996_);
  nor _82174_ (_31916_, _05777_, _11236_);
  nor _82175_ (_31917_, _31916_, _31892_);
  nor _82176_ (_31918_, _31917_, _03996_);
  nor _82177_ (_31919_, _31918_, _31915_);
  nor _82178_ (_31920_, _31919_, _03729_);
  or _82179_ (_31921_, _31920_, _07390_);
  nor _82180_ (_31922_, _31921_, _31905_);
  and _82181_ (_31923_, _31917_, _07390_);
  nor _82182_ (_31925_, _31923_, _31922_);
  nor _82183_ (_31926_, _31925_, _04481_);
  and _82184_ (_31927_, _06730_, _05286_);
  nor _82185_ (_31928_, _31892_, _07400_);
  not _82186_ (_31929_, _31928_);
  nor _82187_ (_31930_, _31929_, _31927_);
  or _82188_ (_31931_, _31930_, _03222_);
  nor _82189_ (_31932_, _31931_, _31926_);
  nor _82190_ (_31933_, _12933_, _11236_);
  nor _82191_ (_31934_, _31933_, _31892_);
  nor _82192_ (_31936_, _31934_, _03589_);
  or _82193_ (_31937_, _31936_, _03601_);
  nor _82194_ (_31938_, _31937_, _31932_);
  nor _82195_ (_31939_, _31938_, _31901_);
  or _82196_ (_31940_, _31939_, _03600_);
  and _82197_ (_31941_, _12821_, _05286_);
  or _82198_ (_31942_, _31941_, _31892_);
  or _82199_ (_31943_, _31942_, _07766_);
  and _82200_ (_31944_, _31943_, _07778_);
  and _82201_ (_31945_, _31944_, _31940_);
  nor _82202_ (_31947_, _31945_, _31898_);
  nor _82203_ (_31948_, _31947_, _03622_);
  nor _82204_ (_31949_, _31892_, _05825_);
  not _82205_ (_31950_, _31949_);
  nor _82206_ (_31951_, _31900_, _07777_);
  and _82207_ (_31952_, _31951_, _31950_);
  nor _82208_ (_31953_, _31952_, _31948_);
  nor _82209_ (_31954_, _31953_, _03790_);
  nor _82210_ (_31955_, _31904_, _06828_);
  and _82211_ (_31956_, _31955_, _31950_);
  nor _82212_ (_31958_, _31956_, _03624_);
  not _82213_ (_31959_, _31958_);
  nor _82214_ (_31960_, _31959_, _31954_);
  nor _82215_ (_31961_, _12819_, _11236_);
  or _82216_ (_31962_, _31892_, _07795_);
  nor _82217_ (_31963_, _31962_, _31961_);
  or _82218_ (_31964_, _31963_, _03785_);
  nor _82219_ (_31965_, _31964_, _31960_);
  nor _82220_ (_31966_, _31965_, _31895_);
  nor _82221_ (_31967_, _31966_, _03815_);
  nor _82222_ (_31969_, _31911_, _04246_);
  or _82223_ (_31970_, _31969_, _03447_);
  nor _82224_ (_31971_, _31970_, _31967_);
  and _82225_ (_31972_, _13003_, _05286_);
  or _82226_ (_31973_, _31892_, _03514_);
  nor _82227_ (_31974_, _31973_, _31972_);
  nor _82228_ (_31975_, _31974_, _31971_);
  or _82229_ (_31976_, _31975_, _43004_);
  or _82230_ (_31977_, _43000_, \oc8051_golden_model_1.TMOD [4]);
  and _82231_ (_31978_, _31977_, _41806_);
  and _82232_ (_43664_, _31978_, _31976_);
  not _82233_ (_31980_, \oc8051_golden_model_1.TMOD [5]);
  nor _82234_ (_31981_, _05286_, _31980_);
  nor _82235_ (_31982_, _13146_, _11236_);
  nor _82236_ (_31983_, _31982_, _31981_);
  nor _82237_ (_31984_, _31983_, _07793_);
  and _82238_ (_31985_, _13147_, _05286_);
  nor _82239_ (_31986_, _31985_, _31981_);
  nor _82240_ (_31987_, _31986_, _07778_);
  and _82241_ (_31988_, _06684_, _05286_);
  or _82242_ (_31990_, _31988_, _31981_);
  and _82243_ (_31991_, _31990_, _04481_);
  and _82244_ (_31992_, _05286_, \oc8051_golden_model_1.ACC [5]);
  nor _82245_ (_31993_, _31992_, _31981_);
  nor _82246_ (_31994_, _31993_, _03737_);
  nor _82247_ (_31995_, _31993_, _09029_);
  nor _82248_ (_31996_, _04409_, _31980_);
  or _82249_ (_31997_, _31996_, _31995_);
  and _82250_ (_31998_, _31997_, _04081_);
  nor _82251_ (_31999_, _13014_, _11236_);
  nor _82252_ (_32001_, _31999_, _31981_);
  nor _82253_ (_32002_, _32001_, _04081_);
  or _82254_ (_32003_, _32002_, _31998_);
  and _82255_ (_32004_, _32003_, _03996_);
  nor _82256_ (_32005_, _05469_, _11236_);
  nor _82257_ (_32006_, _32005_, _31981_);
  nor _82258_ (_32007_, _32006_, _03996_);
  nor _82259_ (_32008_, _32007_, _32004_);
  nor _82260_ (_32009_, _32008_, _03729_);
  or _82261_ (_32010_, _32009_, _07390_);
  nor _82262_ (_32012_, _32010_, _31994_);
  and _82263_ (_32013_, _32006_, _07390_);
  or _82264_ (_32014_, _32013_, _04481_);
  nor _82265_ (_32015_, _32014_, _32012_);
  or _82266_ (_32016_, _32015_, _31991_);
  and _82267_ (_32017_, _32016_, _03589_);
  nor _82268_ (_32018_, _13127_, _11236_);
  nor _82269_ (_32019_, _32018_, _31981_);
  nor _82270_ (_32020_, _32019_, _03589_);
  or _82271_ (_32021_, _32020_, _08828_);
  or _82272_ (_32023_, _32021_, _32017_);
  and _82273_ (_32024_, _13141_, _05286_);
  or _82274_ (_32025_, _31981_, _07766_);
  or _82275_ (_32026_, _32025_, _32024_);
  and _82276_ (_32027_, _06306_, _05286_);
  nor _82277_ (_32028_, _32027_, _31981_);
  and _82278_ (_32029_, _32028_, _03601_);
  nor _82279_ (_32030_, _32029_, _03780_);
  and _82280_ (_32031_, _32030_, _32026_);
  and _82281_ (_32032_, _32031_, _32023_);
  nor _82282_ (_32034_, _32032_, _31987_);
  nor _82283_ (_32035_, _32034_, _03622_);
  nor _82284_ (_32036_, _31981_, _05518_);
  not _82285_ (_32037_, _32036_);
  nor _82286_ (_32038_, _32028_, _07777_);
  and _82287_ (_32039_, _32038_, _32037_);
  nor _82288_ (_32040_, _32039_, _32035_);
  nor _82289_ (_32041_, _32040_, _03790_);
  nor _82290_ (_32042_, _31993_, _06828_);
  and _82291_ (_32043_, _32042_, _32037_);
  or _82292_ (_32045_, _32043_, _32041_);
  and _82293_ (_32046_, _32045_, _07795_);
  nor _82294_ (_32047_, _13140_, _11236_);
  nor _82295_ (_32048_, _32047_, _31981_);
  nor _82296_ (_32049_, _32048_, _07795_);
  or _82297_ (_32050_, _32049_, _32046_);
  and _82298_ (_32051_, _32050_, _07793_);
  nor _82299_ (_32052_, _32051_, _31984_);
  nor _82300_ (_32053_, _32052_, _03815_);
  nor _82301_ (_32054_, _32001_, _04246_);
  or _82302_ (_32056_, _32054_, _03447_);
  nor _82303_ (_32057_, _32056_, _32053_);
  and _82304_ (_32058_, _13199_, _05286_);
  or _82305_ (_32059_, _31981_, _03514_);
  nor _82306_ (_32060_, _32059_, _32058_);
  nor _82307_ (_32061_, _32060_, _32057_);
  or _82308_ (_32062_, _32061_, _43004_);
  or _82309_ (_32063_, _43000_, \oc8051_golden_model_1.TMOD [5]);
  and _82310_ (_32064_, _32063_, _41806_);
  and _82311_ (_43665_, _32064_, _32062_);
  not _82312_ (_32066_, \oc8051_golden_model_1.TMOD [6]);
  nor _82313_ (_32067_, _05286_, _32066_);
  nor _82314_ (_32068_, _13352_, _11236_);
  nor _82315_ (_32069_, _32068_, _32067_);
  nor _82316_ (_32070_, _32069_, _07793_);
  and _82317_ (_32071_, _13353_, _05286_);
  nor _82318_ (_32072_, _32071_, _32067_);
  nor _82319_ (_32073_, _32072_, _07778_);
  and _82320_ (_32074_, _06455_, _05286_);
  or _82321_ (_32075_, _32074_, _32067_);
  and _82322_ (_32077_, _32075_, _04481_);
  and _82323_ (_32078_, _05286_, \oc8051_golden_model_1.ACC [6]);
  nor _82324_ (_32079_, _32078_, _32067_);
  nor _82325_ (_32080_, _32079_, _03737_);
  nor _82326_ (_32081_, _32079_, _09029_);
  nor _82327_ (_32082_, _04409_, _32066_);
  or _82328_ (_32083_, _32082_, _32081_);
  and _82329_ (_32084_, _32083_, _04081_);
  nor _82330_ (_32085_, _13242_, _11236_);
  nor _82331_ (_32086_, _32085_, _32067_);
  nor _82332_ (_32088_, _32086_, _04081_);
  or _82333_ (_32089_, _32088_, _32084_);
  and _82334_ (_32090_, _32089_, _03996_);
  nor _82335_ (_32091_, _05363_, _11236_);
  nor _82336_ (_32092_, _32091_, _32067_);
  nor _82337_ (_32093_, _32092_, _03996_);
  nor _82338_ (_32094_, _32093_, _32090_);
  nor _82339_ (_32095_, _32094_, _03729_);
  or _82340_ (_32096_, _32095_, _07390_);
  nor _82341_ (_32097_, _32096_, _32080_);
  and _82342_ (_32099_, _32092_, _07390_);
  or _82343_ (_32100_, _32099_, _04481_);
  nor _82344_ (_32101_, _32100_, _32097_);
  or _82345_ (_32102_, _32101_, _32077_);
  and _82346_ (_32103_, _32102_, _03589_);
  nor _82347_ (_32104_, _13332_, _11236_);
  nor _82348_ (_32105_, _32104_, _32067_);
  nor _82349_ (_32106_, _32105_, _03589_);
  or _82350_ (_32107_, _32106_, _08828_);
  or _82351_ (_32108_, _32107_, _32103_);
  and _82352_ (_32110_, _13347_, _05286_);
  or _82353_ (_32111_, _32067_, _07766_);
  or _82354_ (_32112_, _32111_, _32110_);
  and _82355_ (_32113_, _13339_, _05286_);
  nor _82356_ (_32114_, _32113_, _32067_);
  and _82357_ (_32115_, _32114_, _03601_);
  nor _82358_ (_32116_, _32115_, _03780_);
  and _82359_ (_32117_, _32116_, _32112_);
  and _82360_ (_32118_, _32117_, _32108_);
  nor _82361_ (_32119_, _32118_, _32073_);
  nor _82362_ (_32121_, _32119_, _03622_);
  nor _82363_ (_32122_, _32067_, _05412_);
  not _82364_ (_32123_, _32122_);
  nor _82365_ (_32124_, _32114_, _07777_);
  and _82366_ (_32125_, _32124_, _32123_);
  nor _82367_ (_32126_, _32125_, _32121_);
  nor _82368_ (_32127_, _32126_, _03790_);
  nor _82369_ (_32128_, _32079_, _06828_);
  and _82370_ (_32129_, _32128_, _32123_);
  or _82371_ (_32130_, _32129_, _32127_);
  and _82372_ (_32132_, _32130_, _07795_);
  nor _82373_ (_32133_, _13346_, _11236_);
  nor _82374_ (_32134_, _32133_, _32067_);
  nor _82375_ (_32135_, _32134_, _07795_);
  or _82376_ (_32136_, _32135_, _32132_);
  and _82377_ (_32137_, _32136_, _07793_);
  nor _82378_ (_32138_, _32137_, _32070_);
  nor _82379_ (_32139_, _32138_, _03815_);
  nor _82380_ (_32140_, _32086_, _04246_);
  or _82381_ (_32141_, _32140_, _03447_);
  nor _82382_ (_32143_, _32141_, _32139_);
  and _82383_ (_32144_, _13402_, _05286_);
  or _82384_ (_32145_, _32067_, _03514_);
  nor _82385_ (_32146_, _32145_, _32144_);
  nor _82386_ (_32147_, _32146_, _32143_);
  or _82387_ (_32148_, _32147_, _43004_);
  or _82388_ (_32149_, _43000_, \oc8051_golden_model_1.TMOD [6]);
  and _82389_ (_32150_, _32149_, _41806_);
  and _82390_ (_43666_, _32150_, _32148_);
  and _82391_ (_32151_, _11975_, _02905_);
  nor _82392_ (_32153_, _03631_, _03196_);
  not _82393_ (_32154_, _32153_);
  and _82394_ (_32155_, _32154_, _04163_);
  and _82395_ (_32156_, _09854_, \oc8051_golden_model_1.PC [0]);
  and _82396_ (_32157_, _04163_, \oc8051_golden_model_1.PC [0]);
  nor _82397_ (_32158_, _32157_, _11444_);
  nor _82398_ (_32159_, _32158_, _09854_);
  nor _82399_ (_32160_, _32159_, _32156_);
  and _82400_ (_32161_, _32160_, _03453_);
  and _82401_ (_32162_, _11933_, _11940_);
  nor _82402_ (_32164_, _32162_, _02905_);
  not _82403_ (_32165_, _03203_);
  and _82404_ (_32166_, _11328_, _08733_);
  nor _82405_ (_32167_, _32166_, _02905_);
  not _82406_ (_32168_, _03201_);
  and _82407_ (_32169_, _11335_, _07795_);
  nor _82408_ (_32170_, _32169_, _02905_);
  not _82409_ (_32171_, _03192_);
  and _82410_ (_32172_, _11851_, _07777_);
  nor _82411_ (_32173_, _32172_, _02905_);
  not _82412_ (_32175_, _03182_);
  and _82413_ (_32176_, _11345_, _07766_);
  nor _82414_ (_32177_, _32176_, _02905_);
  and _82415_ (_32178_, _03601_, _02905_);
  nor _82416_ (_32179_, _03625_, _03222_);
  and _82417_ (_32180_, _32179_, _11756_);
  nor _82418_ (_32181_, _32180_, _02905_);
  nor _82419_ (_32182_, _04163_, _03227_);
  nor _82420_ (_32183_, _04163_, _03233_);
  and _82421_ (_32184_, _04163_, _03980_);
  nor _82422_ (_32186_, _11630_, _02905_);
  nor _82423_ (_32187_, _11642_, _02905_);
  and _82424_ (_32188_, _11642_, _02905_);
  nor _82425_ (_32189_, _32188_, _32187_);
  and _82426_ (_32190_, _11630_, _04763_);
  not _82427_ (_32191_, _32190_);
  nor _82428_ (_32192_, _32191_, _32189_);
  nor _82429_ (_32193_, _32192_, _32186_);
  not _82430_ (_32194_, _32193_);
  nor _82431_ (_32195_, _32194_, _32184_);
  nor _82432_ (_32197_, _32195_, _06073_);
  and _82433_ (_32198_, _11504_, \oc8051_golden_model_1.PC [0]);
  and _82434_ (_32199_, _04048_, _02905_);
  nor _82435_ (_32200_, _32199_, _11571_);
  and _82436_ (_32201_, _32200_, _11624_);
  or _82437_ (_32202_, _32201_, _32198_);
  nor _82438_ (_32203_, _32202_, _06072_);
  nor _82439_ (_32204_, _32203_, _32197_);
  nor _82440_ (_32205_, _32204_, _04422_);
  and _82441_ (_32206_, _04422_, \oc8051_golden_model_1.PC [0]);
  nor _82442_ (_32208_, _32206_, _03610_);
  not _82443_ (_32209_, _32208_);
  nor _82444_ (_32210_, _32209_, _32205_);
  not _82445_ (_32211_, _32210_);
  not _82446_ (_32212_, _32158_);
  and _82447_ (_32213_, _32212_, _11367_);
  and _82448_ (_32214_, _05666_, _05566_);
  and _82449_ (_32215_, _32214_, _11366_);
  nand _82450_ (_32216_, _32215_, _12413_);
  nor _82451_ (_32217_, _32216_, _02905_);
  or _82452_ (_32219_, _32217_, _04081_);
  or _82453_ (_32220_, _32219_, _32213_);
  and _82454_ (_32221_, _32220_, _11362_);
  and _82455_ (_32222_, _32221_, _32211_);
  nor _82456_ (_32223_, _11362_, _02905_);
  nor _82457_ (_32224_, _32223_, _04768_);
  not _82458_ (_32225_, _32224_);
  nor _82459_ (_32226_, _32225_, _32222_);
  nor _82460_ (_32227_, _04163_, _03230_);
  and _82461_ (_32228_, _11666_, _11659_);
  not _82462_ (_32230_, _32228_);
  nor _82463_ (_32231_, _32230_, _32227_);
  not _82464_ (_32232_, _32231_);
  nor _82465_ (_32233_, _32232_, _32226_);
  nor _82466_ (_32234_, _32228_, _02905_);
  nor _82467_ (_32235_, _32234_, _11670_);
  not _82468_ (_32236_, _32235_);
  nor _82469_ (_32237_, _32236_, _32233_);
  or _82470_ (_32238_, _32237_, _09917_);
  nor _82471_ (_32239_, _32238_, _32183_);
  and _82472_ (_32241_, _09969_, _02905_);
  not _82473_ (_32242_, _32241_);
  nor _82474_ (_32243_, _32212_, _09969_);
  nor _82475_ (_32244_, _32243_, _09921_);
  and _82476_ (_32245_, _32244_, _32242_);
  or _82477_ (_32246_, _32245_, _03615_);
  or _82478_ (_32247_, _32246_, _32239_);
  and _82479_ (_32248_, _32247_, _09920_);
  and _82480_ (_32249_, _11685_, _02905_);
  and _82481_ (_32250_, _32158_, _10018_);
  or _82482_ (_32252_, _32250_, _32249_);
  nor _82483_ (_32253_, _32252_, _09920_);
  nor _82484_ (_32254_, _32253_, _32248_);
  and _82485_ (_32255_, _09876_, _02905_);
  nor _82486_ (_32256_, _32212_, _09876_);
  nor _82487_ (_32257_, _32256_, _32255_);
  nor _82488_ (_32258_, _32257_, _04107_);
  nor _82489_ (_32259_, _32258_, _32254_);
  nor _82490_ (_32260_, _32259_, _03604_);
  and _82491_ (_32261_, _10061_, _02905_);
  nor _82492_ (_32263_, _32212_, _10061_);
  or _82493_ (_32264_, _32263_, _32261_);
  and _82494_ (_32265_, _32264_, _03604_);
  or _82495_ (_32266_, _32265_, _32260_);
  and _82496_ (_32267_, _32266_, _11358_);
  and _82497_ (_32268_, _10025_, _02905_);
  or _82498_ (_32269_, _32268_, _32267_);
  and _82499_ (_32270_, _32269_, _03227_);
  or _82500_ (_32271_, _32270_, _11356_);
  nor _82501_ (_32272_, _32271_, _32182_);
  nor _82502_ (_32274_, _11355_, _02905_);
  nor _82503_ (_32275_, _32274_, _11727_);
  not _82504_ (_32276_, _32275_);
  nor _82505_ (_32277_, _32276_, _32272_);
  nor _82506_ (_32278_, _04163_, _03238_);
  and _82507_ (_32279_, _11350_, _03248_);
  not _82508_ (_32280_, _32279_);
  nor _82509_ (_32281_, _32280_, _32278_);
  not _82510_ (_32282_, _32281_);
  nor _82511_ (_32283_, _32282_, _32277_);
  nor _82512_ (_32284_, _32279_, _02905_);
  nor _82513_ (_32285_, _32284_, _03224_);
  not _82514_ (_32286_, _32285_);
  nor _82515_ (_32287_, _32286_, _32283_);
  nor _82516_ (_32288_, _04163_, _05897_);
  not _82517_ (_32289_, _32180_);
  nor _82518_ (_32290_, _32289_, _32288_);
  not _82519_ (_32291_, _32290_);
  nor _82520_ (_32292_, _32291_, _32287_);
  or _82521_ (_32293_, _32292_, _03169_);
  nor _82522_ (_32295_, _32293_, _32181_);
  nor _82523_ (_32296_, _04163_, _03170_);
  or _82524_ (_32297_, _32296_, _11764_);
  or _82525_ (_32298_, _32297_, _32295_);
  or _82526_ (_32299_, _32200_, _11765_);
  and _82527_ (_32300_, _32299_, _32298_);
  and _82528_ (_32301_, _32300_, _05886_);
  or _82529_ (_32302_, _32301_, _32178_);
  and _82530_ (_32303_, _32302_, _11348_);
  and _82531_ (_32304_, _11347_, _03329_);
  or _82532_ (_32306_, _32304_, _32303_);
  and _82533_ (_32307_, _32306_, _10736_);
  nor _82534_ (_32308_, _04163_, _10736_);
  or _82535_ (_32309_, _32308_, _32307_);
  and _82536_ (_32310_, _32309_, _11820_);
  not _82537_ (_32311_, _32176_);
  and _82538_ (_32312_, _08786_, \oc8051_golden_model_1.PC [0]);
  and _82539_ (_32313_, _32200_, _11826_);
  or _82540_ (_32314_, _32313_, _32312_);
  and _82541_ (_32315_, _32314_, _11819_);
  nor _82542_ (_32316_, _32315_, _32311_);
  not _82543_ (_32317_, _32316_);
  nor _82544_ (_32318_, _32317_, _32310_);
  nor _82545_ (_32319_, _32318_, _32177_);
  and _82546_ (_32320_, _32319_, _32175_);
  nor _82547_ (_32321_, _04163_, _32175_);
  or _82548_ (_32322_, _32321_, _32320_);
  and _82549_ (_32323_, _32322_, _11842_);
  not _82550_ (_32324_, _32172_);
  nor _82551_ (_32325_, _32200_, _11826_);
  nor _82552_ (_32328_, _08786_, \oc8051_golden_model_1.PC [0]);
  nor _82553_ (_32329_, _32328_, _11842_);
  not _82554_ (_32330_, _32329_);
  nor _82555_ (_32331_, _32330_, _32325_);
  nor _82556_ (_32332_, _32331_, _32324_);
  not _82557_ (_32333_, _32332_);
  nor _82558_ (_32334_, _32333_, _32323_);
  nor _82559_ (_32335_, _32334_, _32173_);
  and _82560_ (_32336_, _32335_, _32171_);
  nor _82561_ (_32337_, _04163_, _32171_);
  or _82562_ (_32339_, _32337_, _32336_);
  and _82563_ (_32340_, _32339_, _11338_);
  not _82564_ (_32341_, _32169_);
  and _82565_ (_32342_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and _82566_ (_32343_, _32200_, _07871_);
  or _82567_ (_32344_, _32343_, _32342_);
  and _82568_ (_32345_, _32344_, _11337_);
  nor _82569_ (_32346_, _32345_, _32341_);
  not _82570_ (_32347_, _32346_);
  nor _82571_ (_32348_, _32347_, _32340_);
  nor _82572_ (_32350_, _32348_, _32170_);
  and _82573_ (_32351_, _32350_, _32168_);
  nor _82574_ (_32352_, _04163_, _32168_);
  or _82575_ (_32353_, _32352_, _32351_);
  and _82576_ (_32354_, _32353_, _11881_);
  nor _82577_ (_32355_, _07955_, _02905_);
  and _82578_ (_32356_, _07955_, _02905_);
  nor _82579_ (_32357_, _32356_, _32355_);
  nor _82580_ (_32358_, _32357_, _11881_);
  and _82581_ (_32359_, _11330_, _08588_);
  not _82582_ (_32361_, _32359_);
  nor _82583_ (_32362_, _32361_, _32358_);
  not _82584_ (_32363_, _32362_);
  nor _82585_ (_32364_, _32363_, _32354_);
  nor _82586_ (_32365_, _32359_, _02905_);
  or _82587_ (_32366_, _32365_, _03798_);
  nor _82588_ (_32367_, _32366_, _32364_);
  and _82589_ (_32368_, _06546_, _03798_);
  or _82590_ (_32369_, _32368_, _32367_);
  and _82591_ (_32370_, _32369_, _06399_);
  nor _82592_ (_32372_, _04163_, _06399_);
  or _82593_ (_32373_, _32372_, _32370_);
  and _82594_ (_32374_, _32373_, _11903_);
  and _82595_ (_32375_, _32212_, _09854_);
  nor _82596_ (_32376_, _09854_, _02905_);
  or _82597_ (_32377_, _32376_, _11903_);
  or _82598_ (_32378_, _32377_, _32375_);
  and _82599_ (_32379_, _32378_, _32166_);
  not _82600_ (_32380_, _32379_);
  nor _82601_ (_32381_, _32380_, _32374_);
  nor _82602_ (_32383_, _32381_, _32167_);
  and _82603_ (_32384_, _32383_, _03516_);
  and _82604_ (_32385_, _06546_, _03515_);
  or _82605_ (_32386_, _32385_, _32384_);
  and _82606_ (_32387_, _32386_, _32165_);
  nor _82607_ (_32388_, _04163_, _32165_);
  nor _82608_ (_32389_, _32388_, _32387_);
  nor _82609_ (_32390_, _32389_, _03628_);
  not _82610_ (_32391_, _32162_);
  and _82611_ (_32392_, _32160_, _03628_);
  nor _82612_ (_32394_, _32392_, _32391_);
  not _82613_ (_32395_, _32394_);
  nor _82614_ (_32396_, _32395_, _32390_);
  nor _82615_ (_32397_, _32396_, _32164_);
  nor _82616_ (_32398_, _32397_, _05103_);
  and _82617_ (_32399_, _05103_, _04163_);
  nor _82618_ (_32400_, _32399_, _03453_);
  not _82619_ (_32401_, _32400_);
  nor _82620_ (_32402_, _32401_, _32398_);
  nor _82621_ (_32403_, _32402_, _32161_);
  and _82622_ (_32405_, _11957_, _11964_);
  not _82623_ (_32406_, _32405_);
  nor _82624_ (_32407_, _32406_, _32403_);
  nor _82625_ (_32408_, _32405_, \oc8051_golden_model_1.PC [0]);
  nor _82626_ (_32409_, _32408_, _32154_);
  not _82627_ (_32410_, _32409_);
  nor _82628_ (_32411_, _32410_, _32407_);
  or _82629_ (_32412_, _32411_, _11975_);
  nor _82630_ (_32413_, _32412_, _32155_);
  or _82631_ (_32414_, _32413_, _32151_);
  or _82632_ (_32416_, _32414_, _43004_);
  or _82633_ (_32417_, _43000_, \oc8051_golden_model_1.PC [0]);
  and _82634_ (_32418_, _32417_, _41806_);
  and _82635_ (_43667_, _32418_, _32416_);
  and _82636_ (_32419_, _11975_, _11442_);
  and _82637_ (_32420_, _03447_, _02878_);
  and _82638_ (_32421_, _09854_, _11442_);
  nor _82639_ (_32422_, _11446_, _11444_);
  nor _82640_ (_32423_, _32422_, _11447_);
  nor _82641_ (_32424_, _32423_, _09854_);
  nor _82642_ (_32426_, _32424_, _32421_);
  and _82643_ (_32427_, _32426_, _03453_);
  nor _82644_ (_32428_, _11940_, _11442_);
  nor _82645_ (_32429_, _05848_, _11442_);
  nor _82646_ (_32430_, _11328_, _11442_);
  nor _82647_ (_32431_, _11330_, _11442_);
  and _82648_ (_32432_, _15120_, _03275_);
  nor _82649_ (_32433_, _11851_, _11442_);
  nor _82650_ (_32434_, _11345_, _11442_);
  not _82651_ (_32435_, _04066_);
  nand _82652_ (_32437_, _08070_, _32435_);
  and _82653_ (_32438_, _32437_, _03223_);
  and _82654_ (_32439_, _08055_, _03275_);
  and _82655_ (_32440_, _10025_, _03275_);
  nor _82656_ (_32441_, _03617_, _03606_);
  nand _82657_ (_32442_, _09969_, _03275_);
  not _82658_ (_32443_, _32423_);
  or _82659_ (_32444_, _32443_, _09969_);
  and _82660_ (_32445_, _32444_, _32442_);
  and _82661_ (_32446_, _32445_, _09917_);
  nor _82662_ (_32448_, _11666_, _11442_);
  or _82663_ (_32449_, _32216_, _11442_);
  or _82664_ (_32450_, _32443_, _11369_);
  and _82665_ (_32451_, _32450_, _03610_);
  and _82666_ (_32452_, _32451_, _32449_);
  or _82667_ (_32453_, _11624_, \oc8051_golden_model_1.PC [1]);
  nor _82668_ (_32454_, _11573_, _11571_);
  nor _82669_ (_32455_, _32454_, _11574_);
  nand _82670_ (_32456_, _32455_, _11624_);
  and _82671_ (_32457_, _32456_, _06073_);
  and _82672_ (_32459_, _32457_, _32453_);
  nor _82673_ (_32460_, _11630_, _11442_);
  or _82674_ (_32461_, _04303_, _04763_);
  and _82675_ (_32462_, _04064_, _03275_);
  and _82676_ (_32463_, _04729_, \oc8051_golden_model_1.PC [0]);
  nor _82677_ (_32464_, _32463_, _04409_);
  nand _82678_ (_32465_, _32464_, \oc8051_golden_model_1.PC [1]);
  or _82679_ (_32466_, _32464_, \oc8051_golden_model_1.PC [1]);
  nand _82680_ (_32467_, _32466_, _32465_);
  nor _82681_ (_32468_, _32467_, _04064_);
  or _82682_ (_32470_, _32468_, _32462_);
  or _82683_ (_32471_, _32470_, _03980_);
  and _82684_ (_32472_, _32471_, _11630_);
  and _82685_ (_32473_, _32472_, _32461_);
  or _82686_ (_32474_, _32473_, _32460_);
  and _82687_ (_32475_, _32474_, _06072_);
  or _82688_ (_32476_, _32475_, _04422_);
  or _82689_ (_32477_, _32476_, _32459_);
  nand _82690_ (_32478_, _04422_, _11442_);
  and _82691_ (_32479_, _32478_, _04081_);
  and _82692_ (_32481_, _32479_, _32477_);
  or _82693_ (_32482_, _32481_, _32452_);
  and _82694_ (_32483_, _32482_, _11362_);
  nor _82695_ (_32484_, _11362_, _11442_);
  or _82696_ (_32485_, _32484_, _03715_);
  or _82697_ (_32486_, _32485_, _32483_);
  nand _82698_ (_32487_, _03715_, _02878_);
  and _82699_ (_32488_, _32487_, _03230_);
  and _82700_ (_32489_, _32488_, _32486_);
  and _82701_ (_32490_, _04303_, _04768_);
  or _82702_ (_32492_, _32490_, _03723_);
  or _82703_ (_32493_, _32492_, _32489_);
  nand _82704_ (_32494_, _03723_, _02878_);
  and _82705_ (_32495_, _32494_, _11659_);
  and _82706_ (_32496_, _32495_, _32493_);
  nor _82707_ (_32497_, _11659_, _11442_);
  or _82708_ (_32498_, _32497_, _03729_);
  or _82709_ (_32499_, _32498_, _32496_);
  nand _82710_ (_32500_, _03729_, _02878_);
  and _82711_ (_32501_, _32500_, _11666_);
  and _82712_ (_32503_, _32501_, _32499_);
  or _82713_ (_32504_, _32503_, _32448_);
  and _82714_ (_32505_, _32504_, _03736_);
  and _82715_ (_32506_, _03714_, \oc8051_golden_model_1.PC [1]);
  or _82716_ (_32507_, _32506_, _11670_);
  or _82717_ (_32508_, _32507_, _32505_);
  or _82718_ (_32509_, _04303_, _03233_);
  and _82719_ (_32510_, _32509_, _32508_);
  or _82720_ (_32511_, _32510_, _03508_);
  nand _82721_ (_32512_, _03508_, _02878_);
  and _82722_ (_32514_, _32512_, _09921_);
  and _82723_ (_32515_, _32514_, _32511_);
  or _82724_ (_32516_, _32515_, _32446_);
  and _82725_ (_32517_, _32516_, _32441_);
  or _82726_ (_32518_, _10018_, _11442_);
  not _82727_ (_32519_, _32441_);
  or _82728_ (_32520_, _32443_, _11685_);
  and _82729_ (_32521_, _32520_, _32519_);
  and _82730_ (_32522_, _32521_, _32518_);
  or _82731_ (_32523_, _32522_, _03615_);
  or _82732_ (_32525_, _32523_, _32517_);
  or _82733_ (_32526_, _32443_, _09876_);
  nand _82734_ (_32527_, _09876_, _03275_);
  and _82735_ (_32528_, _32527_, _32526_);
  or _82736_ (_32529_, _32528_, _04107_);
  and _82737_ (_32530_, _32529_, _32525_);
  or _82738_ (_32531_, _32530_, _03604_);
  and _82739_ (_32532_, _10061_, _11442_);
  nor _82740_ (_32533_, _32423_, _10061_);
  or _82741_ (_32534_, _32533_, _09856_);
  or _82742_ (_32536_, _32534_, _32532_);
  and _82743_ (_32537_, _32536_, _11358_);
  and _82744_ (_32538_, _32537_, _32531_);
  or _82745_ (_32539_, _32538_, _32440_);
  and _82746_ (_32540_, _32539_, _06840_);
  and _82747_ (_32541_, _03719_, \oc8051_golden_model_1.PC [1]);
  or _82748_ (_32542_, _32541_, _04766_);
  or _82749_ (_32543_, _32542_, _32540_);
  or _82750_ (_32544_, _04303_, _03227_);
  and _82751_ (_32545_, _23519_, _11706_);
  and _82752_ (_32547_, _32545_, _23262_);
  and _82753_ (_32548_, _32547_, _32544_);
  and _82754_ (_32549_, _32548_, _32543_);
  nor _82755_ (_32550_, _32547_, _02878_);
  or _82756_ (_32551_, _32550_, _32549_);
  and _82757_ (_32552_, _32551_, _11355_);
  nor _82758_ (_32553_, _11355_, _11442_);
  or _82759_ (_32554_, _32553_, _03753_);
  or _82760_ (_32555_, _32554_, _32552_);
  nand _82761_ (_32556_, _03753_, _02878_);
  and _82762_ (_32558_, _32556_, _03238_);
  and _82763_ (_32559_, _32558_, _32555_);
  and _82764_ (_32560_, _04303_, _11727_);
  or _82765_ (_32561_, _32560_, _03752_);
  or _82766_ (_32562_, _32561_, _32559_);
  and _82767_ (_32563_, _03752_, _02878_);
  nor _82768_ (_32564_, _32563_, _08055_);
  and _82769_ (_32565_, _32564_, _32562_);
  nor _82770_ (_32566_, _32565_, _32439_);
  nor _82771_ (_32567_, _32566_, _32438_);
  and _82772_ (_32569_, _32438_, _03275_);
  nor _82773_ (_32570_, _04727_, _03247_);
  or _82774_ (_32571_, _32570_, _32569_);
  or _82775_ (_32572_, _32571_, _32567_);
  nand _82776_ (_32573_, _32570_, _11442_);
  and _82777_ (_32574_, _32573_, _08186_);
  and _82778_ (_32575_, _32574_, _32572_);
  nor _82779_ (_32576_, _08186_, _02878_);
  or _82780_ (_32577_, _32576_, _07912_);
  or _82781_ (_32578_, _32577_, _32575_);
  or _82782_ (_32580_, _03275_, _03248_);
  and _82783_ (_32581_, _32580_, _03710_);
  and _82784_ (_32582_, _32581_, _32578_);
  and _82785_ (_32583_, _03505_, \oc8051_golden_model_1.PC [1]);
  or _82786_ (_32584_, _32583_, _32582_);
  and _82787_ (_32585_, _32584_, _05897_);
  and _82788_ (_32586_, _04303_, _03224_);
  or _82789_ (_32587_, _32586_, _03625_);
  or _82790_ (_32588_, _32587_, _32585_);
  nand _82791_ (_32589_, _03625_, _03275_);
  and _82792_ (_32591_, _32589_, _11749_);
  and _82793_ (_32592_, _32591_, _32588_);
  nor _82794_ (_32593_, _11749_, _02878_);
  or _82795_ (_32594_, _32593_, _03222_);
  or _82796_ (_32595_, _32594_, _32592_);
  nand _82797_ (_32596_, _03275_, _03222_);
  and _82798_ (_32597_, _32596_, _11756_);
  and _82799_ (_32598_, _32597_, _32595_);
  nor _82800_ (_32599_, _11756_, _11442_);
  or _82801_ (_32600_, _32599_, _03585_);
  or _82802_ (_32602_, _32600_, _32598_);
  nand _82803_ (_32603_, _03585_, _02878_);
  and _82804_ (_32604_, _32603_, _03170_);
  and _82805_ (_32605_, _32604_, _32602_);
  and _82806_ (_32606_, _04303_, _03169_);
  or _82807_ (_32607_, _32606_, _11764_);
  or _82808_ (_32608_, _32607_, _32605_);
  nand _82809_ (_32609_, _32455_, _11764_);
  and _82810_ (_32610_, _32609_, _05894_);
  and _82811_ (_32611_, _32610_, _32608_);
  nor _82812_ (_32613_, _03601_, \oc8051_golden_model_1.PC [1]);
  nor _82813_ (_32614_, _32613_, _05895_);
  or _82814_ (_32615_, _32614_, _32611_);
  nand _82815_ (_32616_, _03601_, _03275_);
  and _82816_ (_32617_, _32616_, _08364_);
  and _82817_ (_32618_, _32617_, _32615_);
  and _82818_ (_32619_, _08363_, \oc8051_golden_model_1.PC [1]);
  or _82819_ (_32620_, _32619_, _32618_);
  nand _82820_ (_32621_, _32620_, _11348_);
  nor _82821_ (_32622_, _11348_, _03345_);
  nor _82822_ (_32623_, _32622_, _03584_);
  nand _82823_ (_32624_, _32623_, _32621_);
  and _82824_ (_32625_, _03584_, _02878_);
  nor _82825_ (_32626_, _32625_, _03178_);
  nand _82826_ (_32627_, _32626_, _32624_);
  and _82827_ (_32628_, _04303_, _03178_);
  nor _82828_ (_32629_, _32628_, _11819_);
  nand _82829_ (_32630_, _32629_, _32627_);
  nor _82830_ (_32631_, _32455_, _08786_);
  and _82831_ (_32632_, _08786_, \oc8051_golden_model_1.PC [1]);
  nor _82832_ (_32635_, _32632_, _11820_);
  not _82833_ (_32636_, _32635_);
  nor _82834_ (_32637_, _32636_, _32631_);
  nor _82835_ (_32638_, _32637_, _11824_);
  and _82836_ (_32639_, _32638_, _32630_);
  or _82837_ (_32640_, _32639_, _32434_);
  nand _82838_ (_32641_, _32640_, _11341_);
  nor _82839_ (_32642_, _11341_, _02878_);
  nor _82840_ (_32643_, _32642_, _03600_);
  nand _82841_ (_32644_, _32643_, _32641_);
  and _82842_ (_32646_, _03600_, _03275_);
  nor _82843_ (_32647_, _32646_, _03780_);
  and _82844_ (_32648_, _32647_, _32644_);
  and _82845_ (_32649_, _03780_, \oc8051_golden_model_1.PC [1]);
  or _82846_ (_32650_, _32649_, _32648_);
  nand _82847_ (_32651_, _32650_, _32175_);
  and _82848_ (_32652_, _04303_, _03182_);
  nor _82849_ (_32653_, _32652_, _11841_);
  nand _82850_ (_32654_, _32653_, _32651_);
  nor _82851_ (_32655_, _32455_, _11826_);
  nor _82852_ (_32657_, _08786_, _02878_);
  nor _82853_ (_32658_, _32657_, _11842_);
  not _82854_ (_32659_, _32658_);
  nor _82855_ (_32660_, _32659_, _32655_);
  nor _82856_ (_32661_, _32660_, _11853_);
  and _82857_ (_32662_, _32661_, _32654_);
  or _82858_ (_32663_, _32662_, _32433_);
  nand _82859_ (_32664_, _32663_, _08430_);
  nor _82860_ (_32665_, _08430_, _02878_);
  nor _82861_ (_32666_, _32665_, _03622_);
  nand _82862_ (_32668_, _32666_, _32664_);
  and _82863_ (_32669_, _03622_, _03275_);
  nor _82864_ (_32670_, _32669_, _03790_);
  and _82865_ (_32671_, _32670_, _32668_);
  and _82866_ (_32672_, _03790_, \oc8051_golden_model_1.PC [1]);
  or _82867_ (_32673_, _32672_, _32671_);
  nand _82868_ (_32674_, _32673_, _32171_);
  and _82869_ (_32675_, _04303_, _03192_);
  nor _82870_ (_32676_, _32675_, _11337_);
  nand _82871_ (_32677_, _32676_, _32674_);
  and _82872_ (_32679_, \oc8051_golden_model_1.PSW [7], _02878_);
  and _82873_ (_32680_, _32455_, _07871_);
  or _82874_ (_32681_, _32680_, _32679_);
  and _82875_ (_32682_, _32681_, _11337_);
  nor _82876_ (_32683_, _32682_, _15120_);
  and _82877_ (_32684_, _32683_, _32677_);
  or _82878_ (_32685_, _32684_, _32432_);
  nand _82879_ (_32686_, _08450_, _12559_);
  nor _82880_ (_32687_, _15123_, _15127_);
  and _82881_ (_32688_, _32687_, _32686_);
  nand _82882_ (_32690_, _32688_, _32685_);
  and _82883_ (_32691_, _03605_, _03200_);
  nor _82884_ (_32692_, _32688_, _11442_);
  nor _82885_ (_32693_, _32692_, _32691_);
  nand _82886_ (_32694_, _32693_, _32690_);
  and _82887_ (_32695_, _32691_, _11442_);
  nor _82888_ (_32696_, _32695_, _08460_);
  nand _82889_ (_32697_, _32696_, _32694_);
  nor _82890_ (_32698_, _08459_, _02878_);
  nor _82891_ (_32699_, _32698_, _03624_);
  nand _82892_ (_32701_, _32699_, _32697_);
  and _82893_ (_32702_, _03624_, _03275_);
  nor _82894_ (_32703_, _32702_, _03785_);
  and _82895_ (_32704_, _32703_, _32701_);
  and _82896_ (_32705_, _03785_, \oc8051_golden_model_1.PC [1]);
  or _82897_ (_32706_, _32705_, _32704_);
  nand _82898_ (_32707_, _32706_, _32168_);
  and _82899_ (_32708_, _04303_, _03201_);
  nor _82900_ (_32709_, _32708_, _11880_);
  nand _82901_ (_32710_, _32709_, _32707_);
  nor _82902_ (_32712_, _32455_, _07871_);
  and _82903_ (_32713_, _07871_, \oc8051_golden_model_1.PC [1]);
  nor _82904_ (_32714_, _32713_, _11881_);
  not _82905_ (_32715_, _32714_);
  nor _82906_ (_32716_, _32715_, _32712_);
  nor _82907_ (_32717_, _32716_, _11885_);
  and _82908_ (_32718_, _32717_, _32710_);
  or _82909_ (_32719_, _32718_, _32431_);
  nand _82910_ (_32720_, _32719_, _08507_);
  nor _82911_ (_32721_, _08507_, _02878_);
  nor _82912_ (_32723_, _32721_, _08587_);
  nand _82913_ (_32724_, _32723_, _32720_);
  and _82914_ (_32725_, _08587_, _11442_);
  nor _82915_ (_32726_, _32725_, _03798_);
  and _82916_ (_32727_, _32726_, _32724_);
  nor _82917_ (_32728_, _06501_, _10652_);
  or _82918_ (_32729_, _32728_, _32727_);
  nand _82919_ (_32730_, _32729_, _06399_);
  and _82920_ (_32731_, _04303_, _03188_);
  nor _82921_ (_32732_, _32731_, _03621_);
  nand _82922_ (_32734_, _32732_, _32730_);
  nor _82923_ (_32735_, _09854_, _03275_);
  and _82924_ (_32736_, _32443_, _09854_);
  or _82925_ (_32737_, _32736_, _11903_);
  nor _82926_ (_32738_, _32737_, _32735_);
  nor _82927_ (_32739_, _32738_, _11907_);
  and _82928_ (_32740_, _32739_, _32734_);
  or _82929_ (_32741_, _32740_, _32430_);
  nand _82930_ (_32742_, _32741_, _08702_);
  nor _82931_ (_32743_, _08702_, _02878_);
  nor _82932_ (_32745_, _32743_, _08732_);
  nand _82933_ (_32746_, _32745_, _32742_);
  and _82934_ (_32747_, _08732_, _11442_);
  nor _82935_ (_32748_, _32747_, _03515_);
  and _82936_ (_32749_, _32748_, _32746_);
  nor _82937_ (_32750_, _06501_, _03516_);
  or _82938_ (_32751_, _32750_, _32749_);
  nand _82939_ (_32752_, _32751_, _32165_);
  and _82940_ (_32753_, _04303_, _03203_);
  nor _82941_ (_32754_, _32753_, _03628_);
  nand _82942_ (_32756_, _32754_, _32752_);
  and _82943_ (_32757_, _32426_, _03628_);
  nor _82944_ (_32758_, _32757_, _12561_);
  and _82945_ (_32759_, _32758_, _32756_);
  or _82946_ (_32760_, _32759_, _32429_);
  nand _82947_ (_32761_, _32760_, _06409_);
  and _82948_ (_32762_, _04533_, _03275_);
  nor _82949_ (_32763_, _32762_, _03815_);
  nand _82950_ (_32764_, _32763_, _32761_);
  not _82951_ (_32765_, _11940_);
  and _82952_ (_32767_, _03815_, _02878_);
  nor _82953_ (_32768_, _32767_, _32765_);
  and _82954_ (_32769_, _32768_, _32764_);
  or _82955_ (_32770_, _32769_, _32428_);
  nand _82956_ (_32771_, _32770_, _04540_);
  and _82957_ (_32772_, _05103_, _04303_);
  nor _82958_ (_32773_, _32772_, _03453_);
  and _82959_ (_32774_, _32773_, _32771_);
  or _82960_ (_32775_, _32774_, _32427_);
  nand _82961_ (_32776_, _32775_, _11955_);
  nor _82962_ (_32778_, _11955_, _03275_);
  nor _82963_ (_32779_, _32778_, _04552_);
  nand _82964_ (_32780_, _32779_, _32776_);
  and _82965_ (_32781_, _04552_, _03275_);
  nor _82966_ (_32782_, _32781_, _03447_);
  and _82967_ (_32783_, _32782_, _32780_);
  or _82968_ (_32784_, _32783_, _32420_);
  nand _82969_ (_32785_, _32784_, _11964_);
  nor _82970_ (_32786_, _11964_, _03275_);
  nor _82971_ (_32787_, _32786_, _32154_);
  nand _82972_ (_32789_, _32787_, _32785_);
  and _82973_ (_32790_, _32154_, _04303_);
  nor _82974_ (_32791_, _32790_, _11975_);
  and _82975_ (_32792_, _32791_, _32789_);
  or _82976_ (_32793_, _32792_, _32419_);
  or _82977_ (_32794_, _32793_, _43004_);
  or _82978_ (_32795_, _43000_, \oc8051_golden_model_1.PC [1]);
  and _82979_ (_32796_, _32795_, _41806_);
  and _82980_ (_43670_, _32796_, _32794_);
  and _82981_ (_32797_, _03447_, _03210_);
  nor _82982_ (_32799_, _11328_, _03266_);
  nor _82983_ (_32800_, _11330_, _03266_);
  nor _82984_ (_32801_, _11335_, _03266_);
  nor _82985_ (_32802_, _11851_, _03266_);
  nor _82986_ (_32803_, _11345_, _03266_);
  and _82987_ (_32804_, _03505_, _03245_);
  nor _82988_ (_32805_, _32547_, _03210_);
  not _82989_ (_32806_, _03266_);
  and _82990_ (_32807_, _10025_, _32806_);
  and _82991_ (_32808_, _03980_, _03946_);
  nor _82992_ (_32810_, _11643_, _03266_);
  and _82993_ (_32811_, _03979_, _03245_);
  or _82994_ (_32812_, _04409_, \oc8051_golden_model_1.PC [2]);
  nor _82995_ (_32813_, _32812_, _04729_);
  or _82996_ (_32814_, _32813_, _32811_);
  not _82997_ (_32815_, _11632_);
  and _82998_ (_32816_, _32190_, _32815_);
  and _82999_ (_32817_, _32816_, _32814_);
  or _83000_ (_32818_, _32817_, _32810_);
  or _83001_ (_32819_, _32818_, _32808_);
  and _83002_ (_32821_, _32819_, _06072_);
  and _83003_ (_32822_, _11578_, _11575_);
  nor _83004_ (_32823_, _32822_, _11579_);
  nand _83005_ (_32824_, _32823_, _11624_);
  or _83006_ (_32825_, _11624_, _03245_);
  and _83007_ (_32826_, _32825_, _06073_);
  and _83008_ (_32827_, _32826_, _32824_);
  or _83009_ (_32828_, _32827_, _32821_);
  and _83010_ (_32829_, _32828_, _05966_);
  and _83011_ (_32830_, _04422_, _32806_);
  or _83012_ (_32832_, _32830_, _03610_);
  or _83013_ (_32833_, _32832_, _32829_);
  and _83014_ (_32834_, _11451_, _11448_);
  nor _83015_ (_32835_, _32834_, _11452_);
  not _83016_ (_32836_, _32835_);
  and _83017_ (_32837_, _32836_, _11367_);
  and _83018_ (_32838_, _11440_, _11369_);
  or _83019_ (_32839_, _32838_, _04081_);
  or _83020_ (_32840_, _32839_, _32837_);
  and _83021_ (_32841_, _32840_, _11362_);
  and _83022_ (_32843_, _32841_, _32833_);
  nor _83023_ (_32844_, _11362_, _03266_);
  or _83024_ (_32845_, _32844_, _03715_);
  or _83025_ (_32846_, _32845_, _32843_);
  nand _83026_ (_32847_, _03715_, _03210_);
  and _83027_ (_32848_, _32847_, _03230_);
  and _83028_ (_32849_, _32848_, _32846_);
  and _83029_ (_32850_, _03946_, _04768_);
  or _83030_ (_32851_, _32850_, _03723_);
  or _83031_ (_32852_, _32851_, _32849_);
  nand _83032_ (_32854_, _03723_, _03210_);
  and _83033_ (_32855_, _32854_, _11659_);
  and _83034_ (_32856_, _32855_, _32852_);
  nor _83035_ (_32857_, _11659_, _03266_);
  or _83036_ (_32858_, _32857_, _03729_);
  or _83037_ (_32859_, _32858_, _32856_);
  nand _83038_ (_32860_, _03729_, _03210_);
  and _83039_ (_32861_, _32860_, _11666_);
  and _83040_ (_32862_, _32861_, _32859_);
  nor _83041_ (_32863_, _11666_, _03266_);
  or _83042_ (_32865_, _32863_, _03714_);
  or _83043_ (_32866_, _32865_, _32862_);
  nand _83044_ (_32867_, _03714_, _03210_);
  and _83045_ (_32868_, _32867_, _03233_);
  and _83046_ (_32869_, _32868_, _32866_);
  and _83047_ (_32870_, _03946_, _11670_);
  or _83048_ (_32871_, _32870_, _03508_);
  or _83049_ (_32872_, _32871_, _32869_);
  nand _83050_ (_32873_, _03508_, _03210_);
  and _83051_ (_32874_, _32873_, _09921_);
  and _83052_ (_32876_, _32874_, _32872_);
  or _83053_ (_32877_, _32836_, _09969_);
  nand _83054_ (_32878_, _11439_, _09969_);
  and _83055_ (_32879_, _32878_, _09917_);
  nand _83056_ (_32880_, _32879_, _32877_);
  nand _83057_ (_32881_, _32880_, _23483_);
  or _83058_ (_32882_, _32881_, _32876_);
  or _83059_ (_32883_, _32836_, _09876_);
  nand _83060_ (_32884_, _11439_, _09876_);
  and _83061_ (_32885_, _32884_, _32883_);
  or _83062_ (_32887_, _32885_, _04107_);
  or _83063_ (_32888_, _32836_, _11685_);
  or _83064_ (_32889_, _11440_, _10018_);
  and _83065_ (_32890_, _32889_, _32888_);
  or _83066_ (_32891_, _32890_, _09920_);
  and _83067_ (_32892_, _32891_, _32887_);
  and _83068_ (_32893_, _32892_, _32882_);
  or _83069_ (_32894_, _32893_, _03604_);
  and _83070_ (_32895_, _11440_, _10061_);
  nor _83071_ (_32896_, _32835_, _10061_);
  or _83072_ (_32898_, _32896_, _09856_);
  or _83073_ (_32899_, _32898_, _32895_);
  and _83074_ (_32900_, _32899_, _11358_);
  and _83075_ (_32901_, _32900_, _32894_);
  or _83076_ (_32902_, _32901_, _32807_);
  and _83077_ (_32903_, _32902_, _06840_);
  and _83078_ (_32904_, _03719_, _03245_);
  or _83079_ (_32905_, _32904_, _04766_);
  or _83080_ (_32906_, _32905_, _32903_);
  or _83081_ (_32907_, _03946_, _03227_);
  and _83082_ (_32909_, _32907_, _32547_);
  and _83083_ (_32910_, _32909_, _32906_);
  or _83084_ (_32911_, _32910_, _32805_);
  and _83085_ (_32912_, _32911_, _11355_);
  nor _83086_ (_32913_, _11355_, _03266_);
  or _83087_ (_32914_, _32913_, _03753_);
  or _83088_ (_32915_, _32914_, _32912_);
  nand _83089_ (_32916_, _03753_, _03210_);
  and _83090_ (_32917_, _32916_, _03238_);
  and _83091_ (_32918_, _32917_, _32915_);
  and _83092_ (_32920_, _03946_, _11727_);
  or _83093_ (_32921_, _32920_, _03752_);
  or _83094_ (_32922_, _32921_, _32918_);
  nand _83095_ (_32923_, _03752_, _03210_);
  and _83096_ (_32924_, _32923_, _11350_);
  and _83097_ (_32925_, _32924_, _32922_);
  nor _83098_ (_32926_, _11350_, _03266_);
  or _83099_ (_32927_, _32926_, _32925_);
  and _83100_ (_32928_, _32927_, _08186_);
  nor _83101_ (_32929_, _08186_, _03210_);
  or _83102_ (_32931_, _32929_, _07912_);
  or _83103_ (_32932_, _32931_, _32928_);
  or _83104_ (_32933_, _32806_, _03248_);
  and _83105_ (_32934_, _32933_, _03710_);
  and _83106_ (_32935_, _32934_, _32932_);
  or _83107_ (_32936_, _32935_, _32804_);
  and _83108_ (_32937_, _32936_, _05897_);
  and _83109_ (_32938_, _03946_, _03224_);
  or _83110_ (_32939_, _32938_, _03625_);
  or _83111_ (_32940_, _32939_, _32937_);
  and _83112_ (_32942_, _11439_, _03625_);
  nor _83113_ (_32943_, _32942_, _04475_);
  and _83114_ (_32944_, _32943_, _32940_);
  and _83115_ (_32945_, _04475_, _03245_);
  or _83116_ (_32946_, _06835_, _03969_);
  or _83117_ (_32947_, _32946_, _32945_);
  or _83118_ (_32948_, _32947_, _32944_);
  nand _83119_ (_32949_, _32946_, _03210_);
  and _83120_ (_32950_, _32949_, _11748_);
  and _83121_ (_32951_, _32950_, _32948_);
  nor _83122_ (_32953_, _11748_, _03210_);
  or _83123_ (_32954_, _32953_, _03222_);
  or _83124_ (_32955_, _32954_, _32951_);
  nand _83125_ (_32956_, _11439_, _03222_);
  and _83126_ (_32957_, _32956_, _11756_);
  and _83127_ (_32958_, _32957_, _32955_);
  nor _83128_ (_32959_, _11756_, _03266_);
  or _83129_ (_32960_, _32959_, _03585_);
  or _83130_ (_32961_, _32960_, _32958_);
  nand _83131_ (_32962_, _03585_, _03210_);
  and _83132_ (_32964_, _32962_, _03170_);
  and _83133_ (_32965_, _32964_, _32961_);
  and _83134_ (_32966_, _03946_, _03169_);
  or _83135_ (_32967_, _32966_, _32965_);
  and _83136_ (_32968_, _32967_, _11765_);
  nor _83137_ (_32969_, _32823_, _11765_);
  or _83138_ (_32970_, _32969_, _06168_);
  or _83139_ (_32971_, _32970_, _32968_);
  or _83140_ (_32972_, _05894_, _03245_);
  and _83141_ (_32973_, _32972_, _05886_);
  and _83142_ (_32974_, _32973_, _32971_);
  and _83143_ (_32975_, _11440_, _03601_);
  or _83144_ (_32976_, _32975_, _08363_);
  or _83145_ (_32977_, _32976_, _32974_);
  and _83146_ (_32978_, _08363_, _03210_);
  nor _83147_ (_32979_, _32978_, _11347_);
  and _83148_ (_32980_, _32979_, _32977_);
  and _83149_ (_32981_, _11347_, _03262_);
  or _83150_ (_32982_, _32981_, _03584_);
  or _83151_ (_32983_, _32982_, _32980_);
  nand _83152_ (_32986_, _03584_, _03210_);
  and _83153_ (_32987_, _32986_, _10736_);
  and _83154_ (_32988_, _32987_, _32983_);
  and _83155_ (_32989_, _03946_, _03178_);
  or _83156_ (_32990_, _32989_, _11819_);
  or _83157_ (_32991_, _32990_, _32988_);
  nor _83158_ (_32992_, _32823_, _08786_);
  nand _83159_ (_32993_, _08786_, _03245_);
  nand _83160_ (_32994_, _32993_, _11819_);
  or _83161_ (_32995_, _32994_, _32992_);
  and _83162_ (_32997_, _32995_, _11345_);
  and _83163_ (_32998_, _32997_, _32991_);
  or _83164_ (_32999_, _32998_, _32803_);
  and _83165_ (_33000_, _32999_, _11341_);
  nor _83166_ (_33001_, _11341_, _03210_);
  or _83167_ (_33002_, _33001_, _03600_);
  or _83168_ (_33003_, _33002_, _33000_);
  nand _83169_ (_33004_, _11439_, _03600_);
  and _83170_ (_33005_, _33004_, _07778_);
  and _83171_ (_33006_, _33005_, _33003_);
  and _83172_ (_33008_, _03780_, _03245_);
  or _83173_ (_33009_, _33008_, _33006_);
  and _83174_ (_33010_, _33009_, _32175_);
  and _83175_ (_33011_, _03946_, _03182_);
  or _83176_ (_33012_, _33011_, _11841_);
  or _83177_ (_33013_, _33012_, _33010_);
  or _83178_ (_33014_, _32823_, _11826_);
  or _83179_ (_33015_, _08786_, _03210_);
  and _83180_ (_33016_, _33015_, _11841_);
  and _83181_ (_33017_, _33016_, _33014_);
  nor _83182_ (_33019_, _33017_, _11853_);
  and _83183_ (_33020_, _33019_, _33013_);
  or _83184_ (_33021_, _33020_, _32802_);
  and _83185_ (_33022_, _33021_, _08430_);
  nor _83186_ (_33023_, _08430_, _03210_);
  or _83187_ (_33024_, _33023_, _03622_);
  or _83188_ (_33025_, _33024_, _33022_);
  nand _83189_ (_33026_, _11439_, _03622_);
  and _83190_ (_33027_, _33026_, _06828_);
  and _83191_ (_33028_, _33027_, _33025_);
  and _83192_ (_33029_, _03790_, _03245_);
  or _83193_ (_33030_, _33029_, _33028_);
  and _83194_ (_33031_, _33030_, _32171_);
  and _83195_ (_33032_, _03946_, _03192_);
  or _83196_ (_33033_, _33032_, _11337_);
  or _83197_ (_33034_, _33033_, _33031_);
  nor _83198_ (_33035_, _32823_, \oc8051_golden_model_1.PSW [7]);
  or _83199_ (_33036_, _03210_, _07871_);
  nand _83200_ (_33037_, _33036_, _11337_);
  or _83201_ (_33038_, _33037_, _33035_);
  and _83202_ (_33040_, _33038_, _11335_);
  and _83203_ (_33041_, _33040_, _33034_);
  or _83204_ (_33042_, _33041_, _32801_);
  and _83205_ (_33043_, _33042_, _08459_);
  nor _83206_ (_33044_, _08459_, _03210_);
  or _83207_ (_33045_, _33044_, _03624_);
  or _83208_ (_33046_, _33045_, _33043_);
  nand _83209_ (_33047_, _11439_, _03624_);
  and _83210_ (_33048_, _33047_, _07793_);
  and _83211_ (_33049_, _33048_, _33046_);
  and _83212_ (_33051_, _03785_, _03245_);
  or _83213_ (_33052_, _33051_, _33049_);
  and _83214_ (_33053_, _33052_, _32168_);
  and _83215_ (_33054_, _03946_, _03201_);
  or _83216_ (_33055_, _33054_, _11880_);
  or _83217_ (_33056_, _33055_, _33053_);
  nor _83218_ (_33057_, _32823_, _07871_);
  or _83219_ (_33058_, _03210_, \oc8051_golden_model_1.PSW [7]);
  nand _83220_ (_33059_, _33058_, _11880_);
  or _83221_ (_33060_, _33059_, _33057_);
  and _83222_ (_33062_, _33060_, _11330_);
  and _83223_ (_33063_, _33062_, _33056_);
  or _83224_ (_33064_, _33063_, _32800_);
  and _83225_ (_33065_, _33064_, _08507_);
  nor _83226_ (_33066_, _08507_, _03210_);
  or _83227_ (_33067_, _33066_, _08587_);
  or _83228_ (_33068_, _33067_, _33065_);
  nand _83229_ (_33069_, _08587_, _03266_);
  and _83230_ (_33070_, _33069_, _10652_);
  and _83231_ (_33071_, _33070_, _33068_);
  nor _83232_ (_33073_, _06637_, _10652_);
  or _83233_ (_33074_, _33073_, _33071_);
  and _83234_ (_33075_, _33074_, _06399_);
  and _83235_ (_33076_, _03946_, _03188_);
  or _83236_ (_33077_, _33076_, _03621_);
  or _83237_ (_33078_, _33077_, _33075_);
  and _83238_ (_33079_, _32836_, _09854_);
  nor _83239_ (_33080_, _11439_, _09854_);
  or _83240_ (_33081_, _33080_, _11903_);
  or _83241_ (_33082_, _33081_, _33079_);
  and _83242_ (_33084_, _33082_, _11328_);
  and _83243_ (_33085_, _33084_, _33078_);
  or _83244_ (_33086_, _33085_, _32799_);
  and _83245_ (_33087_, _33086_, _08702_);
  nor _83246_ (_33088_, _08702_, _03210_);
  or _83247_ (_33089_, _33088_, _08732_);
  or _83248_ (_33090_, _33089_, _33087_);
  nand _83249_ (_33091_, _08732_, _03266_);
  and _83250_ (_33092_, _33091_, _03516_);
  and _83251_ (_33093_, _33092_, _33090_);
  nor _83252_ (_33095_, _06637_, _03516_);
  or _83253_ (_33096_, _33095_, _33093_);
  and _83254_ (_33097_, _33096_, _32165_);
  and _83255_ (_33098_, _03946_, _03203_);
  or _83256_ (_33099_, _33098_, _03628_);
  or _83257_ (_33100_, _33099_, _33097_);
  nor _83258_ (_33101_, _32835_, _09854_);
  and _83259_ (_33102_, _11440_, _09854_);
  nor _83260_ (_33103_, _33102_, _33101_);
  nand _83261_ (_33104_, _33103_, _03628_);
  and _83262_ (_33106_, _33104_, _11933_);
  and _83263_ (_33107_, _33106_, _33100_);
  nor _83264_ (_33108_, _11933_, _03266_);
  or _83265_ (_33109_, _33108_, _03815_);
  or _83266_ (_33110_, _33109_, _33107_);
  and _83267_ (_33111_, _03815_, _03210_);
  nor _83268_ (_33112_, _33111_, _32765_);
  and _83269_ (_33113_, _33112_, _33110_);
  nor _83270_ (_33114_, _11940_, _03266_);
  or _83271_ (_33115_, _33114_, _33113_);
  and _83272_ (_33117_, _33115_, _04540_);
  and _83273_ (_33118_, _05103_, _03946_);
  nor _83274_ (_33119_, _33118_, _03453_);
  not _83275_ (_33120_, _33119_);
  or _83276_ (_33121_, _33120_, _33117_);
  and _83277_ (_33122_, _33103_, _03453_);
  nor _83278_ (_33123_, _33122_, _11958_);
  nand _83279_ (_33124_, _33123_, _33121_);
  nor _83280_ (_33125_, _11957_, _03266_);
  nor _83281_ (_33126_, _33125_, _03447_);
  and _83282_ (_33128_, _33126_, _33124_);
  or _83283_ (_33129_, _33128_, _32797_);
  nand _83284_ (_33130_, _33129_, _11964_);
  nor _83285_ (_33131_, _11964_, _32806_);
  nor _83286_ (_33132_, _33131_, _32154_);
  nand _83287_ (_33133_, _33132_, _33130_);
  and _83288_ (_33134_, _32154_, _03946_);
  nor _83289_ (_33135_, _33134_, _11975_);
  and _83290_ (_33136_, _33135_, _33133_);
  and _83291_ (_33137_, _11975_, _03266_);
  or _83292_ (_33139_, _33137_, _33136_);
  or _83293_ (_33140_, _33139_, _43004_);
  or _83294_ (_33141_, _43000_, \oc8051_golden_model_1.PC [2]);
  and _83295_ (_33142_, _33141_, _41806_);
  and _83296_ (_43671_, _33142_, _33140_);
  and _83297_ (_33143_, _03447_, _03297_);
  and _83298_ (_33144_, _03815_, _03297_);
  nor _83299_ (_33145_, _11328_, _03650_);
  nor _83300_ (_33146_, _11330_, _03650_);
  nor _83301_ (_33147_, _11335_, _03650_);
  nor _83302_ (_33149_, _11851_, _03650_);
  nor _83303_ (_33150_, _11345_, _03650_);
  and _83304_ (_33151_, _08363_, _03648_);
  and _83305_ (_33152_, _03505_, _03648_);
  nor _83306_ (_33153_, _11350_, _03650_);
  nor _83307_ (_33154_, _32547_, _03297_);
  and _83308_ (_33155_, _10025_, _03311_);
  and _83309_ (_33156_, _11504_, _03648_);
  or _83310_ (_33157_, _11568_, _11567_);
  and _83311_ (_33158_, _33157_, _11580_);
  nor _83312_ (_33160_, _33157_, _11580_);
  nor _83313_ (_33161_, _33160_, _33158_);
  not _83314_ (_33162_, _33161_);
  and _83315_ (_33163_, _33162_, _11624_);
  or _83316_ (_33164_, _33163_, _06072_);
  or _83317_ (_33165_, _33164_, _33156_);
  and _83318_ (_33166_, _03980_, _03708_);
  nor _83319_ (_33167_, _11642_, _03650_);
  and _83320_ (_33168_, _03979_, _03648_);
  not _83321_ (_33169_, _04729_);
  nor _83322_ (_33171_, _04409_, \oc8051_golden_model_1.PC [3]);
  and _83323_ (_33172_, _33171_, _33169_);
  nor _83324_ (_33173_, _33172_, _33168_);
  nor _83325_ (_33174_, _33173_, _11632_);
  nor _83326_ (_33175_, _33174_, _33167_);
  nor _83327_ (_33176_, _33175_, _32191_);
  nor _83328_ (_33177_, _11630_, _03650_);
  or _83329_ (_33178_, _33177_, _06073_);
  or _83330_ (_33179_, _33178_, _33176_);
  or _83331_ (_33180_, _33179_, _33166_);
  and _83332_ (_33182_, _33180_, _33165_);
  nand _83333_ (_33183_, _33182_, _05966_);
  and _83334_ (_33184_, _04422_, _03311_);
  nor _83335_ (_33185_, _33184_, _03610_);
  and _83336_ (_33186_, _33185_, _33183_);
  or _83337_ (_33187_, _11435_, _11367_);
  or _83338_ (_33188_, _11437_, _11436_);
  and _83339_ (_33189_, _33188_, _11453_);
  nor _83340_ (_33190_, _33188_, _11453_);
  nor _83341_ (_33191_, _33190_, _33189_);
  not _83342_ (_33193_, _33191_);
  or _83343_ (_33194_, _33193_, _11369_);
  nand _83344_ (_33195_, _33194_, _33187_);
  and _83345_ (_33196_, _33195_, _03610_);
  nor _83346_ (_33197_, _33196_, _33186_);
  nand _83347_ (_33198_, _33197_, _11362_);
  nor _83348_ (_33199_, _11362_, _03650_);
  nor _83349_ (_33200_, _33199_, _03715_);
  nand _83350_ (_33201_, _33200_, _33198_);
  and _83351_ (_33202_, _03715_, _03297_);
  nor _83352_ (_33204_, _33202_, _04768_);
  nand _83353_ (_33205_, _33204_, _33201_);
  and _83354_ (_33206_, _03708_, _04768_);
  nor _83355_ (_33207_, _33206_, _03723_);
  nand _83356_ (_33208_, _33207_, _33205_);
  and _83357_ (_33209_, _03723_, _03297_);
  nor _83358_ (_33210_, _33209_, _11660_);
  nand _83359_ (_33211_, _33210_, _33208_);
  nor _83360_ (_33212_, _11659_, _03650_);
  nor _83361_ (_33213_, _33212_, _03729_);
  nand _83362_ (_33215_, _33213_, _33211_);
  and _83363_ (_33216_, _03729_, _03297_);
  nor _83364_ (_33217_, _33216_, _11668_);
  nand _83365_ (_33218_, _33217_, _33215_);
  nor _83366_ (_33219_, _11666_, _03650_);
  nor _83367_ (_33220_, _33219_, _03714_);
  nand _83368_ (_33221_, _33220_, _33218_);
  and _83369_ (_33222_, _03714_, _03297_);
  nor _83370_ (_33223_, _33222_, _11670_);
  nand _83371_ (_33224_, _33223_, _33221_);
  and _83372_ (_33226_, _03708_, _11670_);
  nor _83373_ (_33227_, _33226_, _03508_);
  nand _83374_ (_33228_, _33227_, _33224_);
  and _83375_ (_33229_, _03508_, _03297_);
  nor _83376_ (_33230_, _33229_, _09917_);
  nand _83377_ (_33231_, _33230_, _33228_);
  not _83378_ (_33232_, _23483_);
  and _83379_ (_33233_, _11434_, _09969_);
  nor _83380_ (_33234_, _33193_, _09969_);
  or _83381_ (_33235_, _33234_, _09921_);
  nor _83382_ (_33237_, _33235_, _33233_);
  nor _83383_ (_33238_, _33237_, _33232_);
  nand _83384_ (_33239_, _33238_, _33231_);
  and _83385_ (_33240_, _11434_, _09876_);
  nor _83386_ (_33241_, _33193_, _09876_);
  nor _83387_ (_33242_, _33241_, _33240_);
  nor _83388_ (_33243_, _33242_, _04107_);
  or _83389_ (_33244_, _11435_, _10018_);
  or _83390_ (_33245_, _33193_, _11685_);
  nand _83391_ (_33246_, _33245_, _33244_);
  and _83392_ (_33248_, _33246_, _09919_);
  nor _83393_ (_33249_, _33248_, _33243_);
  nand _83394_ (_33250_, _33249_, _33239_);
  nand _83395_ (_33251_, _33250_, _09856_);
  nor _83396_ (_33252_, _33191_, _10061_);
  and _83397_ (_33253_, _11435_, _10061_);
  or _83398_ (_33254_, _33253_, _09856_);
  nor _83399_ (_33255_, _33254_, _33252_);
  nor _83400_ (_33256_, _33255_, _10025_);
  and _83401_ (_33257_, _33256_, _33251_);
  or _83402_ (_33259_, _33257_, _33155_);
  nand _83403_ (_33260_, _33259_, _06840_);
  and _83404_ (_33261_, _03719_, _03648_);
  nor _83405_ (_33262_, _33261_, _04766_);
  nand _83406_ (_33263_, _33262_, _33260_);
  not _83407_ (_33264_, _32547_);
  nor _83408_ (_33265_, _03708_, _03227_);
  nor _83409_ (_33266_, _33265_, _33264_);
  and _83410_ (_33267_, _33266_, _33263_);
  or _83411_ (_33268_, _33267_, _33154_);
  nand _83412_ (_33270_, _33268_, _11355_);
  nor _83413_ (_33271_, _11355_, _03650_);
  nor _83414_ (_33272_, _33271_, _03753_);
  nand _83415_ (_33273_, _33272_, _33270_);
  and _83416_ (_33274_, _03753_, _03297_);
  nor _83417_ (_33275_, _33274_, _11727_);
  nand _83418_ (_33276_, _33275_, _33273_);
  and _83419_ (_33277_, _03708_, _11727_);
  nor _83420_ (_33278_, _33277_, _03752_);
  nand _83421_ (_33279_, _33278_, _33276_);
  and _83422_ (_33281_, _03752_, _03297_);
  not _83423_ (_33282_, _33281_);
  and _83424_ (_33283_, _33282_, _11350_);
  and _83425_ (_33284_, _33283_, _33279_);
  or _83426_ (_33285_, _33284_, _33153_);
  nand _83427_ (_33286_, _33285_, _08186_);
  nor _83428_ (_33287_, _08186_, _03297_);
  nor _83429_ (_33288_, _33287_, _07912_);
  nand _83430_ (_33289_, _33288_, _33286_);
  nor _83431_ (_33290_, _03248_, _03311_);
  nor _83432_ (_33292_, _33290_, _03505_);
  and _83433_ (_33293_, _33292_, _33289_);
  or _83434_ (_33294_, _33293_, _33152_);
  nand _83435_ (_33295_, _33294_, _05897_);
  and _83436_ (_33296_, _03708_, _03224_);
  nor _83437_ (_33297_, _33296_, _03625_);
  nand _83438_ (_33298_, _33297_, _33295_);
  not _83439_ (_33299_, _11749_);
  and _83440_ (_33300_, _11434_, _03625_);
  nor _83441_ (_33301_, _33300_, _33299_);
  nand _83442_ (_33303_, _33301_, _33298_);
  nor _83443_ (_33304_, _11749_, _03297_);
  nor _83444_ (_33305_, _33304_, _03222_);
  nand _83445_ (_33306_, _33305_, _33303_);
  and _83446_ (_33307_, _11434_, _03222_);
  nor _83447_ (_33308_, _33307_, _11758_);
  nand _83448_ (_33309_, _33308_, _33306_);
  nor _83449_ (_33310_, _11756_, _03650_);
  nor _83450_ (_33311_, _33310_, _03585_);
  and _83451_ (_33312_, _33311_, _33309_);
  and _83452_ (_33314_, _03585_, _03297_);
  or _83453_ (_33315_, _33314_, _03169_);
  or _83454_ (_33316_, _33315_, _33312_);
  and _83455_ (_33317_, _03708_, _03169_);
  nor _83456_ (_33318_, _33317_, _11764_);
  nand _83457_ (_33319_, _33318_, _33316_);
  and _83458_ (_33320_, _33161_, _11764_);
  nor _83459_ (_33321_, _33320_, _06168_);
  nand _83460_ (_33322_, _33321_, _33319_);
  nor _83461_ (_33323_, _05894_, _03297_);
  nor _83462_ (_33325_, _33323_, _03601_);
  nand _83463_ (_33326_, _33325_, _33322_);
  and _83464_ (_33327_, _11434_, _03601_);
  nor _83465_ (_33328_, _33327_, _08363_);
  and _83466_ (_33329_, _33328_, _33326_);
  or _83467_ (_33330_, _33329_, _33151_);
  nand _83468_ (_33331_, _33330_, _11348_);
  nor _83469_ (_33332_, _11348_, _03307_);
  nor _83470_ (_33333_, _33332_, _03584_);
  nand _83471_ (_33334_, _33333_, _33331_);
  and _83472_ (_33336_, _03584_, _03297_);
  nor _83473_ (_33337_, _33336_, _03178_);
  nand _83474_ (_33338_, _33337_, _33334_);
  and _83475_ (_33339_, _03708_, _03178_);
  nor _83476_ (_33340_, _33339_, _11819_);
  nand _83477_ (_33341_, _33340_, _33338_);
  and _83478_ (_33342_, _08786_, _03297_);
  and _83479_ (_33343_, _33161_, _11826_);
  or _83480_ (_33344_, _33343_, _33342_);
  and _83481_ (_33345_, _33344_, _11819_);
  nor _83482_ (_33346_, _33345_, _11824_);
  and _83483_ (_33347_, _33346_, _33341_);
  or _83484_ (_33348_, _33347_, _33150_);
  nand _83485_ (_33349_, _33348_, _11341_);
  nor _83486_ (_33350_, _11341_, _03297_);
  nor _83487_ (_33351_, _33350_, _03600_);
  and _83488_ (_33352_, _33351_, _33349_);
  and _83489_ (_33353_, _11434_, _03600_);
  or _83490_ (_33354_, _33353_, _03780_);
  nor _83491_ (_33355_, _33354_, _33352_);
  and _83492_ (_33358_, _03780_, _03648_);
  or _83493_ (_33359_, _33358_, _33355_);
  nand _83494_ (_33360_, _33359_, _32175_);
  and _83495_ (_33361_, _03708_, _03182_);
  nor _83496_ (_33362_, _33361_, _11841_);
  nand _83497_ (_33363_, _33362_, _33360_);
  or _83498_ (_33364_, _33161_, _11826_);
  or _83499_ (_33365_, _08786_, _03297_);
  and _83500_ (_33366_, _33365_, _11841_);
  and _83501_ (_33367_, _33366_, _33364_);
  nor _83502_ (_33369_, _33367_, _11853_);
  and _83503_ (_33370_, _33369_, _33363_);
  or _83504_ (_33371_, _33370_, _33149_);
  nand _83505_ (_33372_, _33371_, _08430_);
  nor _83506_ (_33373_, _08430_, _03297_);
  nor _83507_ (_33374_, _33373_, _03622_);
  and _83508_ (_33375_, _33374_, _33372_);
  and _83509_ (_33376_, _11434_, _03622_);
  or _83510_ (_33377_, _33376_, _03790_);
  nor _83511_ (_33378_, _33377_, _33375_);
  and _83512_ (_33380_, _03790_, _03648_);
  or _83513_ (_33381_, _33380_, _33378_);
  nand _83514_ (_33382_, _33381_, _32171_);
  and _83515_ (_33383_, _03708_, _03192_);
  nor _83516_ (_33384_, _33383_, _11337_);
  nand _83517_ (_33385_, _33384_, _33382_);
  and _83518_ (_33386_, _03297_, \oc8051_golden_model_1.PSW [7]);
  and _83519_ (_33387_, _33161_, _07871_);
  or _83520_ (_33388_, _33387_, _33386_);
  and _83521_ (_33389_, _33388_, _11337_);
  nor _83522_ (_33391_, _33389_, _11864_);
  and _83523_ (_33392_, _33391_, _33385_);
  or _83524_ (_33393_, _33392_, _33147_);
  nand _83525_ (_33394_, _33393_, _08459_);
  nor _83526_ (_33395_, _08459_, _03297_);
  nor _83527_ (_33396_, _33395_, _03624_);
  and _83528_ (_33397_, _33396_, _33394_);
  and _83529_ (_33398_, _11434_, _03624_);
  or _83530_ (_33399_, _33398_, _03785_);
  nor _83531_ (_33400_, _33399_, _33397_);
  and _83532_ (_33402_, _03785_, _03648_);
  or _83533_ (_33403_, _33402_, _33400_);
  nand _83534_ (_33404_, _33403_, _32168_);
  and _83535_ (_33405_, _03708_, _03201_);
  nor _83536_ (_33406_, _33405_, _11880_);
  nand _83537_ (_33407_, _33406_, _33404_);
  nor _83538_ (_33408_, _33161_, _07871_);
  nor _83539_ (_33409_, _03297_, \oc8051_golden_model_1.PSW [7]);
  nor _83540_ (_33410_, _33409_, _11881_);
  not _83541_ (_33411_, _33410_);
  nor _83542_ (_33413_, _33411_, _33408_);
  nor _83543_ (_33414_, _33413_, _11885_);
  and _83544_ (_33415_, _33414_, _33407_);
  or _83545_ (_33416_, _33415_, _33146_);
  nand _83546_ (_33417_, _33416_, _08507_);
  nor _83547_ (_33418_, _08507_, _03297_);
  nor _83548_ (_33419_, _33418_, _08587_);
  and _83549_ (_33420_, _33419_, _33417_);
  and _83550_ (_33421_, _08587_, _03650_);
  or _83551_ (_33422_, _33421_, _03798_);
  nor _83552_ (_33424_, _33422_, _33420_);
  and _83553_ (_33425_, _08636_, _03798_);
  or _83554_ (_33426_, _33425_, _33424_);
  nand _83555_ (_33427_, _33426_, _06399_);
  and _83556_ (_33428_, _03708_, _03188_);
  nor _83557_ (_33429_, _33428_, _03621_);
  nand _83558_ (_33430_, _33429_, _33427_);
  and _83559_ (_33431_, _33193_, _09854_);
  nor _83560_ (_33432_, _11434_, _09854_);
  or _83561_ (_33433_, _33432_, _11903_);
  or _83562_ (_33435_, _33433_, _33431_);
  and _83563_ (_33436_, _33435_, _11328_);
  and _83564_ (_33437_, _33436_, _33430_);
  or _83565_ (_33438_, _33437_, _33145_);
  nand _83566_ (_33439_, _33438_, _08702_);
  nor _83567_ (_33440_, _08702_, _03297_);
  nor _83568_ (_33441_, _33440_, _08732_);
  and _83569_ (_33442_, _33441_, _33439_);
  and _83570_ (_33443_, _08732_, _03650_);
  or _83571_ (_33444_, _33443_, _03515_);
  nor _83572_ (_33446_, _33444_, _33442_);
  and _83573_ (_33447_, _08636_, _03515_);
  or _83574_ (_33448_, _33447_, _33446_);
  nand _83575_ (_33449_, _33448_, _32165_);
  and _83576_ (_33450_, _03708_, _03203_);
  nor _83577_ (_33451_, _33450_, _03628_);
  nand _83578_ (_33452_, _33451_, _33449_);
  nor _83579_ (_33453_, _33191_, _09854_);
  and _83580_ (_33454_, _11435_, _09854_);
  nor _83581_ (_33455_, _33454_, _33453_);
  and _83582_ (_33457_, _33455_, _03628_);
  nor _83583_ (_33458_, _33457_, _11934_);
  nand _83584_ (_33459_, _33458_, _33452_);
  nor _83585_ (_33460_, _11933_, _03650_);
  nor _83586_ (_33461_, _33460_, _03815_);
  and _83587_ (_33462_, _33461_, _33459_);
  or _83588_ (_33463_, _33462_, _33144_);
  nand _83589_ (_33464_, _33463_, _11940_);
  nor _83590_ (_33465_, _11940_, _03311_);
  nor _83591_ (_33466_, _33465_, _05103_);
  nand _83592_ (_33468_, _33466_, _33464_);
  and _83593_ (_33469_, _05103_, _03708_);
  nor _83594_ (_33470_, _33469_, _03453_);
  nand _83595_ (_33471_, _33470_, _33468_);
  and _83596_ (_33472_, _33455_, _03453_);
  nor _83597_ (_33473_, _33472_, _11958_);
  nand _83598_ (_33474_, _33473_, _33471_);
  nor _83599_ (_33475_, _11957_, _03650_);
  nor _83600_ (_33476_, _33475_, _03447_);
  and _83601_ (_33477_, _33476_, _33474_);
  or _83602_ (_33479_, _33477_, _33143_);
  nand _83603_ (_33480_, _33479_, _11964_);
  nor _83604_ (_33481_, _11964_, _03311_);
  nor _83605_ (_33482_, _33481_, _32154_);
  nand _83606_ (_33483_, _33482_, _33480_);
  and _83607_ (_33484_, _32154_, _03708_);
  nor _83608_ (_33485_, _33484_, _11975_);
  and _83609_ (_33486_, _33485_, _33483_);
  and _83610_ (_33487_, _11975_, _03650_);
  or _83611_ (_33488_, _33487_, _33486_);
  or _83612_ (_33490_, _33488_, _43004_);
  or _83613_ (_33491_, _43000_, \oc8051_golden_model_1.PC [3]);
  and _83614_ (_33492_, _33491_, _41806_);
  and _83615_ (_43672_, _33492_, _33490_);
  and _83616_ (_33493_, _06236_, _05103_);
  and _83617_ (_33494_, _11565_, _03780_);
  and _83618_ (_33495_, _11564_, _08786_);
  and _83619_ (_33496_, _11585_, _11582_);
  nor _83620_ (_33497_, _33496_, _11586_);
  and _83621_ (_33498_, _33497_, _11826_);
  or _83622_ (_33500_, _33498_, _33495_);
  and _83623_ (_33501_, _33500_, _11819_);
  nor _83624_ (_33502_, _32547_, _11564_);
  not _83625_ (_33503_, \oc8051_golden_model_1.PC [4]);
  nor _83626_ (_33504_, _02892_, _33503_);
  and _83627_ (_33505_, _02892_, _33503_);
  nor _83628_ (_33506_, _33505_, _33504_);
  not _83629_ (_33507_, _33506_);
  and _83630_ (_33508_, _33507_, _10025_);
  and _83631_ (_33509_, _11565_, _03714_);
  nor _83632_ (_33511_, _33506_, _11659_);
  and _83633_ (_33512_, _11458_, _11455_);
  nor _83634_ (_33513_, _33512_, _11459_);
  or _83635_ (_33514_, _33513_, _11369_);
  and _83636_ (_33515_, _33514_, _03610_);
  or _83637_ (_33516_, _11430_, _11367_);
  and _83638_ (_33517_, _33516_, _33515_);
  nand _83639_ (_33518_, _33497_, _11624_);
  or _83640_ (_33519_, _11624_, _11565_);
  and _83641_ (_33520_, _33519_, _06073_);
  nand _83642_ (_33522_, _33520_, _33518_);
  not _83643_ (_33523_, _11647_);
  and _83644_ (_33524_, _06236_, _03980_);
  nor _83645_ (_33525_, _33506_, _11642_);
  and _83646_ (_33526_, _11565_, _03979_);
  nor _83647_ (_33527_, _04409_, \oc8051_golden_model_1.PC [4]);
  and _83648_ (_33528_, _33527_, _33169_);
  nor _83649_ (_33529_, _33528_, _33526_);
  nor _83650_ (_33530_, _33529_, _11632_);
  nor _83651_ (_33531_, _33530_, _33525_);
  nor _83652_ (_33533_, _33531_, _03980_);
  nor _83653_ (_33534_, _33533_, _11631_);
  not _83654_ (_33535_, _33534_);
  nor _83655_ (_33536_, _33535_, _33524_);
  nor _83656_ (_33537_, _33507_, _11630_);
  nor _83657_ (_33538_, _33537_, _06073_);
  not _83658_ (_33539_, _33538_);
  nor _83659_ (_33540_, _33539_, _33536_);
  nor _83660_ (_33541_, _33540_, _33523_);
  and _83661_ (_33542_, _33541_, _33522_);
  or _83662_ (_33544_, _33542_, _33517_);
  and _83663_ (_33545_, _33544_, _11362_);
  nor _83664_ (_33546_, _33507_, _11653_);
  or _83665_ (_33547_, _33546_, _03715_);
  or _83666_ (_33548_, _33547_, _33545_);
  and _83667_ (_33549_, _11565_, _03715_);
  nor _83668_ (_33550_, _33549_, _04768_);
  and _83669_ (_33551_, _33550_, _33548_);
  nor _83670_ (_33552_, _06236_, _03230_);
  or _83671_ (_33553_, _33552_, _03723_);
  nor _83672_ (_33555_, _33553_, _33551_);
  and _83673_ (_33556_, _11565_, _03723_);
  or _83674_ (_33557_, _33556_, _33555_);
  and _83675_ (_33558_, _33557_, _11659_);
  or _83676_ (_33559_, _33558_, _33511_);
  nand _83677_ (_33560_, _33559_, _03737_);
  and _83678_ (_33561_, _11565_, _03729_);
  nor _83679_ (_33562_, _33561_, _11668_);
  nand _83680_ (_33563_, _33562_, _33560_);
  nor _83681_ (_33564_, _33507_, _11666_);
  nor _83682_ (_33566_, _33564_, _03714_);
  and _83683_ (_33567_, _33566_, _33563_);
  or _83684_ (_33568_, _33567_, _33509_);
  nand _83685_ (_33569_, _33568_, _03233_);
  and _83686_ (_33570_, _06236_, _11670_);
  nor _83687_ (_33571_, _33570_, _03508_);
  nand _83688_ (_33572_, _33571_, _33569_);
  and _83689_ (_33573_, _11564_, _03508_);
  nor _83690_ (_33574_, _33573_, _09917_);
  nand _83691_ (_33575_, _33574_, _33572_);
  and _83692_ (_33577_, _11430_, _09969_);
  not _83693_ (_33578_, _33513_);
  nor _83694_ (_33579_, _33578_, _09969_);
  or _83695_ (_33580_, _33579_, _09921_);
  nor _83696_ (_33581_, _33580_, _33577_);
  nor _83697_ (_33582_, _33581_, _33232_);
  nand _83698_ (_33583_, _33582_, _33575_);
  and _83699_ (_33584_, _11430_, _09876_);
  nor _83700_ (_33585_, _33578_, _09876_);
  nor _83701_ (_33586_, _33585_, _33584_);
  nor _83702_ (_33588_, _33586_, _04107_);
  and _83703_ (_33589_, _33578_, _10018_);
  or _83704_ (_33590_, _11430_, _10018_);
  nand _83705_ (_33591_, _33590_, _09919_);
  nor _83706_ (_33592_, _33591_, _33589_);
  nor _83707_ (_33593_, _33592_, _33588_);
  nand _83708_ (_33594_, _33593_, _33583_);
  nand _83709_ (_33595_, _33594_, _09856_);
  and _83710_ (_33596_, _11430_, _10061_);
  not _83711_ (_33597_, _10061_);
  and _83712_ (_33599_, _33513_, _33597_);
  or _83713_ (_33600_, _33599_, _33596_);
  and _83714_ (_33601_, _33600_, _03604_);
  nor _83715_ (_33602_, _33601_, _10025_);
  and _83716_ (_33603_, _33602_, _33595_);
  or _83717_ (_33604_, _33603_, _33508_);
  nand _83718_ (_33605_, _33604_, _06840_);
  and _83719_ (_33606_, _11565_, _03719_);
  nor _83720_ (_33607_, _33606_, _04766_);
  nand _83721_ (_33608_, _33607_, _33605_);
  nor _83722_ (_33610_, _06236_, _03227_);
  nor _83723_ (_33611_, _33610_, _33264_);
  and _83724_ (_33612_, _33611_, _33608_);
  or _83725_ (_33613_, _33612_, _33502_);
  nand _83726_ (_33614_, _33613_, _11355_);
  nor _83727_ (_33615_, _33506_, _11355_);
  nor _83728_ (_33616_, _33615_, _03753_);
  and _83729_ (_33617_, _33616_, _33614_);
  and _83730_ (_33618_, _11564_, _03753_);
  or _83731_ (_33619_, _33618_, _33617_);
  and _83732_ (_33621_, _33619_, _03238_);
  nor _83733_ (_33622_, _06236_, _03238_);
  or _83734_ (_33623_, _33622_, _03752_);
  or _83735_ (_33624_, _33623_, _33621_);
  and _83736_ (_33625_, _11565_, _03752_);
  not _83737_ (_33626_, _33625_);
  and _83738_ (_33627_, _33626_, _11350_);
  nand _83739_ (_33628_, _33627_, _33624_);
  nor _83740_ (_33629_, _33507_, _11350_);
  nor _83741_ (_33630_, _33629_, _08187_);
  nand _83742_ (_33632_, _33630_, _33628_);
  nor _83743_ (_33633_, _11564_, _08186_);
  nor _83744_ (_33634_, _33633_, _07912_);
  and _83745_ (_33635_, _33634_, _33632_);
  nor _83746_ (_33636_, _33507_, _03248_);
  or _83747_ (_33637_, _33636_, _03505_);
  nor _83748_ (_33638_, _33637_, _33635_);
  and _83749_ (_33639_, _11565_, _03505_);
  or _83750_ (_33640_, _33639_, _33638_);
  nand _83751_ (_33641_, _33640_, _05897_);
  and _83752_ (_33643_, _06236_, _03224_);
  nor _83753_ (_33644_, _33643_, _03625_);
  nand _83754_ (_33645_, _33644_, _33641_);
  and _83755_ (_33646_, _11430_, _03625_);
  nor _83756_ (_33647_, _33646_, _33299_);
  nand _83757_ (_33648_, _33647_, _33645_);
  nor _83758_ (_33649_, _11749_, _11564_);
  nor _83759_ (_33650_, _33649_, _03222_);
  and _83760_ (_33651_, _33650_, _33648_);
  and _83761_ (_33652_, _11430_, _03222_);
  nor _83762_ (_33654_, _33652_, _33651_);
  nand _83763_ (_33655_, _33654_, _11756_);
  nor _83764_ (_33656_, _33506_, _11756_);
  nor _83765_ (_33657_, _33656_, _03585_);
  and _83766_ (_33658_, _33657_, _33655_);
  and _83767_ (_33659_, _11564_, _03585_);
  or _83768_ (_33660_, _33659_, _03169_);
  or _83769_ (_33661_, _33660_, _33658_);
  and _83770_ (_33662_, _06236_, _03169_);
  nor _83771_ (_33663_, _33662_, _11764_);
  nand _83772_ (_33665_, _33663_, _33661_);
  and _83773_ (_33666_, _33497_, _11764_);
  nor _83774_ (_33667_, _33666_, _06168_);
  nand _83775_ (_33668_, _33667_, _33665_);
  nor _83776_ (_33669_, _11564_, _05894_);
  nor _83777_ (_33670_, _33669_, _03601_);
  nand _83778_ (_33671_, _33670_, _33668_);
  and _83779_ (_33672_, _11430_, _03601_);
  nor _83780_ (_33673_, _33672_, _08363_);
  nand _83781_ (_33674_, _33673_, _33671_);
  and _83782_ (_33676_, _11565_, _08363_);
  nor _83783_ (_33677_, _33676_, _11347_);
  nand _83784_ (_33678_, _33677_, _33674_);
  and _83785_ (_33679_, _11795_, _11792_);
  nor _83786_ (_33680_, _33679_, _11796_);
  and _83787_ (_33681_, _33680_, _11347_);
  nor _83788_ (_33682_, _33681_, _03584_);
  and _83789_ (_33683_, _33682_, _33678_);
  and _83790_ (_33684_, _11565_, _03584_);
  or _83791_ (_33685_, _33684_, _33683_);
  nand _83792_ (_33687_, _33685_, _10736_);
  and _83793_ (_33688_, _06236_, _03178_);
  nor _83794_ (_33689_, _33688_, _11819_);
  and _83795_ (_33690_, _33689_, _33687_);
  or _83796_ (_33691_, _33690_, _33501_);
  nand _83797_ (_33692_, _33691_, _11345_);
  nor _83798_ (_33693_, _33507_, _11345_);
  nor _83799_ (_33694_, _33693_, _11342_);
  nand _83800_ (_33695_, _33694_, _33692_);
  nor _83801_ (_33696_, _11564_, _11341_);
  nor _83802_ (_33698_, _33696_, _03600_);
  nand _83803_ (_33699_, _33698_, _33695_);
  and _83804_ (_33700_, _11430_, _03600_);
  nor _83805_ (_33701_, _33700_, _03780_);
  and _83806_ (_33702_, _33701_, _33699_);
  or _83807_ (_33703_, _33702_, _33494_);
  nand _83808_ (_33704_, _33703_, _32175_);
  and _83809_ (_33705_, _06236_, _03182_);
  nor _83810_ (_33706_, _33705_, _11841_);
  nand _83811_ (_33707_, _33706_, _33704_);
  or _83812_ (_33709_, _11565_, _08786_);
  nand _83813_ (_33710_, _33497_, _08786_);
  and _83814_ (_33711_, _33710_, _33709_);
  or _83815_ (_33712_, _33711_, _11842_);
  nand _83816_ (_33713_, _33712_, _33707_);
  nand _83817_ (_33714_, _33713_, _11851_);
  nor _83818_ (_33715_, _33507_, _11851_);
  nor _83819_ (_33716_, _33715_, _08431_);
  nand _83820_ (_33717_, _33716_, _33714_);
  nor _83821_ (_33718_, _11564_, _08430_);
  nor _83822_ (_33720_, _33718_, _03622_);
  nand _83823_ (_33721_, _33720_, _33717_);
  and _83824_ (_33722_, _11430_, _03622_);
  nor _83825_ (_33723_, _33722_, _03790_);
  and _83826_ (_33724_, _33723_, _33721_);
  and _83827_ (_33725_, _11565_, _03790_);
  or _83828_ (_33726_, _33725_, _33724_);
  nand _83829_ (_33727_, _33726_, _32171_);
  and _83830_ (_33728_, _06236_, _03192_);
  nor _83831_ (_33729_, _33728_, _11337_);
  and _83832_ (_33731_, _33729_, _33727_);
  and _83833_ (_33732_, _11564_, \oc8051_golden_model_1.PSW [7]);
  and _83834_ (_33733_, _33497_, _07871_);
  or _83835_ (_33734_, _33733_, _33732_);
  and _83836_ (_33735_, _33734_, _11337_);
  or _83837_ (_33736_, _33735_, _33731_);
  nand _83838_ (_33737_, _33736_, _11335_);
  nor _83839_ (_33738_, _33507_, _11335_);
  nor _83840_ (_33739_, _33738_, _08460_);
  nand _83841_ (_33740_, _33739_, _33737_);
  nor _83842_ (_33742_, _11564_, _08459_);
  nor _83843_ (_33743_, _33742_, _03624_);
  nand _83844_ (_33744_, _33743_, _33740_);
  and _83845_ (_33745_, _11430_, _03624_);
  nor _83846_ (_33746_, _33745_, _03785_);
  and _83847_ (_33747_, _33746_, _33744_);
  and _83848_ (_33748_, _11565_, _03785_);
  or _83849_ (_33749_, _33748_, _33747_);
  nand _83850_ (_33750_, _33749_, _32168_);
  and _83851_ (_33751_, _06236_, _03201_);
  nor _83852_ (_33753_, _33751_, _11880_);
  nand _83853_ (_33754_, _33753_, _33750_);
  nand _83854_ (_33755_, _11564_, _07871_);
  nand _83855_ (_33756_, _33497_, \oc8051_golden_model_1.PSW [7]);
  and _83856_ (_33757_, _33756_, _33755_);
  or _83857_ (_33758_, _33757_, _11881_);
  nand _83858_ (_33759_, _33758_, _33754_);
  nand _83859_ (_33760_, _33759_, _11330_);
  nor _83860_ (_33761_, _33507_, _11330_);
  nor _83861_ (_33762_, _33761_, _08508_);
  nand _83862_ (_33764_, _33762_, _33760_);
  nor _83863_ (_33765_, _11564_, _08507_);
  nor _83864_ (_33766_, _33765_, _08587_);
  nand _83865_ (_33767_, _33766_, _33764_);
  and _83866_ (_33768_, _33506_, _08587_);
  nor _83867_ (_33769_, _33768_, _03798_);
  and _83868_ (_33770_, _33769_, _33767_);
  nor _83869_ (_33771_, _06730_, _10652_);
  or _83870_ (_33772_, _33771_, _33770_);
  nand _83871_ (_33773_, _33772_, _06399_);
  and _83872_ (_33775_, _06236_, _03188_);
  nor _83873_ (_33776_, _33775_, _03621_);
  and _83874_ (_33777_, _33776_, _33773_);
  nor _83875_ (_33778_, _11431_, _09854_);
  and _83876_ (_33779_, _33513_, _09854_);
  nor _83877_ (_33780_, _33779_, _33778_);
  nor _83878_ (_33781_, _33780_, _11903_);
  or _83879_ (_33782_, _33781_, _33777_);
  nand _83880_ (_33783_, _33782_, _11328_);
  nor _83881_ (_33784_, _33507_, _11328_);
  nor _83882_ (_33785_, _33784_, _08703_);
  nand _83883_ (_33786_, _33785_, _33783_);
  nor _83884_ (_33787_, _11564_, _08702_);
  nor _83885_ (_33788_, _33787_, _08732_);
  nand _83886_ (_33789_, _33788_, _33786_);
  and _83887_ (_33790_, _33506_, _08732_);
  nor _83888_ (_33791_, _33790_, _03515_);
  nand _83889_ (_33792_, _33791_, _33789_);
  nor _83890_ (_33793_, _06730_, _03516_);
  nor _83891_ (_33794_, _33793_, _03203_);
  nand _83892_ (_33796_, _33794_, _33792_);
  nor _83893_ (_33797_, _06236_, _32165_);
  nor _83894_ (_33798_, _33797_, _03628_);
  nand _83895_ (_33799_, _33798_, _33796_);
  and _83896_ (_33800_, _11431_, _09854_);
  nor _83897_ (_33801_, _33513_, _09854_);
  nor _83898_ (_33802_, _33801_, _33800_);
  nor _83899_ (_33803_, _33802_, _03816_);
  nor _83900_ (_33804_, _33803_, _11934_);
  nand _83901_ (_33805_, _33804_, _33799_);
  nor _83902_ (_33807_, _33507_, _11933_);
  nor _83903_ (_33808_, _33807_, _03815_);
  nand _83904_ (_33809_, _33808_, _33805_);
  and _83905_ (_33810_, _11565_, _03815_);
  nor _83906_ (_33811_, _33810_, _32765_);
  nand _83907_ (_33812_, _33811_, _33809_);
  nor _83908_ (_33813_, _33507_, _11940_);
  nor _83909_ (_33814_, _33813_, _05103_);
  and _83910_ (_33815_, _33814_, _33812_);
  or _83911_ (_33816_, _33815_, _33493_);
  nand _83912_ (_33818_, _33816_, _03823_);
  nor _83913_ (_33819_, _33802_, _03823_);
  nor _83914_ (_33820_, _33819_, _11958_);
  nand _83915_ (_33821_, _33820_, _33818_);
  nor _83916_ (_33822_, _33507_, _11957_);
  nor _83917_ (_33823_, _33822_, _03447_);
  nand _83918_ (_33824_, _33823_, _33821_);
  not _83919_ (_33825_, _11964_);
  and _83920_ (_33826_, _11565_, _03447_);
  nor _83921_ (_33827_, _33826_, _33825_);
  nand _83922_ (_33829_, _33827_, _33824_);
  nor _83923_ (_33830_, _33507_, _11964_);
  nor _83924_ (_33831_, _33830_, _32154_);
  nand _83925_ (_33832_, _33831_, _33829_);
  and _83926_ (_33833_, _32154_, _06236_);
  nor _83927_ (_33834_, _33833_, _11975_);
  and _83928_ (_33835_, _33834_, _33832_);
  and _83929_ (_33836_, _33506_, _11975_);
  or _83930_ (_33837_, _33836_, _33835_);
  or _83931_ (_33838_, _33837_, _43004_);
  or _83932_ (_33840_, _43000_, \oc8051_golden_model_1.PC [4]);
  and _83933_ (_33841_, _33840_, _41806_);
  and _83934_ (_43673_, _33841_, _33838_);
  nor _83935_ (_33842_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor _83936_ (_33843_, _11559_, _02905_);
  nor _83937_ (_33844_, _33843_, _33842_);
  and _83938_ (_33845_, _33844_, _11975_);
  and _83939_ (_33846_, _11559_, _03447_);
  nor _83940_ (_33847_, _33844_, _11328_);
  nor _83941_ (_33848_, _33844_, _11330_);
  nor _83942_ (_33850_, _33844_, _11335_);
  nor _83943_ (_33851_, _33844_, _11851_);
  nor _83944_ (_33852_, _33844_, _11345_);
  and _83945_ (_33853_, _11560_, _03584_);
  and _83946_ (_33854_, _11560_, _03505_);
  nor _83947_ (_33855_, _32547_, _11559_);
  and _83948_ (_33856_, _11504_, _11560_);
  or _83949_ (_33857_, _11562_, _11561_);
  and _83950_ (_33858_, _33857_, _11587_);
  nor _83951_ (_33859_, _33857_, _11587_);
  or _83952_ (_33861_, _33859_, _33858_);
  and _83953_ (_33862_, _33861_, _11624_);
  or _83954_ (_33863_, _33862_, _06072_);
  or _83955_ (_33864_, _33863_, _33856_);
  and _83956_ (_33865_, _06267_, _03980_);
  nor _83957_ (_33866_, _33844_, _11643_);
  and _83958_ (_33867_, _11560_, _03979_);
  or _83959_ (_33868_, _04409_, \oc8051_golden_model_1.PC [5]);
  nor _83960_ (_33869_, _33868_, _04729_);
  or _83961_ (_33870_, _33869_, _33867_);
  and _83962_ (_33871_, _33870_, _32816_);
  or _83963_ (_33872_, _33871_, _06073_);
  or _83964_ (_33873_, _33872_, _33866_);
  or _83965_ (_33874_, _33873_, _33865_);
  and _83966_ (_33875_, _33874_, _33864_);
  nand _83967_ (_33876_, _33875_, _05966_);
  not _83968_ (_33877_, _33844_);
  and _83969_ (_33878_, _33877_, _04422_);
  nor _83970_ (_33879_, _33878_, _03610_);
  and _83971_ (_33880_, _33879_, _33876_);
  or _83972_ (_33883_, _11426_, _11367_);
  or _83973_ (_33884_, _11428_, _11427_);
  and _83974_ (_33885_, _33884_, _11460_);
  nor _83975_ (_33886_, _33884_, _11460_);
  or _83976_ (_33887_, _33886_, _33885_);
  or _83977_ (_33888_, _33887_, _11369_);
  nand _83978_ (_33889_, _33888_, _33883_);
  and _83979_ (_33890_, _33889_, _03610_);
  nor _83980_ (_33891_, _33890_, _33880_);
  nand _83981_ (_33892_, _33891_, _11362_);
  nor _83982_ (_33894_, _33844_, _11362_);
  nor _83983_ (_33895_, _33894_, _03715_);
  nand _83984_ (_33896_, _33895_, _33892_);
  and _83985_ (_33897_, _11559_, _03715_);
  nor _83986_ (_33898_, _33897_, _04768_);
  nand _83987_ (_33899_, _33898_, _33896_);
  and _83988_ (_33900_, _06267_, _04768_);
  nor _83989_ (_33901_, _33900_, _03723_);
  nand _83990_ (_33902_, _33901_, _33899_);
  and _83991_ (_33903_, _11559_, _03723_);
  nor _83992_ (_33905_, _33903_, _11660_);
  nand _83993_ (_33906_, _33905_, _33902_);
  nor _83994_ (_33907_, _33844_, _11659_);
  nor _83995_ (_33908_, _33907_, _03729_);
  nand _83996_ (_33909_, _33908_, _33906_);
  and _83997_ (_33910_, _11559_, _03729_);
  nor _83998_ (_33911_, _33910_, _11668_);
  nand _83999_ (_33912_, _33911_, _33909_);
  nor _84000_ (_33913_, _33844_, _11666_);
  nor _84001_ (_33914_, _33913_, _03714_);
  nand _84002_ (_33916_, _33914_, _33912_);
  and _84003_ (_33917_, _11559_, _03714_);
  nor _84004_ (_33918_, _33917_, _11670_);
  nand _84005_ (_33919_, _33918_, _33916_);
  and _84006_ (_33920_, _06267_, _11670_);
  nor _84007_ (_33921_, _33920_, _03508_);
  nand _84008_ (_33922_, _33921_, _33919_);
  and _84009_ (_33923_, _11559_, _03508_);
  nor _84010_ (_33924_, _33923_, _09917_);
  nand _84011_ (_33925_, _33924_, _33922_);
  and _84012_ (_33927_, _11425_, _09969_);
  not _84013_ (_33928_, _33927_);
  nor _84014_ (_33929_, _33887_, _09969_);
  nor _84015_ (_33930_, _33929_, _09921_);
  and _84016_ (_33931_, _33930_, _33928_);
  nor _84017_ (_33932_, _33931_, _33232_);
  nand _84018_ (_33933_, _33932_, _33925_);
  and _84019_ (_33934_, _11425_, _09876_);
  nor _84020_ (_33935_, _33887_, _09876_);
  nor _84021_ (_33936_, _33935_, _33934_);
  nor _84022_ (_33938_, _33936_, _04107_);
  or _84023_ (_33939_, _11426_, _10018_);
  or _84024_ (_33940_, _33887_, _11685_);
  nand _84025_ (_33941_, _33940_, _33939_);
  and _84026_ (_33942_, _33941_, _09919_);
  nor _84027_ (_33943_, _33942_, _33938_);
  nand _84028_ (_33944_, _33943_, _33933_);
  nand _84029_ (_33945_, _33944_, _09856_);
  nand _84030_ (_33946_, _11425_, _10061_);
  or _84031_ (_33947_, _33887_, _10061_);
  and _84032_ (_33949_, _33947_, _33946_);
  or _84033_ (_33950_, _33949_, _09856_);
  and _84034_ (_33951_, _33950_, _33945_);
  or _84035_ (_33952_, _33951_, _10025_);
  nand _84036_ (_33953_, _33844_, _10025_);
  and _84037_ (_33954_, _33953_, _33952_);
  nand _84038_ (_33955_, _33954_, _06840_);
  and _84039_ (_33956_, _11560_, _03719_);
  nor _84040_ (_33957_, _33956_, _04766_);
  nand _84041_ (_33958_, _33957_, _33955_);
  nor _84042_ (_33960_, _06267_, _03227_);
  nor _84043_ (_33961_, _33960_, _33264_);
  and _84044_ (_33962_, _33961_, _33958_);
  or _84045_ (_33963_, _33962_, _33855_);
  nand _84046_ (_33964_, _33963_, _11355_);
  nor _84047_ (_33965_, _33844_, _11355_);
  nor _84048_ (_33966_, _33965_, _03753_);
  nand _84049_ (_33967_, _33966_, _33964_);
  and _84050_ (_33968_, _11559_, _03753_);
  nor _84051_ (_33969_, _33968_, _11727_);
  nand _84052_ (_33971_, _33969_, _33967_);
  and _84053_ (_33972_, _06267_, _11727_);
  nor _84054_ (_33973_, _33972_, _03752_);
  nand _84055_ (_33974_, _33973_, _33971_);
  and _84056_ (_33975_, _11559_, _03752_);
  not _84057_ (_33976_, _33975_);
  and _84058_ (_33977_, _33976_, _11350_);
  and _84059_ (_33978_, _33977_, _33974_);
  nor _84060_ (_33979_, _33844_, _11350_);
  or _84061_ (_33980_, _33979_, _33978_);
  nand _84062_ (_33982_, _33980_, _08186_);
  nor _84063_ (_33983_, _11559_, _08186_);
  nor _84064_ (_33984_, _33983_, _07912_);
  nand _84065_ (_33985_, _33984_, _33982_);
  nor _84066_ (_33986_, _33877_, _03248_);
  nor _84067_ (_33987_, _33986_, _03505_);
  and _84068_ (_33988_, _33987_, _33985_);
  or _84069_ (_33989_, _33988_, _33854_);
  nand _84070_ (_33990_, _33989_, _05897_);
  and _84071_ (_33991_, _06267_, _03224_);
  nor _84072_ (_33993_, _33991_, _03625_);
  nand _84073_ (_33994_, _33993_, _33990_);
  and _84074_ (_33995_, _11425_, _03625_);
  nor _84075_ (_33996_, _33995_, _33299_);
  nand _84076_ (_33997_, _33996_, _33994_);
  nor _84077_ (_33998_, _11749_, _11559_);
  nor _84078_ (_33999_, _33998_, _03222_);
  nand _84079_ (_34000_, _33999_, _33997_);
  and _84080_ (_34001_, _11425_, _03222_);
  nor _84081_ (_34002_, _34001_, _11758_);
  nand _84082_ (_34004_, _34002_, _34000_);
  nor _84083_ (_34005_, _33844_, _11756_);
  nor _84084_ (_34006_, _34005_, _03585_);
  nand _84085_ (_34007_, _34006_, _34004_);
  nor _84086_ (_34008_, _11559_, _03169_);
  or _84087_ (_34009_, _34008_, _11760_);
  nand _84088_ (_34010_, _34009_, _34007_);
  and _84089_ (_34011_, _06267_, _03169_);
  nor _84090_ (_34012_, _34011_, _11764_);
  nand _84091_ (_34013_, _34012_, _34010_);
  nor _84092_ (_34015_, _33861_, _11765_);
  nor _84093_ (_34016_, _34015_, _06168_);
  nand _84094_ (_34017_, _34016_, _34013_);
  nor _84095_ (_34018_, _11559_, _05894_);
  nor _84096_ (_34019_, _34018_, _03601_);
  nand _84097_ (_34020_, _34019_, _34017_);
  and _84098_ (_34021_, _11425_, _03601_);
  nor _84099_ (_34022_, _34021_, _08363_);
  nand _84100_ (_34023_, _34022_, _34020_);
  and _84101_ (_34024_, _11560_, _08363_);
  nor _84102_ (_34026_, _34024_, _11347_);
  nand _84103_ (_34027_, _34026_, _34023_);
  and _84104_ (_34028_, _11797_, _11790_);
  not _84105_ (_34029_, _34028_);
  nor _84106_ (_34030_, _11798_, _11348_);
  and _84107_ (_34031_, _34030_, _34029_);
  nor _84108_ (_34032_, _34031_, _03584_);
  and _84109_ (_34033_, _34032_, _34027_);
  or _84110_ (_34034_, _34033_, _33853_);
  nand _84111_ (_34035_, _34034_, _10736_);
  and _84112_ (_34037_, _06267_, _03178_);
  nor _84113_ (_34038_, _34037_, _11819_);
  nand _84114_ (_34039_, _34038_, _34035_);
  and _84115_ (_34040_, _11559_, _08786_);
  nor _84116_ (_34041_, _33861_, _08786_);
  or _84117_ (_34042_, _34041_, _34040_);
  and _84118_ (_34043_, _34042_, _11819_);
  nor _84119_ (_34044_, _34043_, _11824_);
  and _84120_ (_34045_, _34044_, _34039_);
  or _84121_ (_34046_, _34045_, _33852_);
  nand _84122_ (_34048_, _34046_, _11341_);
  nor _84123_ (_34049_, _11559_, _11341_);
  nor _84124_ (_34050_, _34049_, _03600_);
  and _84125_ (_34051_, _34050_, _34048_);
  and _84126_ (_34052_, _11425_, _03600_);
  or _84127_ (_34053_, _34052_, _03780_);
  nor _84128_ (_34054_, _34053_, _34051_);
  and _84129_ (_34055_, _11560_, _03780_);
  or _84130_ (_34056_, _34055_, _34054_);
  nand _84131_ (_34057_, _34056_, _32175_);
  and _84132_ (_34059_, _06267_, _03182_);
  nor _84133_ (_34060_, _34059_, _11841_);
  nand _84134_ (_34061_, _34060_, _34057_);
  nand _84135_ (_34062_, _33861_, _08786_);
  or _84136_ (_34063_, _11559_, _08786_);
  and _84137_ (_34064_, _34063_, _11841_);
  and _84138_ (_34065_, _34064_, _34062_);
  nor _84139_ (_34066_, _34065_, _11853_);
  and _84140_ (_34067_, _34066_, _34061_);
  or _84141_ (_34068_, _34067_, _33851_);
  nand _84142_ (_34070_, _34068_, _08430_);
  nor _84143_ (_34071_, _11559_, _08430_);
  nor _84144_ (_34072_, _34071_, _03622_);
  and _84145_ (_34073_, _34072_, _34070_);
  and _84146_ (_34074_, _11425_, _03622_);
  or _84147_ (_34075_, _34074_, _03790_);
  nor _84148_ (_34076_, _34075_, _34073_);
  and _84149_ (_34077_, _11560_, _03790_);
  or _84150_ (_34078_, _34077_, _34076_);
  nand _84151_ (_34079_, _34078_, _32171_);
  and _84152_ (_34081_, _06267_, _03192_);
  nor _84153_ (_34082_, _34081_, _11337_);
  nand _84154_ (_34083_, _34082_, _34079_);
  and _84155_ (_34084_, _33861_, _07871_);
  nor _84156_ (_34085_, _11559_, _07871_);
  nor _84157_ (_34086_, _34085_, _11338_);
  not _84158_ (_34087_, _34086_);
  nor _84159_ (_34088_, _34087_, _34084_);
  nor _84160_ (_34089_, _34088_, _11864_);
  and _84161_ (_34090_, _34089_, _34083_);
  or _84162_ (_34092_, _34090_, _33850_);
  nand _84163_ (_34093_, _34092_, _08459_);
  nor _84164_ (_34094_, _11559_, _08459_);
  nor _84165_ (_34095_, _34094_, _03624_);
  and _84166_ (_34096_, _34095_, _34093_);
  and _84167_ (_34097_, _11425_, _03624_);
  or _84168_ (_34098_, _34097_, _03785_);
  nor _84169_ (_34099_, _34098_, _34096_);
  and _84170_ (_34100_, _11560_, _03785_);
  or _84171_ (_34101_, _34100_, _34099_);
  nand _84172_ (_34103_, _34101_, _32168_);
  and _84173_ (_34104_, _06267_, _03201_);
  nor _84174_ (_34105_, _34104_, _11880_);
  nand _84175_ (_34106_, _34105_, _34103_);
  and _84176_ (_34107_, _33861_, \oc8051_golden_model_1.PSW [7]);
  nor _84177_ (_34108_, _11559_, \oc8051_golden_model_1.PSW [7]);
  nor _84178_ (_34109_, _34108_, _11881_);
  not _84179_ (_34110_, _34109_);
  nor _84180_ (_34111_, _34110_, _34107_);
  nor _84181_ (_34112_, _34111_, _11885_);
  and _84182_ (_34114_, _34112_, _34106_);
  or _84183_ (_34115_, _34114_, _33848_);
  nand _84184_ (_34116_, _34115_, _08507_);
  nor _84185_ (_34117_, _11559_, _08507_);
  nor _84186_ (_34118_, _34117_, _08587_);
  nand _84187_ (_34119_, _34118_, _34116_);
  and _84188_ (_34120_, _33844_, _08587_);
  nor _84189_ (_34121_, _34120_, _03798_);
  and _84190_ (_34122_, _34121_, _34119_);
  nor _84191_ (_34123_, _06684_, _10652_);
  or _84192_ (_34125_, _34123_, _34122_);
  nand _84193_ (_34126_, _34125_, _06399_);
  and _84194_ (_34127_, _06267_, _03188_);
  nor _84195_ (_34128_, _34127_, _03621_);
  nand _84196_ (_34129_, _34128_, _34126_);
  and _84197_ (_34130_, _33887_, _09854_);
  nor _84198_ (_34131_, _11425_, _09854_);
  or _84199_ (_34132_, _34131_, _11903_);
  or _84200_ (_34133_, _34132_, _34130_);
  and _84201_ (_34134_, _34133_, _11328_);
  and _84202_ (_34136_, _34134_, _34129_);
  or _84203_ (_34137_, _34136_, _33847_);
  nand _84204_ (_34138_, _34137_, _08702_);
  nor _84205_ (_34139_, _11559_, _08702_);
  nor _84206_ (_34140_, _34139_, _08732_);
  nand _84207_ (_34141_, _34140_, _34138_);
  and _84208_ (_34142_, _33844_, _08732_);
  nor _84209_ (_34143_, _34142_, _03515_);
  and _84210_ (_34144_, _34143_, _34141_);
  nor _84211_ (_34145_, _06684_, _03516_);
  or _84212_ (_34146_, _34145_, _34144_);
  nand _84213_ (_34147_, _34146_, _32165_);
  and _84214_ (_34148_, _06267_, _03203_);
  nor _84215_ (_34149_, _34148_, _03628_);
  nand _84216_ (_34150_, _34149_, _34147_);
  and _84217_ (_34151_, _11425_, _09854_);
  nor _84218_ (_34152_, _33887_, _09854_);
  or _84219_ (_34153_, _34152_, _34151_);
  and _84220_ (_34154_, _34153_, _03628_);
  nor _84221_ (_34155_, _34154_, _11934_);
  nand _84222_ (_34158_, _34155_, _34150_);
  nor _84223_ (_34159_, _33844_, _11933_);
  nor _84224_ (_34160_, _34159_, _03815_);
  nand _84225_ (_34161_, _34160_, _34158_);
  and _84226_ (_34162_, _11559_, _03815_);
  nor _84227_ (_34163_, _34162_, _32765_);
  and _84228_ (_34164_, _34163_, _34161_);
  nor _84229_ (_34165_, _33844_, _11940_);
  or _84230_ (_34166_, _34165_, _34164_);
  nand _84231_ (_34167_, _34166_, _04540_);
  and _84232_ (_34169_, _06267_, _05103_);
  nor _84233_ (_34170_, _34169_, _03453_);
  nand _84234_ (_34171_, _34170_, _34167_);
  and _84235_ (_34172_, _34153_, _03453_);
  nor _84236_ (_34173_, _34172_, _11958_);
  nand _84237_ (_34174_, _34173_, _34171_);
  nor _84238_ (_34175_, _33844_, _11957_);
  nor _84239_ (_34176_, _34175_, _03447_);
  and _84240_ (_34177_, _34176_, _34174_);
  or _84241_ (_34178_, _34177_, _33846_);
  nand _84242_ (_34180_, _34178_, _11964_);
  nor _84243_ (_34181_, _33877_, _11964_);
  nor _84244_ (_34182_, _34181_, _32154_);
  nand _84245_ (_34183_, _34182_, _34180_);
  and _84246_ (_34184_, _32154_, _06267_);
  nor _84247_ (_34185_, _34184_, _11975_);
  and _84248_ (_34186_, _34185_, _34183_);
  or _84249_ (_34187_, _34186_, _33845_);
  or _84250_ (_34188_, _34187_, _43004_);
  or _84251_ (_34189_, _43000_, \oc8051_golden_model_1.PC [5]);
  and _84252_ (_34191_, _34189_, _41806_);
  and _84253_ (_43674_, _34191_, _34188_);
  and _84254_ (_34192_, _06204_, _05103_);
  and _84255_ (_34193_, _06077_, _11315_);
  nor _84256_ (_34194_, _34193_, \oc8051_golden_model_1.PC [6]);
  nor _84257_ (_34195_, _34194_, _11316_);
  not _84258_ (_34196_, _34195_);
  and _84259_ (_34197_, _34196_, _08732_);
  and _84260_ (_34198_, _11418_, _03624_);
  and _84261_ (_34199_, _11418_, _03622_);
  and _84262_ (_34201_, _11418_, _03600_);
  nor _84263_ (_34202_, _34196_, _11350_);
  and _84264_ (_34203_, _11552_, _03714_);
  nor _84265_ (_34204_, _34195_, _11653_);
  and _84266_ (_34205_, _06204_, _03980_);
  nor _84267_ (_34206_, _04729_, \oc8051_golden_model_1.PC [6]);
  or _84268_ (_34207_, _34206_, _04409_);
  and _84269_ (_34208_, _11551_, _04409_);
  nor _84270_ (_34209_, _34208_, _11632_);
  and _84271_ (_34210_, _34209_, _34207_);
  or _84272_ (_34212_, _34195_, _11642_);
  nand _84273_ (_34213_, _34212_, _11630_);
  or _84274_ (_34214_, _34213_, _34210_);
  and _84275_ (_34215_, _34214_, _04763_);
  nor _84276_ (_34216_, _34215_, _34205_);
  nor _84277_ (_34217_, _34196_, _11630_);
  nor _84278_ (_34218_, _34217_, _06073_);
  not _84279_ (_34219_, _34218_);
  nor _84280_ (_34220_, _34219_, _34216_);
  and _84281_ (_34221_, _11589_, _11556_);
  nor _84282_ (_34223_, _34221_, _11590_);
  nand _84283_ (_34224_, _34223_, _11624_);
  or _84284_ (_34225_, _11624_, _11552_);
  and _84285_ (_34226_, _34225_, _06073_);
  and _84286_ (_34227_, _34226_, _34224_);
  or _84287_ (_34228_, _34227_, _34220_);
  nand _84288_ (_34229_, _34228_, _11647_);
  or _84289_ (_34230_, _11418_, _11367_);
  and _84290_ (_34231_, _11462_, _11422_);
  nor _84291_ (_34232_, _34231_, _11463_);
  not _84292_ (_34234_, _34232_);
  or _84293_ (_34235_, _34234_, _11369_);
  and _84294_ (_34236_, _34235_, _03610_);
  nand _84295_ (_34237_, _34236_, _34230_);
  nand _84296_ (_34238_, _34237_, _34229_);
  and _84297_ (_34239_, _34238_, _11362_);
  or _84298_ (_34240_, _34239_, _34204_);
  nand _84299_ (_34241_, _34240_, _04055_);
  and _84300_ (_34242_, _11552_, _03715_);
  nor _84301_ (_34243_, _34242_, _04768_);
  and _84302_ (_34245_, _34243_, _34241_);
  nor _84303_ (_34246_, _06204_, _03230_);
  or _84304_ (_34247_, _34246_, _03723_);
  nor _84305_ (_34248_, _34247_, _34245_);
  and _84306_ (_34249_, _11552_, _03723_);
  or _84307_ (_34250_, _34249_, _34248_);
  and _84308_ (_34251_, _34250_, _11659_);
  nor _84309_ (_34252_, _34195_, _11659_);
  or _84310_ (_34253_, _34252_, _34251_);
  nand _84311_ (_34254_, _34253_, _03737_);
  and _84312_ (_34256_, _11552_, _03729_);
  nor _84313_ (_34257_, _34256_, _11668_);
  nand _84314_ (_34258_, _34257_, _34254_);
  nor _84315_ (_34259_, _34196_, _11666_);
  nor _84316_ (_34260_, _34259_, _03714_);
  and _84317_ (_34261_, _34260_, _34258_);
  or _84318_ (_34262_, _34261_, _34203_);
  nand _84319_ (_34263_, _34262_, _03233_);
  and _84320_ (_34264_, _06204_, _11670_);
  nor _84321_ (_34265_, _34264_, _03508_);
  nand _84322_ (_34267_, _34265_, _34263_);
  and _84323_ (_34268_, _11551_, _03508_);
  nor _84324_ (_34269_, _34268_, _09917_);
  nand _84325_ (_34270_, _34269_, _34267_);
  and _84326_ (_34271_, _11417_, _09969_);
  nor _84327_ (_34272_, _34234_, _09969_);
  or _84328_ (_34273_, _34272_, _09921_);
  nor _84329_ (_34274_, _34273_, _34271_);
  nor _84330_ (_34275_, _34274_, _33232_);
  and _84331_ (_34276_, _34275_, _34270_);
  and _84332_ (_34278_, _34234_, _10018_);
  and _84333_ (_34279_, _11418_, _11685_);
  nor _84334_ (_34280_, _34279_, _34278_);
  and _84335_ (_34281_, _34280_, _32519_);
  nor _84336_ (_34282_, _34281_, _34276_);
  and _84337_ (_34283_, _11418_, _09876_);
  nor _84338_ (_34284_, _34232_, _09876_);
  or _84339_ (_34285_, _34284_, _04107_);
  or _84340_ (_34286_, _34285_, _34283_);
  nand _84341_ (_34287_, _34286_, _34282_);
  nand _84342_ (_34289_, _34287_, _09856_);
  nand _84343_ (_34290_, _11417_, _10061_);
  nand _84344_ (_34291_, _34232_, _33597_);
  and _84345_ (_34292_, _34291_, _34290_);
  or _84346_ (_34293_, _34292_, _09856_);
  and _84347_ (_34294_, _34293_, _34289_);
  or _84348_ (_34295_, _34294_, _10025_);
  nand _84349_ (_34296_, _34195_, _10025_);
  and _84350_ (_34297_, _34296_, _34295_);
  nand _84351_ (_34298_, _34297_, _06840_);
  and _84352_ (_34300_, _11552_, _03719_);
  nor _84353_ (_34301_, _34300_, _04766_);
  nand _84354_ (_34302_, _34301_, _34298_);
  nor _84355_ (_34303_, _06204_, _03227_);
  nor _84356_ (_34304_, _34303_, _33264_);
  and _84357_ (_34305_, _34304_, _34302_);
  nor _84358_ (_34306_, _32547_, _11551_);
  or _84359_ (_34307_, _34306_, _34305_);
  nand _84360_ (_34308_, _34307_, _11355_);
  nor _84361_ (_34309_, _34195_, _11355_);
  nor _84362_ (_34311_, _34309_, _03753_);
  and _84363_ (_34312_, _34311_, _34308_);
  and _84364_ (_34313_, _11551_, _03753_);
  or _84365_ (_34314_, _34313_, _34312_);
  and _84366_ (_34315_, _34314_, _03238_);
  nor _84367_ (_34316_, _06204_, _03238_);
  or _84368_ (_34317_, _34316_, _03752_);
  or _84369_ (_34318_, _34317_, _34315_);
  and _84370_ (_34319_, _11552_, _03752_);
  not _84371_ (_34320_, _34319_);
  and _84372_ (_34322_, _34320_, _11350_);
  and _84373_ (_34323_, _34322_, _34318_);
  or _84374_ (_34324_, _34323_, _34202_);
  and _84375_ (_34325_, _34324_, _08186_);
  nor _84376_ (_34326_, _11552_, _08186_);
  or _84377_ (_34327_, _34326_, _34325_);
  and _84378_ (_34328_, _34327_, _03248_);
  nor _84379_ (_34329_, _34196_, _03248_);
  or _84380_ (_34330_, _34329_, _03505_);
  or _84381_ (_34331_, _34330_, _34328_);
  and _84382_ (_34333_, _11552_, _03505_);
  nor _84383_ (_34334_, _34333_, _03224_);
  nand _84384_ (_34335_, _34334_, _34331_);
  nor _84385_ (_34336_, _06204_, _05897_);
  nor _84386_ (_34337_, _34336_, _03625_);
  nand _84387_ (_34338_, _34337_, _34335_);
  and _84388_ (_34339_, _11418_, _03625_);
  nor _84389_ (_34340_, _34339_, _33299_);
  nand _84390_ (_34341_, _34340_, _34338_);
  nor _84391_ (_34342_, _11749_, _11552_);
  nor _84392_ (_34344_, _34342_, _03222_);
  nand _84393_ (_34345_, _34344_, _34341_);
  and _84394_ (_34346_, _11418_, _03222_);
  nor _84395_ (_34347_, _34346_, _11758_);
  nand _84396_ (_34348_, _34347_, _34345_);
  nor _84397_ (_34349_, _34196_, _11756_);
  nor _84398_ (_34350_, _34349_, _03585_);
  nand _84399_ (_34351_, _34350_, _34348_);
  and _84400_ (_34352_, _11552_, _03585_);
  nor _84401_ (_34353_, _34352_, _03169_);
  and _84402_ (_34355_, _34353_, _34351_);
  nor _84403_ (_34356_, _06204_, _03170_);
  or _84404_ (_34357_, _34356_, _34355_);
  and _84405_ (_34358_, _34357_, _11765_);
  and _84406_ (_34359_, _34223_, _11764_);
  or _84407_ (_34360_, _34359_, _34358_);
  nand _84408_ (_34361_, _34360_, _05894_);
  nor _84409_ (_34362_, _11552_, _05894_);
  nor _84410_ (_34363_, _34362_, _03601_);
  nand _84411_ (_34364_, _34363_, _34361_);
  and _84412_ (_34366_, _11418_, _03601_);
  nor _84413_ (_34367_, _34366_, _08363_);
  nand _84414_ (_34368_, _34367_, _34364_);
  and _84415_ (_34369_, _11551_, _08363_);
  nor _84416_ (_34370_, _34369_, _11347_);
  nand _84417_ (_34371_, _34370_, _34368_);
  and _84418_ (_34372_, _11799_, _11786_);
  nor _84419_ (_34373_, _34372_, _11800_);
  nor _84420_ (_34374_, _34373_, _11348_);
  nor _84421_ (_34375_, _34374_, _03584_);
  nand _84422_ (_34377_, _34375_, _34371_);
  and _84423_ (_34378_, _11551_, _03584_);
  nor _84424_ (_34379_, _34378_, _03178_);
  nand _84425_ (_34380_, _34379_, _34377_);
  and _84426_ (_34381_, _06204_, _03178_);
  nor _84427_ (_34382_, _34381_, _11819_);
  nand _84428_ (_34383_, _34382_, _34380_);
  and _84429_ (_34384_, _11551_, _08786_);
  and _84430_ (_34385_, _34223_, _11826_);
  or _84431_ (_34386_, _34385_, _34384_);
  and _84432_ (_34388_, _34386_, _11819_);
  nor _84433_ (_34389_, _34388_, _11824_);
  nand _84434_ (_34390_, _34389_, _34383_);
  nor _84435_ (_34391_, _34195_, _11345_);
  nor _84436_ (_34392_, _34391_, _11342_);
  nand _84437_ (_34393_, _34392_, _34390_);
  nor _84438_ (_34394_, _11552_, _11341_);
  nor _84439_ (_34395_, _34394_, _03600_);
  and _84440_ (_34396_, _34395_, _34393_);
  or _84441_ (_34397_, _34396_, _34201_);
  nand _84442_ (_34399_, _34397_, _07778_);
  and _84443_ (_34400_, _11552_, _03780_);
  nor _84444_ (_34401_, _34400_, _03182_);
  and _84445_ (_34402_, _34401_, _34399_);
  nor _84446_ (_34403_, _06204_, _32175_);
  or _84447_ (_34404_, _34403_, _34402_);
  nand _84448_ (_34405_, _34404_, _11842_);
  or _84449_ (_34406_, _34223_, _11826_);
  or _84450_ (_34407_, _11551_, _08786_);
  and _84451_ (_34408_, _34407_, _11841_);
  and _84452_ (_34410_, _34408_, _34406_);
  nor _84453_ (_34411_, _34410_, _11853_);
  nand _84454_ (_34412_, _34411_, _34405_);
  nor _84455_ (_34413_, _34195_, _11851_);
  nor _84456_ (_34414_, _34413_, _08431_);
  nand _84457_ (_34415_, _34414_, _34412_);
  nor _84458_ (_34416_, _11552_, _08430_);
  nor _84459_ (_34417_, _34416_, _03622_);
  and _84460_ (_34418_, _34417_, _34415_);
  or _84461_ (_34419_, _34418_, _34199_);
  nand _84462_ (_34421_, _34419_, _06828_);
  and _84463_ (_34422_, _11552_, _03790_);
  nor _84464_ (_34423_, _34422_, _03192_);
  and _84465_ (_34424_, _34423_, _34421_);
  nor _84466_ (_34425_, _06204_, _32171_);
  or _84467_ (_34426_, _34425_, _34424_);
  nand _84468_ (_34427_, _34426_, _11338_);
  and _84469_ (_34428_, _11551_, \oc8051_golden_model_1.PSW [7]);
  and _84470_ (_34429_, _34223_, _07871_);
  or _84471_ (_34430_, _34429_, _34428_);
  and _84472_ (_34432_, _34430_, _11337_);
  nor _84473_ (_34433_, _34432_, _11864_);
  nand _84474_ (_34434_, _34433_, _34427_);
  nor _84475_ (_34435_, _34195_, _11335_);
  nor _84476_ (_34436_, _34435_, _08460_);
  nand _84477_ (_34437_, _34436_, _34434_);
  nor _84478_ (_34438_, _11552_, _08459_);
  nor _84479_ (_34439_, _34438_, _03624_);
  and _84480_ (_34440_, _34439_, _34437_);
  or _84481_ (_34441_, _34440_, _34198_);
  nand _84482_ (_34443_, _34441_, _07793_);
  and _84483_ (_34444_, _11552_, _03785_);
  nor _84484_ (_34445_, _34444_, _03201_);
  and _84485_ (_34446_, _34445_, _34443_);
  nor _84486_ (_34447_, _06204_, _32168_);
  or _84487_ (_34448_, _34447_, _34446_);
  nand _84488_ (_34449_, _34448_, _11881_);
  nor _84489_ (_34450_, _34223_, _07871_);
  nor _84490_ (_34451_, _11551_, \oc8051_golden_model_1.PSW [7]);
  nor _84491_ (_34452_, _34451_, _11881_);
  not _84492_ (_34454_, _34452_);
  nor _84493_ (_34455_, _34454_, _34450_);
  nor _84494_ (_34456_, _34455_, _11885_);
  nand _84495_ (_34457_, _34456_, _34449_);
  nor _84496_ (_34458_, _34195_, _11330_);
  nor _84497_ (_34459_, _34458_, _08508_);
  nand _84498_ (_34460_, _34459_, _34457_);
  nor _84499_ (_34461_, _11552_, _08507_);
  nor _84500_ (_34462_, _34461_, _08587_);
  nand _84501_ (_34463_, _34462_, _34460_);
  and _84502_ (_34465_, _34196_, _08587_);
  nor _84503_ (_34466_, _34465_, _03798_);
  nand _84504_ (_34467_, _34466_, _34463_);
  and _84505_ (_34468_, _06455_, _03798_);
  nor _84506_ (_34469_, _34468_, _03188_);
  nand _84507_ (_34470_, _34469_, _34467_);
  and _84508_ (_34471_, _06204_, _03188_);
  nor _84509_ (_34472_, _34471_, _03621_);
  nand _84510_ (_34473_, _34472_, _34470_);
  nor _84511_ (_34474_, _11417_, _09854_);
  and _84512_ (_34476_, _34234_, _09854_);
  or _84513_ (_34477_, _34476_, _11903_);
  nor _84514_ (_34478_, _34477_, _34474_);
  nor _84515_ (_34479_, _34478_, _11907_);
  nand _84516_ (_34480_, _34479_, _34473_);
  nor _84517_ (_34481_, _34195_, _11328_);
  nor _84518_ (_34482_, _34481_, _08703_);
  nand _84519_ (_34483_, _34482_, _34480_);
  nor _84520_ (_34484_, _11552_, _08702_);
  nor _84521_ (_34485_, _34484_, _08732_);
  and _84522_ (_34487_, _34485_, _34483_);
  or _84523_ (_34488_, _34487_, _34197_);
  nand _84524_ (_34489_, _34488_, _03516_);
  nor _84525_ (_34490_, _06455_, _03516_);
  nor _84526_ (_34491_, _34490_, _03203_);
  nand _84527_ (_34492_, _34491_, _34489_);
  nor _84528_ (_34493_, _06204_, _32165_);
  nor _84529_ (_34494_, _34493_, _03628_);
  and _84530_ (_34495_, _34494_, _34492_);
  nor _84531_ (_34496_, _34232_, _09854_);
  and _84532_ (_34498_, _11418_, _09854_);
  nor _84533_ (_34499_, _34498_, _34496_);
  nor _84534_ (_34500_, _34499_, _03816_);
  or _84535_ (_34501_, _34500_, _34495_);
  and _84536_ (_34502_, _34501_, _11933_);
  nor _84537_ (_34503_, _34195_, _11933_);
  or _84538_ (_34504_, _34503_, _34502_);
  nand _84539_ (_34505_, _34504_, _04246_);
  and _84540_ (_34506_, _11552_, _03815_);
  nor _84541_ (_34507_, _34506_, _32765_);
  nand _84542_ (_34509_, _34507_, _34505_);
  nor _84543_ (_34510_, _34196_, _11940_);
  nor _84544_ (_34511_, _34510_, _05103_);
  and _84545_ (_34512_, _34511_, _34509_);
  or _84546_ (_34513_, _34512_, _34192_);
  nand _84547_ (_34514_, _34513_, _03823_);
  nor _84548_ (_34515_, _34499_, _03823_);
  nor _84549_ (_34516_, _34515_, _11958_);
  nand _84550_ (_34517_, _34516_, _34514_);
  nor _84551_ (_34518_, _34196_, _11957_);
  nor _84552_ (_34520_, _34518_, _03447_);
  nand _84553_ (_34521_, _34520_, _34517_);
  and _84554_ (_34522_, _11552_, _03447_);
  nor _84555_ (_34523_, _34522_, _33825_);
  nand _84556_ (_34524_, _34523_, _34521_);
  nor _84557_ (_34525_, _34196_, _11964_);
  nor _84558_ (_34526_, _34525_, _32154_);
  nand _84559_ (_34527_, _34526_, _34524_);
  and _84560_ (_34528_, _32154_, _06204_);
  nor _84561_ (_34529_, _34528_, _11975_);
  and _84562_ (_34531_, _34529_, _34527_);
  and _84563_ (_34532_, _34195_, _11975_);
  or _84564_ (_34533_, _34532_, _34531_);
  or _84565_ (_34534_, _34533_, _43004_);
  or _84566_ (_34535_, _43000_, \oc8051_golden_model_1.PC [6]);
  and _84567_ (_34536_, _34535_, _41806_);
  and _84568_ (_43675_, _34536_, _34534_);
  and _84569_ (_34537_, _06082_, _03447_);
  and _84570_ (_34538_, _06082_, _03815_);
  nor _84571_ (_34539_, _11316_, \oc8051_golden_model_1.PC [7]);
  nor _84572_ (_34541_, _34539_, _11317_);
  nor _84573_ (_34542_, _34541_, _11328_);
  nor _84574_ (_34543_, _34541_, _11330_);
  nor _84575_ (_34544_, _34541_, _11335_);
  nor _84576_ (_34545_, _34541_, _11851_);
  nor _84577_ (_34546_, _34541_, _11345_);
  and _84578_ (_34547_, _06143_, _03505_);
  nor _84579_ (_34548_, _34541_, _11350_);
  nor _84580_ (_34549_, _32547_, _06082_);
  not _84581_ (_34550_, _34541_);
  and _84582_ (_34552_, _34550_, _10025_);
  and _84583_ (_34553_, _11504_, _06143_);
  or _84584_ (_34554_, _11547_, _11548_);
  and _84585_ (_34555_, _34554_, _11591_);
  nor _84586_ (_34556_, _34554_, _11591_);
  nor _84587_ (_34557_, _34556_, _34555_);
  not _84588_ (_34558_, _34557_);
  and _84589_ (_34559_, _34558_, _11624_);
  or _84590_ (_34560_, _34559_, _06072_);
  or _84591_ (_34561_, _34560_, _34553_);
  and _84592_ (_34563_, _05881_, _03980_);
  nor _84593_ (_34564_, _34541_, _11642_);
  and _84594_ (_34565_, _06143_, _03979_);
  nor _84595_ (_34566_, _04409_, \oc8051_golden_model_1.PC [7]);
  and _84596_ (_34567_, _34566_, _33169_);
  nor _84597_ (_34568_, _34567_, _34565_);
  nor _84598_ (_34569_, _34568_, _11632_);
  nor _84599_ (_34570_, _34569_, _34564_);
  nor _84600_ (_34571_, _34570_, _32191_);
  nor _84601_ (_34572_, _34541_, _11630_);
  or _84602_ (_34574_, _34572_, _06073_);
  or _84603_ (_34575_, _34574_, _34571_);
  or _84604_ (_34576_, _34575_, _34563_);
  and _84605_ (_34577_, _34576_, _34561_);
  nand _84606_ (_34578_, _34577_, _05966_);
  and _84607_ (_34579_, _34550_, _04422_);
  nor _84608_ (_34580_, _34579_, _03610_);
  and _84609_ (_34581_, _34580_, _34578_);
  or _84610_ (_34582_, _11367_, _06749_);
  or _84611_ (_34583_, _11413_, _11414_);
  and _84612_ (_34585_, _34583_, _11464_);
  nor _84613_ (_34586_, _34583_, _11464_);
  nor _84614_ (_34587_, _34586_, _34585_);
  not _84615_ (_34588_, _34587_);
  or _84616_ (_34589_, _34588_, _11369_);
  nand _84617_ (_34590_, _34589_, _34582_);
  and _84618_ (_34591_, _34590_, _03610_);
  nor _84619_ (_34592_, _34591_, _34581_);
  nand _84620_ (_34593_, _34592_, _11362_);
  nor _84621_ (_34594_, _34541_, _11362_);
  nor _84622_ (_34596_, _34594_, _03715_);
  nand _84623_ (_34597_, _34596_, _34593_);
  and _84624_ (_34598_, _06082_, _03715_);
  nor _84625_ (_34599_, _34598_, _04768_);
  nand _84626_ (_34600_, _34599_, _34597_);
  and _84627_ (_34601_, _05881_, _04768_);
  nor _84628_ (_34602_, _34601_, _03723_);
  nand _84629_ (_34603_, _34602_, _34600_);
  and _84630_ (_34604_, _06082_, _03723_);
  nor _84631_ (_34605_, _34604_, _11660_);
  nand _84632_ (_34607_, _34605_, _34603_);
  nor _84633_ (_34608_, _34541_, _11659_);
  nor _84634_ (_34609_, _34608_, _03729_);
  nand _84635_ (_34610_, _34609_, _34607_);
  and _84636_ (_34611_, _06082_, _03729_);
  nor _84637_ (_34612_, _34611_, _11668_);
  nand _84638_ (_34613_, _34612_, _34610_);
  nor _84639_ (_34614_, _34541_, _11666_);
  nor _84640_ (_34615_, _34614_, _03714_);
  nand _84641_ (_34616_, _34615_, _34613_);
  and _84642_ (_34618_, _06082_, _03714_);
  nor _84643_ (_34619_, _34618_, _11670_);
  nand _84644_ (_34620_, _34619_, _34616_);
  and _84645_ (_34621_, _05881_, _11670_);
  nor _84646_ (_34622_, _34621_, _03508_);
  nand _84647_ (_34623_, _34622_, _34620_);
  and _84648_ (_34624_, _06082_, _03508_);
  nor _84649_ (_34625_, _34624_, _09917_);
  nand _84650_ (_34626_, _34625_, _34623_);
  and _84651_ (_34627_, _09969_, _06748_);
  nor _84652_ (_34629_, _34588_, _09969_);
  or _84653_ (_34630_, _34629_, _34627_);
  nor _84654_ (_34631_, _34630_, _09921_);
  nor _84655_ (_34632_, _34631_, _09919_);
  nand _84656_ (_34633_, _34632_, _34626_);
  or _84657_ (_34634_, _10018_, _06749_);
  or _84658_ (_34635_, _34588_, _11685_);
  nand _84659_ (_34636_, _34635_, _34634_);
  nand _84660_ (_34637_, _34636_, _32519_);
  and _84661_ (_34638_, _34637_, _34633_);
  or _84662_ (_34640_, _34638_, _03615_);
  and _84663_ (_34641_, _09876_, _06748_);
  nor _84664_ (_34642_, _34588_, _09876_);
  nor _84665_ (_34643_, _34642_, _34641_);
  or _84666_ (_34644_, _34643_, _04107_);
  and _84667_ (_34645_, _34644_, _34640_);
  or _84668_ (_34646_, _34645_, _03604_);
  and _84669_ (_34647_, _10061_, _06749_);
  nor _84670_ (_34648_, _34587_, _10061_);
  or _84671_ (_34649_, _34648_, _09856_);
  or _84672_ (_34651_, _34649_, _34647_);
  and _84673_ (_34652_, _34651_, _11358_);
  and _84674_ (_34653_, _34652_, _34646_);
  or _84675_ (_34654_, _34653_, _34552_);
  nand _84676_ (_34655_, _34654_, _06840_);
  and _84677_ (_34656_, _06143_, _03719_);
  nor _84678_ (_34657_, _34656_, _04766_);
  nand _84679_ (_34658_, _34657_, _34655_);
  nor _84680_ (_34659_, _05881_, _03227_);
  nor _84681_ (_34660_, _34659_, _33264_);
  and _84682_ (_34662_, _34660_, _34658_);
  or _84683_ (_34663_, _34662_, _34549_);
  nand _84684_ (_34664_, _34663_, _11355_);
  nor _84685_ (_34665_, _34541_, _11355_);
  nor _84686_ (_34666_, _34665_, _03753_);
  nand _84687_ (_34667_, _34666_, _34664_);
  and _84688_ (_34668_, _06082_, _03753_);
  nor _84689_ (_34669_, _34668_, _11727_);
  nand _84690_ (_34670_, _34669_, _34667_);
  and _84691_ (_34671_, _05881_, _11727_);
  nor _84692_ (_34673_, _34671_, _03752_);
  nand _84693_ (_34674_, _34673_, _34670_);
  and _84694_ (_34675_, _06082_, _03752_);
  not _84695_ (_34676_, _34675_);
  and _84696_ (_34677_, _34676_, _11350_);
  and _84697_ (_34678_, _34677_, _34674_);
  or _84698_ (_34679_, _34678_, _34548_);
  nand _84699_ (_34680_, _34679_, _08186_);
  nor _84700_ (_34681_, _08186_, _06082_);
  nor _84701_ (_34682_, _34681_, _07912_);
  nand _84702_ (_34684_, _34682_, _34680_);
  nor _84703_ (_34685_, _34550_, _03248_);
  nor _84704_ (_34686_, _34685_, _03505_);
  and _84705_ (_34687_, _34686_, _34684_);
  or _84706_ (_34688_, _34687_, _34547_);
  nand _84707_ (_34689_, _34688_, _05897_);
  and _84708_ (_34690_, _05881_, _03224_);
  nor _84709_ (_34691_, _34690_, _03625_);
  nand _84710_ (_34692_, _34691_, _34689_);
  and _84711_ (_34693_, _06748_, _03625_);
  nor _84712_ (_34695_, _34693_, _33299_);
  nand _84713_ (_34696_, _34695_, _34692_);
  nor _84714_ (_34697_, _11749_, _06082_);
  nor _84715_ (_34698_, _34697_, _03222_);
  nand _84716_ (_34699_, _34698_, _34696_);
  and _84717_ (_34700_, _06748_, _03222_);
  nor _84718_ (_34701_, _34700_, _11758_);
  nand _84719_ (_34702_, _34701_, _34699_);
  nor _84720_ (_34703_, _34541_, _11756_);
  nor _84721_ (_34704_, _34703_, _03585_);
  nand _84722_ (_34706_, _34704_, _34702_);
  nor _84723_ (_34707_, _06082_, _03169_);
  or _84724_ (_34708_, _34707_, _11760_);
  nand _84725_ (_34709_, _34708_, _34706_);
  and _84726_ (_34710_, _05881_, _03169_);
  nor _84727_ (_34711_, _34710_, _11764_);
  nand _84728_ (_34712_, _34711_, _34709_);
  and _84729_ (_34713_, _34557_, _11764_);
  nor _84730_ (_34714_, _34713_, _06168_);
  nand _84731_ (_34715_, _34714_, _34712_);
  nor _84732_ (_34717_, _06082_, _05894_);
  nor _84733_ (_34718_, _34717_, _03601_);
  nand _84734_ (_34719_, _34718_, _34715_);
  and _84735_ (_34720_, _06748_, _03601_);
  nor _84736_ (_34721_, _34720_, _08363_);
  nand _84737_ (_34722_, _34721_, _34719_);
  and _84738_ (_34723_, _08363_, _06143_);
  nor _84739_ (_34724_, _34723_, _11347_);
  nand _84740_ (_34725_, _34724_, _34722_);
  or _84741_ (_34726_, _11781_, _11782_);
  and _84742_ (_34728_, _34726_, _11801_);
  nor _84743_ (_34729_, _34726_, _11801_);
  or _84744_ (_34730_, _34729_, _34728_);
  nor _84745_ (_34731_, _34730_, _11348_);
  nor _84746_ (_34732_, _34731_, _03584_);
  and _84747_ (_34733_, _34732_, _34725_);
  and _84748_ (_34734_, _06143_, _03584_);
  or _84749_ (_34735_, _34734_, _34733_);
  nand _84750_ (_34736_, _34735_, _10736_);
  and _84751_ (_34737_, _05881_, _03178_);
  nor _84752_ (_34739_, _34737_, _11819_);
  nand _84753_ (_34740_, _34739_, _34736_);
  and _84754_ (_34741_, _08786_, _06082_);
  and _84755_ (_34742_, _34557_, _11826_);
  or _84756_ (_34743_, _34742_, _34741_);
  and _84757_ (_34744_, _34743_, _11819_);
  nor _84758_ (_34745_, _34744_, _11824_);
  and _84759_ (_34746_, _34745_, _34740_);
  or _84760_ (_34747_, _34746_, _34546_);
  nand _84761_ (_34748_, _34747_, _11341_);
  nor _84762_ (_34750_, _11341_, _06082_);
  nor _84763_ (_34751_, _34750_, _03600_);
  and _84764_ (_34752_, _34751_, _34748_);
  and _84765_ (_34753_, _06748_, _03600_);
  or _84766_ (_34754_, _34753_, _03780_);
  nor _84767_ (_34755_, _34754_, _34752_);
  and _84768_ (_34756_, _06143_, _03780_);
  or _84769_ (_34757_, _34756_, _34755_);
  nand _84770_ (_34758_, _34757_, _32175_);
  and _84771_ (_34759_, _05881_, _03182_);
  nor _84772_ (_34761_, _34759_, _11841_);
  nand _84773_ (_34762_, _34761_, _34758_);
  or _84774_ (_34763_, _34557_, _11826_);
  or _84775_ (_34764_, _08786_, _06082_);
  and _84776_ (_34765_, _34764_, _11841_);
  and _84777_ (_34766_, _34765_, _34763_);
  nor _84778_ (_34767_, _34766_, _11853_);
  and _84779_ (_34768_, _34767_, _34762_);
  or _84780_ (_34769_, _34768_, _34545_);
  nand _84781_ (_34770_, _34769_, _08430_);
  nor _84782_ (_34771_, _08430_, _06082_);
  nor _84783_ (_34772_, _34771_, _03622_);
  and _84784_ (_34773_, _34772_, _34770_);
  and _84785_ (_34774_, _06748_, _03622_);
  or _84786_ (_34775_, _34774_, _03790_);
  nor _84787_ (_34776_, _34775_, _34773_);
  and _84788_ (_34777_, _06143_, _03790_);
  or _84789_ (_34778_, _34777_, _34776_);
  nand _84790_ (_34779_, _34778_, _32171_);
  and _84791_ (_34780_, _05881_, _03192_);
  nor _84792_ (_34783_, _34780_, _11337_);
  nand _84793_ (_34784_, _34783_, _34779_);
  and _84794_ (_34785_, _06082_, \oc8051_golden_model_1.PSW [7]);
  and _84795_ (_34786_, _34557_, _07871_);
  or _84796_ (_34787_, _34786_, _34785_);
  and _84797_ (_34788_, _34787_, _11337_);
  nor _84798_ (_34789_, _34788_, _11864_);
  and _84799_ (_34790_, _34789_, _34784_);
  or _84800_ (_34791_, _34790_, _34544_);
  nand _84801_ (_34792_, _34791_, _08459_);
  nor _84802_ (_34794_, _08459_, _06082_);
  nor _84803_ (_34795_, _34794_, _03624_);
  and _84804_ (_34796_, _34795_, _34792_);
  and _84805_ (_34797_, _06748_, _03624_);
  or _84806_ (_34798_, _34797_, _03785_);
  nor _84807_ (_34799_, _34798_, _34796_);
  and _84808_ (_34800_, _06143_, _03785_);
  or _84809_ (_34801_, _34800_, _34799_);
  nand _84810_ (_34802_, _34801_, _32168_);
  and _84811_ (_34803_, _05881_, _03201_);
  nor _84812_ (_34805_, _34803_, _11880_);
  nand _84813_ (_34806_, _34805_, _34802_);
  nor _84814_ (_34807_, _34557_, _07871_);
  nor _84815_ (_34808_, _06082_, \oc8051_golden_model_1.PSW [7]);
  nor _84816_ (_34809_, _34808_, _11881_);
  not _84817_ (_34810_, _34809_);
  nor _84818_ (_34811_, _34810_, _34807_);
  nor _84819_ (_34812_, _34811_, _11885_);
  and _84820_ (_34813_, _34812_, _34806_);
  or _84821_ (_34814_, _34813_, _34543_);
  nand _84822_ (_34816_, _34814_, _08507_);
  nor _84823_ (_34817_, _08507_, _06082_);
  nor _84824_ (_34818_, _34817_, _08587_);
  nand _84825_ (_34819_, _34818_, _34816_);
  and _84826_ (_34820_, _34541_, _08587_);
  nor _84827_ (_34821_, _34820_, _03798_);
  and _84828_ (_34822_, _34821_, _34819_);
  nor _84829_ (_34823_, _06069_, _10652_);
  or _84830_ (_34824_, _34823_, _34822_);
  nand _84831_ (_34825_, _34824_, _06399_);
  and _84832_ (_34827_, _05881_, _03188_);
  nor _84833_ (_34828_, _34827_, _03621_);
  nand _84834_ (_34829_, _34828_, _34825_);
  and _84835_ (_34830_, _34588_, _09854_);
  nor _84836_ (_34831_, _09854_, _06748_);
  or _84837_ (_34832_, _34831_, _11903_);
  or _84838_ (_34833_, _34832_, _34830_);
  and _84839_ (_34834_, _34833_, _11328_);
  and _84840_ (_34835_, _34834_, _34829_);
  or _84841_ (_34836_, _34835_, _34542_);
  nand _84842_ (_34838_, _34836_, _08702_);
  nor _84843_ (_34839_, _08702_, _06082_);
  nor _84844_ (_34840_, _34839_, _08732_);
  nand _84845_ (_34841_, _34840_, _34838_);
  and _84846_ (_34842_, _34541_, _08732_);
  nor _84847_ (_34843_, _34842_, _03515_);
  and _84848_ (_34844_, _34843_, _34841_);
  nor _84849_ (_34845_, _06069_, _03516_);
  or _84850_ (_34846_, _34845_, _34844_);
  nand _84851_ (_34847_, _34846_, _32165_);
  and _84852_ (_34849_, _05881_, _03203_);
  nor _84853_ (_34850_, _34849_, _03628_);
  nand _84854_ (_34851_, _34850_, _34847_);
  and _84855_ (_34852_, _09854_, _06749_);
  nor _84856_ (_34853_, _34587_, _09854_);
  nor _84857_ (_34854_, _34853_, _34852_);
  and _84858_ (_34855_, _34854_, _03628_);
  nor _84859_ (_34856_, _34855_, _11934_);
  nand _84860_ (_34857_, _34856_, _34851_);
  nor _84861_ (_34858_, _34541_, _11933_);
  nor _84862_ (_34860_, _34858_, _03815_);
  and _84863_ (_34861_, _34860_, _34857_);
  or _84864_ (_34862_, _34861_, _34538_);
  nand _84865_ (_34863_, _34862_, _11940_);
  nor _84866_ (_34864_, _34550_, _11940_);
  nor _84867_ (_34865_, _34864_, _05103_);
  nand _84868_ (_34866_, _34865_, _34863_);
  and _84869_ (_34867_, _05881_, _05103_);
  nor _84870_ (_34868_, _34867_, _03453_);
  nand _84871_ (_34869_, _34868_, _34866_);
  and _84872_ (_34871_, _34854_, _03453_);
  nor _84873_ (_34872_, _34871_, _11958_);
  nand _84874_ (_34873_, _34872_, _34869_);
  nor _84875_ (_34874_, _34541_, _11957_);
  nor _84876_ (_34875_, _34874_, _03447_);
  and _84877_ (_34876_, _34875_, _34873_);
  or _84878_ (_34877_, _34876_, _34537_);
  nand _84879_ (_34878_, _34877_, _11964_);
  nor _84880_ (_34879_, _34550_, _11964_);
  nor _84881_ (_34880_, _34879_, _32154_);
  nand _84882_ (_34882_, _34880_, _34878_);
  and _84883_ (_34883_, _32154_, _05881_);
  nor _84884_ (_34884_, _34883_, _11975_);
  and _84885_ (_34885_, _34884_, _34882_);
  and _84886_ (_34886_, _34541_, _11975_);
  or _84887_ (_34887_, _34886_, _34885_);
  or _84888_ (_34888_, _34887_, _43004_);
  or _84889_ (_34889_, _43000_, \oc8051_golden_model_1.PC [7]);
  and _84890_ (_34890_, _34889_, _41806_);
  and _84891_ (_43676_, _34890_, _34888_);
  nor _84892_ (_34892_, _04048_, _11968_);
  nor _84893_ (_34893_, _04048_, _11944_);
  and _84894_ (_34894_, _11469_, _03624_);
  nor _84895_ (_34895_, _11337_, _03192_);
  nor _84896_ (_34896_, _11595_, _05894_);
  and _84897_ (_34897_, _11595_, _03585_);
  or _84898_ (_34898_, _11468_, _10018_);
  nor _84899_ (_34899_, _11472_, _11466_);
  nor _84900_ (_34900_, _34899_, _11473_);
  or _84901_ (_34901_, _34900_, _11685_);
  nand _84902_ (_34903_, _34901_, _34898_);
  nand _84903_ (_34904_, _34903_, _09919_);
  and _84904_ (_34905_, _11468_, _09969_);
  not _84905_ (_34906_, _34900_);
  nor _84906_ (_34907_, _34906_, _09969_);
  or _84907_ (_34908_, _34907_, _34905_);
  nor _84908_ (_34909_, _34908_, _09921_);
  and _84909_ (_34910_, _11595_, _03714_);
  nor _84910_ (_34911_, _03723_, _04768_);
  and _84911_ (_34912_, _11595_, _03715_);
  or _84912_ (_34914_, _11468_, _11367_);
  or _84913_ (_34915_, _34900_, _11369_);
  and _84914_ (_34916_, _34915_, _34914_);
  or _84915_ (_34917_, _34916_, _04081_);
  and _84916_ (_34918_, _11504_, _11595_);
  nor _84917_ (_34919_, _11599_, _11593_);
  nor _84918_ (_34920_, _34919_, _11600_);
  and _84919_ (_34921_, _34920_, _11624_);
  nor _84920_ (_34922_, _34921_, _34918_);
  nand _84921_ (_34923_, _34922_, _06073_);
  nand _84922_ (_34925_, _11596_, _03979_);
  or _84923_ (_34926_, _04409_, \oc8051_golden_model_1.PC [8]);
  or _84924_ (_34927_, _34926_, _04729_);
  and _84925_ (_34928_, _34927_, _34925_);
  or _84926_ (_34929_, _34928_, _11632_);
  nor _84927_ (_34930_, _11317_, \oc8051_golden_model_1.PC [8]);
  nor _84928_ (_34931_, _34930_, _11318_);
  or _84929_ (_34932_, _34931_, _11642_);
  and _84930_ (_34933_, _34932_, _34929_);
  nor _84931_ (_34934_, _34933_, _32191_);
  nor _84932_ (_34936_, _34931_, _11630_);
  nor _84933_ (_34937_, _34936_, _34934_);
  nor _84934_ (_34938_, _34937_, _06073_);
  nor _84935_ (_34939_, _34938_, _04422_);
  and _84936_ (_34940_, _34939_, _34923_);
  and _84937_ (_34941_, _34931_, _04422_);
  or _84938_ (_34942_, _34941_, _03610_);
  or _84939_ (_34943_, _34942_, _34940_);
  nand _84940_ (_34944_, _34943_, _34917_);
  nand _84941_ (_34945_, _34944_, _11362_);
  nor _84942_ (_34947_, _34931_, _11362_);
  nor _84943_ (_34948_, _34947_, _03715_);
  and _84944_ (_34949_, _34948_, _34945_);
  or _84945_ (_34950_, _34949_, _34912_);
  nand _84946_ (_34951_, _34950_, _34911_);
  and _84947_ (_34952_, _11595_, _03723_);
  nor _84948_ (_34953_, _34952_, _11660_);
  nand _84949_ (_34954_, _34953_, _34951_);
  nor _84950_ (_34955_, _34931_, _11659_);
  nor _84951_ (_34956_, _34955_, _03729_);
  nand _84952_ (_34958_, _34956_, _34954_);
  and _84953_ (_34959_, _11595_, _03729_);
  nor _84954_ (_34960_, _34959_, _11668_);
  nand _84955_ (_34961_, _34960_, _34958_);
  nor _84956_ (_34962_, _34931_, _11666_);
  nor _84957_ (_34963_, _34962_, _03714_);
  and _84958_ (_34964_, _34963_, _34961_);
  or _84959_ (_34965_, _34964_, _34910_);
  nand _84960_ (_34966_, _34965_, _11671_);
  and _84961_ (_34967_, _11595_, _03508_);
  nor _84962_ (_34969_, _34967_, _09917_);
  and _84963_ (_34970_, _34969_, _34966_);
  or _84964_ (_34971_, _34970_, _34909_);
  nand _84965_ (_34972_, _34971_, _09920_);
  nand _84966_ (_34973_, _34972_, _34904_);
  or _84967_ (_34974_, _34973_, _03615_);
  nor _84968_ (_34975_, _34906_, _09876_);
  and _84969_ (_34976_, _11468_, _09876_);
  nor _84970_ (_34977_, _34976_, _34975_);
  or _84971_ (_34978_, _34977_, _04107_);
  and _84972_ (_34980_, _34978_, _34974_);
  or _84973_ (_34981_, _34980_, _03604_);
  and _84974_ (_34982_, _11468_, _10061_);
  and _84975_ (_34983_, _34900_, _33597_);
  or _84976_ (_34984_, _34983_, _34982_);
  and _84977_ (_34985_, _34984_, _03604_);
  nor _84978_ (_34986_, _34985_, _10025_);
  nand _84979_ (_34987_, _34986_, _34981_);
  not _84980_ (_34988_, _34931_);
  and _84981_ (_34989_, _34988_, _10025_);
  nor _84982_ (_34991_, _34989_, _03719_);
  nand _84983_ (_34992_, _34991_, _34987_);
  and _84984_ (_34993_, _11595_, _03719_);
  nor _84985_ (_34994_, _34993_, _04766_);
  nand _84986_ (_34995_, _34994_, _34992_);
  nand _84987_ (_34996_, _34995_, _32547_);
  nor _84988_ (_34997_, _32547_, _11596_);
  nor _84989_ (_34998_, _34997_, _11356_);
  nand _84990_ (_34999_, _34998_, _34996_);
  nor _84991_ (_35000_, _34931_, _11355_);
  nor _84992_ (_35002_, _35000_, _03753_);
  nand _84993_ (_35003_, _35002_, _34999_);
  and _84994_ (_35004_, _11595_, _03753_);
  nor _84995_ (_35005_, _35004_, _11727_);
  nand _84996_ (_35006_, _35005_, _35003_);
  nand _84997_ (_35007_, _35006_, _09668_);
  and _84998_ (_35008_, _11595_, _03752_);
  not _84999_ (_35009_, _35008_);
  and _85000_ (_35010_, _35009_, _11350_);
  nand _85001_ (_35011_, _35010_, _35007_);
  nor _85002_ (_35013_, _34931_, _11350_);
  nor _85003_ (_35014_, _35013_, _08187_);
  and _85004_ (_35015_, _35014_, _35011_);
  nor _85005_ (_35016_, _11596_, _08186_);
  or _85006_ (_35017_, _35016_, _07912_);
  nor _85007_ (_35018_, _35017_, _35015_);
  nor _85008_ (_35019_, _34931_, _03248_);
  or _85009_ (_35020_, _35019_, _35018_);
  nand _85010_ (_35021_, _35020_, _03710_);
  and _85011_ (_35022_, _11596_, _03505_);
  nor _85012_ (_35024_, _35022_, _23690_);
  and _85013_ (_35025_, _35024_, _35021_);
  and _85014_ (_35026_, _11468_, _03625_);
  nor _85015_ (_35027_, _35026_, _35025_);
  nand _85016_ (_35028_, _35027_, _11749_);
  nor _85017_ (_35029_, _11749_, _11595_);
  nor _85018_ (_35030_, _35029_, _03222_);
  nand _85019_ (_35031_, _35030_, _35028_);
  and _85020_ (_35032_, _11468_, _03222_);
  nor _85021_ (_35033_, _35032_, _11758_);
  nand _85022_ (_35035_, _35033_, _35031_);
  nor _85023_ (_35036_, _34931_, _11756_);
  nor _85024_ (_35037_, _35036_, _03585_);
  and _85025_ (_35038_, _35037_, _35035_);
  or _85026_ (_35039_, _35038_, _34897_);
  nor _85027_ (_35040_, _11764_, _03169_);
  nand _85028_ (_35041_, _35040_, _35039_);
  and _85029_ (_35042_, _34920_, _11764_);
  nor _85030_ (_35043_, _35042_, _06168_);
  and _85031_ (_35044_, _35043_, _35041_);
  or _85032_ (_35046_, _35044_, _34896_);
  nand _85033_ (_35047_, _35046_, _05886_);
  and _85034_ (_35048_, _11469_, _03601_);
  nor _85035_ (_35049_, _35048_, _08363_);
  nand _85036_ (_35050_, _35049_, _35047_);
  and _85037_ (_35051_, _11595_, _08363_);
  nor _85038_ (_35052_, _35051_, _11347_);
  nand _85039_ (_35053_, _35052_, _35050_);
  nor _85040_ (_35054_, _11803_, \oc8051_golden_model_1.DPH [0]);
  nor _85041_ (_35055_, _35054_, _11804_);
  nor _85042_ (_35057_, _35055_, _11348_);
  nor _85043_ (_35058_, _35057_, _03584_);
  nand _85044_ (_35059_, _35058_, _35053_);
  and _85045_ (_35060_, _11595_, _03584_);
  nor _85046_ (_35061_, _35060_, _03178_);
  nand _85047_ (_35062_, _35061_, _35059_);
  nand _85048_ (_35063_, _35062_, _11820_);
  and _85049_ (_35064_, _11595_, _08786_);
  and _85050_ (_35065_, _34920_, _11826_);
  or _85051_ (_35066_, _35065_, _35064_);
  and _85052_ (_35068_, _35066_, _11819_);
  nor _85053_ (_35069_, _35068_, _11824_);
  nand _85054_ (_35070_, _35069_, _35063_);
  nor _85055_ (_35071_, _34931_, _11345_);
  nor _85056_ (_35072_, _35071_, _11342_);
  nand _85057_ (_35073_, _35072_, _35070_);
  nor _85058_ (_35074_, _11596_, _11341_);
  nor _85059_ (_35075_, _35074_, _03600_);
  nand _85060_ (_35076_, _35075_, _35073_);
  and _85061_ (_35077_, _11469_, _03600_);
  nor _85062_ (_35079_, _35077_, _03780_);
  nand _85063_ (_35080_, _35079_, _35076_);
  and _85064_ (_35081_, _11595_, _03780_);
  nor _85065_ (_35082_, _35081_, _03182_);
  nand _85066_ (_35083_, _35082_, _35080_);
  nand _85067_ (_35084_, _35083_, _11842_);
  or _85068_ (_35085_, _34920_, _11826_);
  or _85069_ (_35086_, _11595_, _08786_);
  and _85070_ (_35087_, _35086_, _11841_);
  and _85071_ (_35088_, _35087_, _35085_);
  nor _85072_ (_35090_, _35088_, _11853_);
  nand _85073_ (_35091_, _35090_, _35084_);
  nor _85074_ (_35092_, _34931_, _11851_);
  nor _85075_ (_35093_, _35092_, _08431_);
  and _85076_ (_35094_, _35093_, _35091_);
  nor _85077_ (_35095_, _11596_, _08430_);
  or _85078_ (_35096_, _35095_, _03622_);
  or _85079_ (_35097_, _35096_, _35094_);
  and _85080_ (_35098_, _11469_, _03622_);
  nor _85081_ (_35099_, _35098_, _03790_);
  and _85082_ (_35101_, _35099_, _35097_);
  and _85083_ (_35102_, _11595_, _03790_);
  or _85084_ (_35103_, _35102_, _35101_);
  nand _85085_ (_35104_, _35103_, _34895_);
  and _85086_ (_35105_, _11595_, \oc8051_golden_model_1.PSW [7]);
  and _85087_ (_35106_, _34920_, _07871_);
  or _85088_ (_35107_, _35106_, _35105_);
  and _85089_ (_35108_, _35107_, _11337_);
  nor _85090_ (_35109_, _35108_, _11864_);
  nand _85091_ (_35110_, _35109_, _35104_);
  nor _85092_ (_35112_, _34931_, _11335_);
  nor _85093_ (_35113_, _35112_, _08460_);
  nand _85094_ (_35114_, _35113_, _35110_);
  nor _85095_ (_35115_, _11596_, _08459_);
  nor _85096_ (_35116_, _35115_, _03624_);
  and _85097_ (_35117_, _35116_, _35114_);
  or _85098_ (_35118_, _35117_, _34894_);
  nand _85099_ (_35119_, _35118_, _07793_);
  nor _85100_ (_35120_, _11880_, _03201_);
  and _85101_ (_35121_, _11596_, _03785_);
  not _85102_ (_35123_, _35121_);
  and _85103_ (_35124_, _35123_, _35120_);
  nand _85104_ (_35125_, _35124_, _35119_);
  nor _85105_ (_35126_, _34920_, _07871_);
  nor _85106_ (_35127_, _11595_, \oc8051_golden_model_1.PSW [7]);
  nor _85107_ (_35128_, _35127_, _11881_);
  not _85108_ (_35129_, _35128_);
  nor _85109_ (_35130_, _35129_, _35126_);
  nor _85110_ (_35131_, _35130_, _11885_);
  nand _85111_ (_35132_, _35131_, _35125_);
  nor _85112_ (_35134_, _34931_, _11330_);
  nor _85113_ (_35135_, _35134_, _08508_);
  and _85114_ (_35136_, _35135_, _35132_);
  nor _85115_ (_35137_, _11596_, _08507_);
  or _85116_ (_35138_, _35137_, _08587_);
  or _85117_ (_35139_, _35138_, _35136_);
  and _85118_ (_35140_, _34988_, _08587_);
  nor _85119_ (_35141_, _35140_, _03798_);
  nand _85120_ (_35142_, _35141_, _35139_);
  and _85121_ (_35143_, _04620_, _03798_);
  nor _85122_ (_35145_, _35143_, _03188_);
  nand _85123_ (_35146_, _35145_, _35142_);
  nand _85124_ (_35147_, _35146_, _11903_);
  and _85125_ (_35148_, _34906_, _09854_);
  nor _85126_ (_35149_, _11468_, _09854_);
  or _85127_ (_35150_, _35149_, _11903_);
  or _85128_ (_35151_, _35150_, _35148_);
  and _85129_ (_35152_, _35151_, _11328_);
  nand _85130_ (_35153_, _35152_, _35147_);
  nor _85131_ (_35154_, _34931_, _11328_);
  nor _85132_ (_35156_, _35154_, _08703_);
  and _85133_ (_35157_, _35156_, _35153_);
  nor _85134_ (_35158_, _11596_, _08702_);
  or _85135_ (_35159_, _35158_, _08732_);
  or _85136_ (_35160_, _35159_, _35157_);
  and _85137_ (_35161_, _34988_, _08732_);
  nor _85138_ (_35162_, _35161_, _03515_);
  nand _85139_ (_35163_, _35162_, _35160_);
  and _85140_ (_35164_, _04620_, _03515_);
  nor _85141_ (_35165_, _35164_, _03203_);
  nand _85142_ (_35167_, _35165_, _35163_);
  nand _85143_ (_35168_, _35167_, _03816_);
  and _85144_ (_35169_, _11469_, _09854_);
  nor _85145_ (_35170_, _34900_, _09854_);
  nor _85146_ (_35171_, _35170_, _35169_);
  and _85147_ (_35172_, _35171_, _03628_);
  nor _85148_ (_35173_, _35172_, _11934_);
  nand _85149_ (_35174_, _35173_, _35168_);
  nor _85150_ (_35175_, _34931_, _11933_);
  nor _85151_ (_35176_, _35175_, _03815_);
  nand _85152_ (_35178_, _35176_, _35174_);
  and _85153_ (_35179_, _11595_, _03815_);
  nor _85154_ (_35180_, _35179_, _32765_);
  nand _85155_ (_35181_, _35180_, _35178_);
  nor _85156_ (_35182_, _34931_, _11940_);
  nor _85157_ (_35183_, _35182_, _03629_);
  and _85158_ (_35184_, _35183_, _35181_);
  or _85159_ (_35185_, _35184_, _34893_);
  nor _85160_ (_35186_, _03198_, _03453_);
  nand _85161_ (_35187_, _35186_, _35185_);
  and _85162_ (_35189_, _35171_, _03453_);
  nor _85163_ (_35190_, _35189_, _11958_);
  nand _85164_ (_35191_, _35190_, _35187_);
  nor _85165_ (_35192_, _34931_, _11957_);
  nor _85166_ (_35193_, _35192_, _03447_);
  nand _85167_ (_35194_, _35193_, _35191_);
  and _85168_ (_35195_, _11595_, _03447_);
  nor _85169_ (_35196_, _35195_, _33825_);
  nand _85170_ (_35197_, _35196_, _35194_);
  nor _85171_ (_35198_, _34931_, _11964_);
  nor _85172_ (_35200_, _35198_, _03631_);
  and _85173_ (_35201_, _35200_, _35197_);
  or _85174_ (_35202_, _35201_, _34892_);
  and _85175_ (_35203_, _35202_, _24553_);
  and _85176_ (_35204_, _34931_, _11975_);
  or _85177_ (_35205_, _35204_, _35203_);
  or _85178_ (_35206_, _35205_, _43004_);
  or _85179_ (_35207_, _43000_, \oc8051_golden_model_1.PC [8]);
  and _85180_ (_35208_, _35207_, _41806_);
  and _85181_ (_43677_, _35208_, _35206_);
  nor _85182_ (_35210_, _03414_, _11968_);
  nor _85183_ (_35211_, _03414_, _11944_);
  nor _85184_ (_35212_, _11318_, \oc8051_golden_model_1.PC [9]);
  nor _85185_ (_35213_, _35212_, _11319_);
  nor _85186_ (_35214_, _35213_, _11328_);
  nor _85187_ (_35215_, _35213_, _11330_);
  and _85188_ (_35216_, _11408_, _03624_);
  nor _85189_ (_35217_, _35213_, _11335_);
  and _85190_ (_35218_, _11408_, _03622_);
  nor _85191_ (_35219_, _35213_, _11851_);
  and _85192_ (_35221_, _11408_, _03600_);
  nor _85193_ (_35222_, _35213_, _11345_);
  and _85194_ (_35223_, _11542_, _03585_);
  nor _85195_ (_35224_, _35213_, _11350_);
  not _85196_ (_35225_, _35213_);
  and _85197_ (_35226_, _35225_, _10025_);
  and _85198_ (_35227_, _11408_, _09876_);
  nor _85199_ (_35228_, _11473_, _11470_);
  and _85200_ (_35229_, _35228_, _11412_);
  nor _85201_ (_35230_, _35228_, _11412_);
  nor _85202_ (_35232_, _35230_, _35229_);
  nor _85203_ (_35233_, _35232_, _09876_);
  nor _85204_ (_35234_, _35233_, _35227_);
  or _85205_ (_35235_, _35234_, _04107_);
  and _85206_ (_35236_, _35213_, _04422_);
  and _85207_ (_35237_, _11504_, _11542_);
  nor _85208_ (_35238_, _11600_, _11597_);
  and _85209_ (_35239_, _35238_, _11546_);
  nor _85210_ (_35240_, _35238_, _11546_);
  nor _85211_ (_35241_, _35240_, _35239_);
  nor _85212_ (_35243_, _35241_, _11504_);
  or _85213_ (_35244_, _35243_, _35237_);
  nor _85214_ (_35245_, _35244_, _06072_);
  nand _85215_ (_35246_, _35213_, _04064_);
  and _85216_ (_35247_, _11630_, _33169_);
  or _85217_ (_35248_, _35247_, _35213_);
  and _85218_ (_35249_, _11543_, _03979_);
  nor _85219_ (_35250_, _35249_, _11632_);
  or _85220_ (_35251_, _04409_, \oc8051_golden_model_1.PC [9]);
  or _85221_ (_35252_, _35251_, _04729_);
  nand _85222_ (_35254_, _35252_, _35250_);
  nand _85223_ (_35255_, _35254_, _32190_);
  and _85224_ (_35256_, _35255_, _35248_);
  nor _85225_ (_35257_, _35256_, _06073_);
  and _85226_ (_35258_, _35257_, _35246_);
  or _85227_ (_35259_, _35258_, _04422_);
  nor _85228_ (_35260_, _35259_, _35245_);
  or _85229_ (_35261_, _35260_, _35236_);
  and _85230_ (_35262_, _35261_, _04081_);
  not _85231_ (_35263_, _35262_);
  not _85232_ (_35265_, _11362_);
  and _85233_ (_35266_, _11408_, _11369_);
  not _85234_ (_35267_, _35232_);
  and _85235_ (_35268_, _35267_, _11367_);
  nor _85236_ (_35269_, _35268_, _35266_);
  nor _85237_ (_35270_, _35269_, _04081_);
  nor _85238_ (_35271_, _35270_, _35265_);
  and _85239_ (_35272_, _35271_, _35263_);
  nor _85240_ (_35273_, _35213_, _11362_);
  nor _85241_ (_35274_, _35273_, _03715_);
  not _85242_ (_35276_, _35274_);
  nor _85243_ (_35277_, _35276_, _35272_);
  and _85244_ (_35278_, _11542_, _03715_);
  or _85245_ (_35279_, _35278_, _04768_);
  nor _85246_ (_35280_, _35279_, _35277_);
  nor _85247_ (_35281_, _35280_, _03723_);
  and _85248_ (_35282_, _11542_, _03723_);
  nor _85249_ (_35283_, _35282_, _11660_);
  not _85250_ (_35284_, _35283_);
  nor _85251_ (_35285_, _35284_, _35281_);
  nor _85252_ (_35287_, _35213_, _11659_);
  nor _85253_ (_35288_, _35287_, _03729_);
  not _85254_ (_35289_, _35288_);
  or _85255_ (_35290_, _35289_, _35285_);
  and _85256_ (_35291_, _11542_, _03729_);
  nor _85257_ (_35292_, _35291_, _11668_);
  nand _85258_ (_35293_, _35292_, _35290_);
  nor _85259_ (_35294_, _35213_, _11666_);
  nor _85260_ (_35295_, _35294_, _03714_);
  nand _85261_ (_35296_, _35295_, _35293_);
  and _85262_ (_35298_, _11542_, _03714_);
  nor _85263_ (_35299_, _35298_, _11670_);
  nand _85264_ (_35300_, _35299_, _35296_);
  nand _85265_ (_35301_, _35300_, _03510_);
  and _85266_ (_35302_, _11542_, _03508_);
  nor _85267_ (_35303_, _35302_, _09917_);
  and _85268_ (_35304_, _35303_, _35301_);
  and _85269_ (_35305_, _11408_, _09969_);
  nor _85270_ (_35306_, _35232_, _09969_);
  or _85271_ (_35307_, _35306_, _35305_);
  nor _85272_ (_35309_, _35307_, _09921_);
  or _85273_ (_35310_, _35309_, _35304_);
  nand _85274_ (_35311_, _35310_, _09920_);
  and _85275_ (_35312_, _35267_, _10018_);
  and _85276_ (_35313_, _11408_, _11685_);
  or _85277_ (_35314_, _35313_, _09920_);
  or _85278_ (_35315_, _35314_, _35312_);
  nand _85279_ (_35316_, _35315_, _35311_);
  or _85280_ (_35317_, _35316_, _03615_);
  and _85281_ (_35318_, _35317_, _35235_);
  or _85282_ (_35320_, _35318_, _03604_);
  and _85283_ (_35321_, _11408_, _10061_);
  nor _85284_ (_35322_, _35232_, _10061_);
  or _85285_ (_35323_, _35322_, _35321_);
  and _85286_ (_35324_, _35323_, _03604_);
  nor _85287_ (_35325_, _35324_, _10025_);
  and _85288_ (_35326_, _35325_, _35320_);
  or _85289_ (_35327_, _35326_, _35226_);
  nand _85290_ (_35328_, _35327_, _06840_);
  and _85291_ (_35329_, _11543_, _03719_);
  not _85292_ (_35331_, _35329_);
  not _85293_ (_35332_, _11715_);
  and _85294_ (_35333_, _23519_, _35332_);
  and _85295_ (_35334_, _35333_, _35331_);
  and _85296_ (_35335_, _35334_, _11712_);
  and _85297_ (_35336_, _35335_, _11710_);
  nand _85298_ (_35337_, _35336_, _35328_);
  nor _85299_ (_35338_, _32547_, _11543_);
  nor _85300_ (_35339_, _35338_, _11356_);
  nand _85301_ (_35340_, _35339_, _35337_);
  nor _85302_ (_35342_, _35213_, _11355_);
  nor _85303_ (_35343_, _35342_, _03753_);
  and _85304_ (_35344_, _35343_, _35340_);
  and _85305_ (_35345_, _11542_, _03753_);
  or _85306_ (_35346_, _35345_, _35344_);
  nand _85307_ (_35347_, _35346_, _11728_);
  and _85308_ (_35348_, _11542_, _03752_);
  not _85309_ (_35349_, _35348_);
  and _85310_ (_35350_, _35349_, _11350_);
  and _85311_ (_35351_, _35350_, _35347_);
  or _85312_ (_35353_, _35351_, _35224_);
  nand _85313_ (_35354_, _35353_, _08186_);
  nor _85314_ (_35355_, _11542_, _08186_);
  nor _85315_ (_35356_, _35355_, _07912_);
  nand _85316_ (_35357_, _35356_, _35354_);
  nor _85317_ (_35358_, _35225_, _03248_);
  nor _85318_ (_35359_, _35358_, _03505_);
  nand _85319_ (_35360_, _35359_, _35357_);
  and _85320_ (_35361_, _11543_, _03505_);
  nor _85321_ (_35362_, _35361_, _23690_);
  nand _85322_ (_35364_, _35362_, _35360_);
  and _85323_ (_35365_, _11408_, _03625_);
  nor _85324_ (_35366_, _35365_, _33299_);
  nand _85325_ (_35367_, _35366_, _35364_);
  nor _85326_ (_35368_, _11749_, _11542_);
  nor _85327_ (_35369_, _35368_, _03222_);
  nand _85328_ (_35370_, _35369_, _35367_);
  and _85329_ (_35371_, _11408_, _03222_);
  nor _85330_ (_35372_, _35371_, _11758_);
  nand _85331_ (_35373_, _35372_, _35370_);
  nor _85332_ (_35375_, _35213_, _11756_);
  nor _85333_ (_35376_, _35375_, _03585_);
  and _85334_ (_35377_, _35376_, _35373_);
  or _85335_ (_35378_, _35377_, _35223_);
  nand _85336_ (_35379_, _35378_, _35040_);
  nor _85337_ (_35380_, _35241_, _11765_);
  nor _85338_ (_35381_, _35380_, _06168_);
  nand _85339_ (_35382_, _35381_, _35379_);
  nor _85340_ (_35383_, _11542_, _05894_);
  nor _85341_ (_35384_, _35383_, _03601_);
  nand _85342_ (_35386_, _35384_, _35382_);
  and _85343_ (_35387_, _11408_, _03601_);
  nor _85344_ (_35388_, _35387_, _08363_);
  nand _85345_ (_35389_, _35388_, _35386_);
  and _85346_ (_35390_, _11543_, _08363_);
  nor _85347_ (_35391_, _35390_, _11347_);
  and _85348_ (_35392_, _35391_, _35389_);
  nor _85349_ (_35393_, _11804_, \oc8051_golden_model_1.DPH [1]);
  not _85350_ (_35394_, _35393_);
  nor _85351_ (_35395_, _11805_, _11348_);
  and _85352_ (_35397_, _35395_, _35394_);
  or _85353_ (_35398_, _35397_, _35392_);
  nand _85354_ (_35399_, _35398_, _10263_);
  and _85355_ (_35400_, _11542_, _03584_);
  nor _85356_ (_35401_, _35400_, _03178_);
  nand _85357_ (_35402_, _35401_, _35399_);
  nand _85358_ (_35403_, _35402_, _11820_);
  and _85359_ (_35404_, _11542_, _08786_);
  nor _85360_ (_35405_, _35241_, _08786_);
  or _85361_ (_35406_, _35405_, _35404_);
  and _85362_ (_35408_, _35406_, _11819_);
  nor _85363_ (_35409_, _35408_, _11824_);
  and _85364_ (_35410_, _35409_, _35403_);
  or _85365_ (_35411_, _35410_, _35222_);
  nand _85366_ (_35412_, _35411_, _11341_);
  nor _85367_ (_35413_, _11542_, _11341_);
  nor _85368_ (_35414_, _35413_, _03600_);
  and _85369_ (_35415_, _35414_, _35412_);
  or _85370_ (_35416_, _35415_, _35221_);
  nand _85371_ (_35417_, _35416_, _07778_);
  and _85372_ (_35419_, _11542_, _03780_);
  nor _85373_ (_35420_, _35419_, _03182_);
  nand _85374_ (_35421_, _35420_, _35417_);
  nand _85375_ (_35422_, _35421_, _11842_);
  nand _85376_ (_35423_, _35241_, _08786_);
  or _85377_ (_35424_, _11542_, _08786_);
  and _85378_ (_35425_, _35424_, _11841_);
  and _85379_ (_35426_, _35425_, _35423_);
  nor _85380_ (_35427_, _35426_, _11853_);
  and _85381_ (_35428_, _35427_, _35422_);
  or _85382_ (_35430_, _35428_, _35219_);
  nand _85383_ (_35431_, _35430_, _08430_);
  nor _85384_ (_35432_, _11542_, _08430_);
  nor _85385_ (_35433_, _35432_, _03622_);
  and _85386_ (_35434_, _35433_, _35431_);
  or _85387_ (_35435_, _35434_, _35218_);
  nand _85388_ (_35436_, _35435_, _06828_);
  and _85389_ (_35437_, _11542_, _03790_);
  nor _85390_ (_35438_, _35437_, _03192_);
  nand _85391_ (_35439_, _35438_, _35436_);
  nand _85392_ (_35441_, _35439_, _11338_);
  and _85393_ (_35442_, _11542_, \oc8051_golden_model_1.PSW [7]);
  nor _85394_ (_35443_, _35241_, \oc8051_golden_model_1.PSW [7]);
  or _85395_ (_35444_, _35443_, _35442_);
  and _85396_ (_35445_, _35444_, _11337_);
  nor _85397_ (_35446_, _35445_, _11864_);
  and _85398_ (_35447_, _35446_, _35441_);
  or _85399_ (_35448_, _35447_, _35217_);
  nand _85400_ (_35449_, _35448_, _08459_);
  nor _85401_ (_35450_, _11542_, _08459_);
  nor _85402_ (_35452_, _35450_, _03624_);
  and _85403_ (_35453_, _35452_, _35449_);
  or _85404_ (_35454_, _35453_, _35216_);
  nand _85405_ (_35455_, _35454_, _07793_);
  and _85406_ (_35456_, _11542_, _03785_);
  nor _85407_ (_35457_, _35456_, _03201_);
  nand _85408_ (_35458_, _35457_, _35455_);
  nand _85409_ (_35459_, _35458_, _11881_);
  and _85410_ (_35460_, _35241_, \oc8051_golden_model_1.PSW [7]);
  nor _85411_ (_35461_, _11542_, \oc8051_golden_model_1.PSW [7]);
  nor _85412_ (_35463_, _35461_, _11881_);
  not _85413_ (_35464_, _35463_);
  nor _85414_ (_35465_, _35464_, _35460_);
  nor _85415_ (_35466_, _35465_, _11885_);
  and _85416_ (_35467_, _35466_, _35459_);
  or _85417_ (_35468_, _35467_, _35215_);
  nand _85418_ (_35469_, _35468_, _08507_);
  nor _85419_ (_35470_, _11542_, _08507_);
  nor _85420_ (_35471_, _35470_, _08587_);
  nand _85421_ (_35472_, _35471_, _35469_);
  and _85422_ (_35474_, _35213_, _08587_);
  nor _85423_ (_35475_, _35474_, _03798_);
  nand _85424_ (_35476_, _35475_, _35472_);
  nor _85425_ (_35477_, _03621_, _03188_);
  not _85426_ (_35478_, _35477_);
  and _85427_ (_35479_, _04406_, _03798_);
  nor _85428_ (_35480_, _35479_, _35478_);
  nand _85429_ (_35481_, _35480_, _35476_);
  and _85430_ (_35482_, _35267_, _09854_);
  nor _85431_ (_35483_, _11409_, _09854_);
  nor _85432_ (_35485_, _35483_, _35482_);
  nor _85433_ (_35486_, _35485_, _11903_);
  nor _85434_ (_35487_, _35486_, _11907_);
  and _85435_ (_35488_, _35487_, _35481_);
  or _85436_ (_35489_, _35488_, _35214_);
  nand _85437_ (_35490_, _35489_, _08702_);
  nor _85438_ (_35491_, _11542_, _08702_);
  nor _85439_ (_35492_, _35491_, _08732_);
  nand _85440_ (_35493_, _35492_, _35490_);
  and _85441_ (_35494_, _35213_, _08732_);
  nor _85442_ (_35497_, _35494_, _03515_);
  nand _85443_ (_35498_, _35497_, _35493_);
  not _85444_ (_35499_, _23212_);
  and _85445_ (_35500_, _04406_, _03515_);
  nor _85446_ (_35501_, _35500_, _35499_);
  nand _85447_ (_35502_, _35501_, _35498_);
  nor _85448_ (_35503_, _35267_, _09854_);
  and _85449_ (_35504_, _11409_, _09854_);
  nor _85450_ (_35505_, _35504_, _35503_);
  and _85451_ (_35506_, _35505_, _03628_);
  nor _85452_ (_35508_, _35506_, _11934_);
  nand _85453_ (_35509_, _35508_, _35502_);
  nor _85454_ (_35510_, _35213_, _11933_);
  nor _85455_ (_35511_, _35510_, _03815_);
  nand _85456_ (_35512_, _35511_, _35509_);
  and _85457_ (_35513_, _11542_, _03815_);
  nor _85458_ (_35514_, _35513_, _32765_);
  nand _85459_ (_35515_, _35514_, _35512_);
  nor _85460_ (_35516_, _35213_, _11940_);
  nor _85461_ (_35517_, _35516_, _03629_);
  and _85462_ (_35520_, _35517_, _35515_);
  or _85463_ (_35521_, _35520_, _35211_);
  nand _85464_ (_35522_, _35521_, _35186_);
  and _85465_ (_35523_, _35505_, _03453_);
  nor _85466_ (_35524_, _35523_, _11958_);
  nand _85467_ (_35525_, _35524_, _35522_);
  nor _85468_ (_35526_, _35213_, _11957_);
  nor _85469_ (_35527_, _35526_, _03447_);
  nand _85470_ (_35528_, _35527_, _35525_);
  and _85471_ (_35529_, _11542_, _03447_);
  nor _85472_ (_35531_, _35529_, _33825_);
  nand _85473_ (_35532_, _35531_, _35528_);
  nor _85474_ (_35533_, _35213_, _11964_);
  nor _85475_ (_35534_, _35533_, _03631_);
  and _85476_ (_35535_, _35534_, _35532_);
  or _85477_ (_35536_, _35535_, _35210_);
  and _85478_ (_35537_, _35536_, _24553_);
  and _85479_ (_35538_, _35213_, _11975_);
  or _85480_ (_35539_, _35538_, _35537_);
  or _85481_ (_35540_, _35539_, _43004_);
  or _85482_ (_35543_, _43000_, \oc8051_golden_model_1.PC [9]);
  and _85483_ (_35544_, _35543_, _41806_);
  and _85484_ (_43678_, _35544_, _35540_);
  nor _85485_ (_35545_, _11319_, \oc8051_golden_model_1.PC [10]);
  nor _85486_ (_35546_, _35545_, _11320_);
  and _85487_ (_35547_, _35546_, _11975_);
  or _85488_ (_35548_, _35546_, _11957_);
  not _85489_ (_35549_, _35546_);
  nand _85490_ (_35550_, _35549_, _08732_);
  nand _85491_ (_35551_, _35549_, _08587_);
  nand _85492_ (_35553_, _11395_, _03624_);
  nand _85493_ (_35554_, _11395_, _03622_);
  nor _85494_ (_35555_, _35549_, _11756_);
  or _85495_ (_35556_, _11529_, _08186_);
  nor _85496_ (_35557_, _35549_, _11666_);
  or _85497_ (_35558_, _35546_, _11659_);
  nor _85498_ (_35559_, _35549_, _11653_);
  nor _85499_ (_35560_, _11477_, _11474_);
  not _85500_ (_35561_, _35560_);
  and _85501_ (_35562_, _35561_, _11405_);
  nor _85502_ (_35565_, _35561_, _11405_);
  nor _85503_ (_35566_, _35565_, _35562_);
  or _85504_ (_35567_, _35566_, _11369_);
  or _85505_ (_35568_, _11394_, _11367_);
  and _85506_ (_35569_, _35568_, _03610_);
  and _85507_ (_35570_, _35569_, _35567_);
  nor _85508_ (_35571_, _11604_, _11601_);
  not _85509_ (_35572_, _35571_);
  and _85510_ (_35573_, _35572_, _11539_);
  nor _85511_ (_35574_, _35572_, _11539_);
  nor _85512_ (_35576_, _35574_, _35573_);
  and _85513_ (_35577_, _35576_, _11624_);
  and _85514_ (_35578_, _11504_, _11529_);
  or _85515_ (_35579_, _35578_, _06072_);
  or _85516_ (_35580_, _35579_, _35577_);
  or _85517_ (_35581_, _35546_, _11643_);
  not _85518_ (_35582_, _03979_);
  or _85519_ (_35583_, _11529_, _35582_);
  or _85520_ (_35584_, _04409_, \oc8051_golden_model_1.PC [10]);
  or _85521_ (_35585_, _35584_, _04729_);
  and _85522_ (_35587_, _35585_, _35583_);
  nand _85523_ (_35588_, _11630_, _32815_);
  or _85524_ (_35589_, _35588_, _35587_);
  and _85525_ (_35590_, _35589_, _35581_);
  or _85526_ (_35591_, _06073_, _03980_);
  or _85527_ (_35592_, _35591_, _35590_);
  and _85528_ (_35593_, _35592_, _11647_);
  and _85529_ (_35594_, _35593_, _35580_);
  or _85530_ (_35595_, _35594_, _35570_);
  and _85531_ (_35596_, _35595_, _11362_);
  or _85532_ (_35598_, _35596_, _35559_);
  and _85533_ (_35599_, _35598_, _03730_);
  and _85534_ (_35600_, _11529_, _14265_);
  nor _85535_ (_35601_, _35600_, _04768_);
  nand _85536_ (_35602_, _35601_, _11659_);
  or _85537_ (_35603_, _35602_, _35599_);
  and _85538_ (_35604_, _35603_, _35558_);
  or _85539_ (_35605_, _35604_, _03729_);
  or _85540_ (_35606_, _11529_, _03737_);
  and _85541_ (_35607_, _35606_, _11666_);
  and _85542_ (_35609_, _35607_, _35605_);
  or _85543_ (_35610_, _35609_, _35557_);
  and _85544_ (_35611_, _35610_, _03736_);
  and _85545_ (_35612_, _11529_, _03714_);
  or _85546_ (_35613_, _35612_, _11670_);
  or _85547_ (_35614_, _35613_, _35611_);
  and _85548_ (_35615_, _35614_, _03510_);
  and _85549_ (_35616_, _11529_, _03508_);
  or _85550_ (_35617_, _35616_, _09917_);
  or _85551_ (_35618_, _35617_, _35615_);
  or _85552_ (_35620_, _35566_, _09969_);
  nand _85553_ (_35621_, _11395_, _09969_);
  and _85554_ (_35622_, _35621_, _35620_);
  or _85555_ (_35623_, _35622_, _09921_);
  and _85556_ (_35624_, _35623_, _35618_);
  or _85557_ (_35625_, _35624_, _32519_);
  and _85558_ (_35626_, _11394_, _11685_);
  and _85559_ (_35627_, _35566_, _10018_);
  or _85560_ (_35628_, _35627_, _35626_);
  or _85561_ (_35629_, _35628_, _09920_);
  and _85562_ (_35631_, _35629_, _35625_);
  or _85563_ (_35632_, _35631_, _03615_);
  and _85564_ (_35633_, _11394_, _09876_);
  and _85565_ (_35634_, _35566_, _11693_);
  or _85566_ (_35635_, _35634_, _04107_);
  or _85567_ (_35636_, _35635_, _35633_);
  and _85568_ (_35637_, _35636_, _09856_);
  and _85569_ (_35638_, _35637_, _35632_);
  or _85570_ (_35639_, _35566_, _10061_);
  nand _85571_ (_35640_, _11395_, _10061_);
  and _85572_ (_35642_, _35640_, _03604_);
  and _85573_ (_35643_, _35642_, _35639_);
  or _85574_ (_35644_, _35643_, _10025_);
  or _85575_ (_35645_, _35644_, _35638_);
  nand _85576_ (_35646_, _35549_, _10025_);
  and _85577_ (_35647_, _32547_, _06840_);
  and _85578_ (_35648_, _35647_, _35646_);
  and _85579_ (_35649_, _35648_, _35645_);
  not _85580_ (_35650_, _11529_);
  nor _85581_ (_35651_, _35647_, _35650_);
  nand _85582_ (_35653_, _11355_, _03227_);
  or _85583_ (_35654_, _35653_, _35651_);
  or _85584_ (_35655_, _35654_, _35649_);
  or _85585_ (_35656_, _35546_, _11355_);
  and _85586_ (_35657_, _35656_, _09669_);
  and _85587_ (_35658_, _35657_, _35655_);
  nand _85588_ (_35659_, _11529_, _03753_);
  nand _85589_ (_35660_, _35659_, _11728_);
  or _85590_ (_35661_, _35660_, _35658_);
  nand _85591_ (_35662_, _35650_, _03752_);
  and _85592_ (_35664_, _35662_, _11350_);
  and _85593_ (_35665_, _35664_, _35661_);
  nor _85594_ (_35666_, _35549_, _11350_);
  or _85595_ (_35667_, _35666_, _08187_);
  or _85596_ (_35668_, _35667_, _35665_);
  and _85597_ (_35669_, _35668_, _35556_);
  or _85598_ (_35670_, _35669_, _07912_);
  or _85599_ (_35671_, _35546_, _03248_);
  and _85600_ (_35672_, _35671_, _03710_);
  and _85601_ (_35673_, _35672_, _35670_);
  nand _85602_ (_35675_, _11529_, _03505_);
  nand _85603_ (_35676_, _35675_, _23689_);
  or _85604_ (_35677_, _35676_, _35673_);
  nand _85605_ (_35678_, _11395_, _03625_);
  and _85606_ (_35679_, _35678_, _11749_);
  and _85607_ (_35680_, _35679_, _35677_);
  nor _85608_ (_35681_, _11749_, _35650_);
  or _85609_ (_35682_, _35681_, _03222_);
  or _85610_ (_35683_, _35682_, _35680_);
  nand _85611_ (_35684_, _11395_, _03222_);
  and _85612_ (_35686_, _35684_, _11756_);
  and _85613_ (_35687_, _35686_, _35683_);
  nor _85614_ (_35688_, _35687_, _35555_);
  nor _85615_ (_35689_, _35688_, _03585_);
  nand _85616_ (_35690_, _11529_, _03585_);
  nand _85617_ (_35691_, _35690_, _35040_);
  or _85618_ (_35692_, _35691_, _35689_);
  or _85619_ (_35693_, _35576_, _11765_);
  and _85620_ (_35694_, _35693_, _05894_);
  and _85621_ (_35695_, _35694_, _35692_);
  nor _85622_ (_35697_, _35650_, _05894_);
  or _85623_ (_35698_, _35697_, _03601_);
  or _85624_ (_35699_, _35698_, _35695_);
  nand _85625_ (_35700_, _11395_, _03601_);
  and _85626_ (_35701_, _35700_, _08364_);
  and _85627_ (_35702_, _35701_, _35699_);
  and _85628_ (_35703_, _11529_, _08363_);
  or _85629_ (_35704_, _35703_, _11347_);
  or _85630_ (_35705_, _35704_, _35702_);
  nor _85631_ (_35706_, _11805_, \oc8051_golden_model_1.DPH [2]);
  nor _85632_ (_35708_, _35706_, _11806_);
  or _85633_ (_35709_, _35708_, _11348_);
  and _85634_ (_35710_, _35709_, _10263_);
  and _85635_ (_35711_, _35710_, _35705_);
  and _85636_ (_35712_, _11529_, _03584_);
  or _85637_ (_35713_, _35712_, _35711_);
  nor _85638_ (_35714_, _11819_, _03178_);
  and _85639_ (_35715_, _35714_, _35713_);
  or _85640_ (_35716_, _35576_, _08786_);
  or _85641_ (_35717_, _11529_, _11826_);
  and _85642_ (_35719_, _35717_, _11819_);
  and _85643_ (_35720_, _35719_, _35716_);
  or _85644_ (_35721_, _35720_, _11824_);
  or _85645_ (_35722_, _35721_, _35715_);
  or _85646_ (_35723_, _35546_, _11345_);
  and _85647_ (_35724_, _35723_, _11341_);
  and _85648_ (_35725_, _35724_, _35722_);
  and _85649_ (_35726_, _11529_, _11342_);
  or _85650_ (_35727_, _35726_, _03600_);
  or _85651_ (_35728_, _35727_, _35725_);
  nand _85652_ (_35730_, _11395_, _03600_);
  and _85653_ (_35731_, _35730_, _35728_);
  or _85654_ (_35732_, _35731_, _03780_);
  nand _85655_ (_35733_, _35650_, _03780_);
  and _85656_ (_35734_, _35733_, _23991_);
  and _85657_ (_35735_, _35734_, _35732_);
  or _85658_ (_35736_, _35576_, _11826_);
  or _85659_ (_35737_, _11529_, _08786_);
  and _85660_ (_35738_, _35737_, _11841_);
  and _85661_ (_35739_, _35738_, _35736_);
  or _85662_ (_35741_, _35739_, _11853_);
  or _85663_ (_35742_, _35741_, _35735_);
  or _85664_ (_35743_, _35546_, _11851_);
  and _85665_ (_35744_, _35743_, _08430_);
  and _85666_ (_35745_, _35744_, _35742_);
  nor _85667_ (_35746_, _35650_, _08430_);
  or _85668_ (_35747_, _35746_, _03622_);
  or _85669_ (_35748_, _35747_, _35745_);
  and _85670_ (_35749_, _35748_, _35554_);
  or _85671_ (_35750_, _35749_, _03790_);
  nand _85672_ (_35752_, _35650_, _03790_);
  and _85673_ (_35753_, _35752_, _34895_);
  and _85674_ (_35754_, _35753_, _35750_);
  or _85675_ (_35755_, _35576_, \oc8051_golden_model_1.PSW [7]);
  or _85676_ (_35756_, _11529_, _07871_);
  and _85677_ (_35757_, _35756_, _11337_);
  and _85678_ (_35758_, _35757_, _35755_);
  or _85679_ (_35759_, _35758_, _11864_);
  or _85680_ (_35760_, _35759_, _35754_);
  or _85681_ (_35761_, _35546_, _11335_);
  and _85682_ (_35763_, _35761_, _08459_);
  and _85683_ (_35764_, _35763_, _35760_);
  nor _85684_ (_35765_, _35650_, _08459_);
  or _85685_ (_35766_, _35765_, _03624_);
  or _85686_ (_35767_, _35766_, _35764_);
  and _85687_ (_35768_, _35767_, _35553_);
  or _85688_ (_35769_, _35768_, _03785_);
  nand _85689_ (_35770_, _35650_, _03785_);
  and _85690_ (_35771_, _35770_, _35120_);
  and _85691_ (_35772_, _35771_, _35769_);
  or _85692_ (_35774_, _35576_, _07871_);
  or _85693_ (_35775_, _11529_, \oc8051_golden_model_1.PSW [7]);
  and _85694_ (_35776_, _35775_, _11880_);
  and _85695_ (_35777_, _35776_, _35774_);
  or _85696_ (_35778_, _35777_, _11885_);
  or _85697_ (_35779_, _35778_, _35772_);
  or _85698_ (_35780_, _35546_, _11330_);
  and _85699_ (_35781_, _35780_, _08507_);
  and _85700_ (_35782_, _35781_, _35779_);
  nor _85701_ (_35783_, _35650_, _08507_);
  or _85702_ (_35785_, _35783_, _08587_);
  or _85703_ (_35786_, _35785_, _35782_);
  and _85704_ (_35787_, _35786_, _35551_);
  or _85705_ (_35788_, _35787_, _03798_);
  nand _85706_ (_35789_, _04875_, _03798_);
  and _85707_ (_35790_, _35789_, _35477_);
  and _85708_ (_35791_, _35790_, _35788_);
  or _85709_ (_35792_, _35566_, _11908_);
  or _85710_ (_35793_, _11394_, _09854_);
  and _85711_ (_35794_, _35793_, _03621_);
  and _85712_ (_35796_, _35794_, _35792_);
  or _85713_ (_35797_, _35796_, _11907_);
  or _85714_ (_35798_, _35797_, _35791_);
  or _85715_ (_35799_, _35546_, _11328_);
  and _85716_ (_35800_, _35799_, _08702_);
  and _85717_ (_35801_, _35800_, _35798_);
  nor _85718_ (_35802_, _35650_, _08702_);
  or _85719_ (_35803_, _35802_, _08732_);
  or _85720_ (_35804_, _35803_, _35801_);
  and _85721_ (_35805_, _35804_, _35550_);
  or _85722_ (_35807_, _35805_, _03515_);
  nand _85723_ (_35808_, _04875_, _03515_);
  and _85724_ (_35809_, _35808_, _23212_);
  and _85725_ (_35810_, _35809_, _35807_);
  or _85726_ (_35811_, _35566_, _09854_);
  nand _85727_ (_35812_, _11395_, _09854_);
  and _85728_ (_35813_, _35812_, _35811_);
  and _85729_ (_35814_, _35813_, _03628_);
  or _85730_ (_35815_, _35814_, _11934_);
  or _85731_ (_35816_, _35815_, _35810_);
  or _85732_ (_35818_, _35546_, _11933_);
  and _85733_ (_35819_, _35818_, _35816_);
  or _85734_ (_35820_, _35819_, _03815_);
  nand _85735_ (_35821_, _35650_, _03815_);
  and _85736_ (_35822_, _35821_, _11940_);
  and _85737_ (_35823_, _35822_, _35820_);
  nor _85738_ (_35824_, _35549_, _11940_);
  or _85739_ (_35825_, _35824_, _03629_);
  or _85740_ (_35826_, _35825_, _35823_);
  nand _85741_ (_35827_, _03904_, _03629_);
  and _85742_ (_35829_, _35827_, _35186_);
  and _85743_ (_35830_, _35829_, _35826_);
  and _85744_ (_35831_, _35813_, _03453_);
  or _85745_ (_35832_, _35831_, _11958_);
  or _85746_ (_35833_, _35832_, _35830_);
  and _85747_ (_35834_, _35833_, _35548_);
  or _85748_ (_35835_, _35834_, _03447_);
  nand _85749_ (_35836_, _35650_, _03447_);
  and _85750_ (_35837_, _35836_, _11964_);
  and _85751_ (_35838_, _35837_, _35835_);
  nor _85752_ (_35840_, _35549_, _11964_);
  or _85753_ (_35841_, _35840_, _03631_);
  or _85754_ (_35842_, _35841_, _35838_);
  nand _85755_ (_35843_, _03904_, _03631_);
  and _85756_ (_35844_, _35843_, _24553_);
  and _85757_ (_35845_, _35844_, _35842_);
  or _85758_ (_35846_, _35845_, _35547_);
  or _85759_ (_35847_, _35846_, _43004_);
  or _85760_ (_35848_, _43000_, \oc8051_golden_model_1.PC [10]);
  and _85761_ (_35849_, _35848_, _41806_);
  and _85762_ (_43679_, _35849_, _35847_);
  nor _85763_ (_35851_, _11320_, \oc8051_golden_model_1.PC [11]);
  nor _85764_ (_35852_, _35851_, _11321_);
  nor _85765_ (_35853_, _35852_, _11328_);
  nor _85766_ (_35854_, _35852_, _11330_);
  nor _85767_ (_35855_, _35852_, _11335_);
  nor _85768_ (_35856_, _35852_, _11851_);
  nor _85769_ (_35857_, _35852_, _11345_);
  nor _85770_ (_35858_, _11533_, _05894_);
  and _85771_ (_35859_, _11399_, _03222_);
  and _85772_ (_35861_, _11399_, _10061_);
  nor _85773_ (_35862_, _35562_, _11396_);
  and _85774_ (_35863_, _35862_, _11403_);
  nor _85775_ (_35864_, _35862_, _11403_);
  nor _85776_ (_35865_, _35864_, _35863_);
  nor _85777_ (_35866_, _35865_, _10061_);
  or _85778_ (_35867_, _35866_, _35861_);
  and _85779_ (_35868_, _35867_, _03604_);
  and _85780_ (_35869_, _11399_, _11685_);
  not _85781_ (_35870_, _35865_);
  and _85782_ (_35872_, _35870_, _10018_);
  or _85783_ (_35873_, _35872_, _35869_);
  nor _85784_ (_35874_, _35873_, _09920_);
  and _85785_ (_35875_, _11533_, _03729_);
  nor _85786_ (_35876_, _11360_, _11533_);
  and _85787_ (_35877_, _11400_, _11369_);
  and _85788_ (_35878_, _35865_, _11367_);
  or _85789_ (_35879_, _35878_, _04081_);
  or _85790_ (_35880_, _35879_, _35877_);
  and _85791_ (_35881_, _11504_, _11533_);
  not _85792_ (_35883_, _35881_);
  nor _85793_ (_35884_, _35573_, _11530_);
  and _85794_ (_35885_, _35884_, _11537_);
  nor _85795_ (_35886_, _35884_, _11537_);
  nor _85796_ (_35887_, _35886_, _35885_);
  nor _85797_ (_35888_, _35887_, _11504_);
  nor _85798_ (_35889_, _35888_, _06072_);
  and _85799_ (_35890_, _35889_, _35883_);
  nor _85800_ (_35891_, _35852_, _11643_);
  and _85801_ (_35892_, _11534_, _03980_);
  and _85802_ (_35894_, _11534_, _03979_);
  nor _85803_ (_35895_, _04409_, \oc8051_golden_model_1.PC [11]);
  and _85804_ (_35896_, _35895_, _11634_);
  nor _85805_ (_35897_, _35896_, _35894_);
  nor _85806_ (_35898_, _35897_, _11632_);
  nor _85807_ (_35899_, _35898_, _35892_);
  nor _85808_ (_35900_, _35899_, _11631_);
  nor _85809_ (_35901_, _35900_, _35891_);
  nor _85810_ (_35902_, _35901_, _06073_);
  or _85811_ (_35903_, _35902_, _33523_);
  or _85812_ (_35905_, _35903_, _35890_);
  and _85813_ (_35906_, _35905_, _35880_);
  or _85814_ (_35907_, _35906_, _35265_);
  not _85815_ (_35908_, _35852_);
  or _85816_ (_35909_, _35908_, _11653_);
  and _85817_ (_35910_, _35909_, _11360_);
  and _85818_ (_35911_, _35910_, _35907_);
  nor _85819_ (_35912_, _35911_, _35876_);
  nor _85820_ (_35913_, _35912_, _11660_);
  nor _85821_ (_35914_, _35852_, _11659_);
  nor _85822_ (_35916_, _35914_, _03729_);
  not _85823_ (_35917_, _35916_);
  nor _85824_ (_35918_, _35917_, _35913_);
  nor _85825_ (_35919_, _35918_, _35875_);
  nor _85826_ (_35920_, _35919_, _11668_);
  nor _85827_ (_35921_, _35908_, _11666_);
  nor _85828_ (_35922_, _35921_, _11673_);
  not _85829_ (_35923_, _35922_);
  or _85830_ (_35924_, _35923_, _35920_);
  nor _85831_ (_35925_, _11672_, _11533_);
  nor _85832_ (_35927_, _35925_, _09917_);
  and _85833_ (_35928_, _35927_, _35924_);
  or _85834_ (_35929_, _35870_, _09969_);
  nand _85835_ (_35930_, _11400_, _09969_);
  and _85836_ (_35931_, _35930_, _09917_);
  and _85837_ (_35932_, _35931_, _35929_);
  or _85838_ (_35933_, _35932_, _09919_);
  nor _85839_ (_35934_, _35933_, _35928_);
  or _85840_ (_35935_, _35934_, _35874_);
  or _85841_ (_35936_, _35935_, _03615_);
  and _85842_ (_35938_, _11399_, _09876_);
  nor _85843_ (_35939_, _35865_, _09876_);
  nor _85844_ (_35940_, _35939_, _35938_);
  or _85845_ (_35941_, _35940_, _04107_);
  and _85846_ (_35942_, _35941_, _35936_);
  nor _85847_ (_35943_, _35942_, _03604_);
  or _85848_ (_35944_, _35943_, _35868_);
  nand _85849_ (_35945_, _35944_, _11358_);
  and _85850_ (_35946_, _35852_, _10025_);
  not _85851_ (_35947_, _35946_);
  and _85852_ (_35949_, _35947_, _11720_);
  nand _85853_ (_35950_, _35949_, _35945_);
  nor _85854_ (_35951_, _11720_, _11533_);
  nor _85855_ (_35952_, _35951_, _11356_);
  nand _85856_ (_35953_, _35952_, _35950_);
  not _85857_ (_35954_, _11729_);
  nor _85858_ (_35955_, _35908_, _11355_);
  nor _85859_ (_35956_, _35955_, _35954_);
  and _85860_ (_35957_, _35956_, _35953_);
  or _85861_ (_35958_, _11729_, _11533_);
  nand _85862_ (_35960_, _35958_, _11350_);
  or _85863_ (_35961_, _35960_, _35957_);
  nor _85864_ (_35962_, _35908_, _11350_);
  nor _85865_ (_35963_, _35962_, _08187_);
  nand _85866_ (_35964_, _35963_, _35961_);
  nor _85867_ (_35965_, _11533_, _08186_);
  nor _85868_ (_35966_, _35965_, _07912_);
  nand _85869_ (_35967_, _35966_, _35964_);
  nor _85870_ (_35968_, _35908_, _03248_);
  nor _85871_ (_35969_, _35968_, _11741_);
  nand _85872_ (_35971_, _35969_, _35967_);
  nor _85873_ (_35972_, _11740_, _11533_);
  nor _85874_ (_35973_, _35972_, _03625_);
  nand _85875_ (_35974_, _35973_, _35971_);
  and _85876_ (_35975_, _11399_, _03625_);
  nor _85877_ (_35976_, _35975_, _33299_);
  nand _85878_ (_35977_, _35976_, _35974_);
  nor _85879_ (_35978_, _11749_, _11533_);
  nor _85880_ (_35979_, _35978_, _03222_);
  and _85881_ (_35980_, _35979_, _35977_);
  or _85882_ (_35982_, _35980_, _35859_);
  nand _85883_ (_35983_, _35982_, _11756_);
  nor _85884_ (_35984_, _35908_, _11756_);
  nor _85885_ (_35985_, _35984_, _11761_);
  nand _85886_ (_35986_, _35985_, _35983_);
  nor _85887_ (_35987_, _11760_, _11533_);
  nor _85888_ (_35988_, _35987_, _11764_);
  nand _85889_ (_35989_, _35988_, _35986_);
  nor _85890_ (_35990_, _35887_, _11765_);
  nor _85891_ (_35991_, _35990_, _06168_);
  and _85892_ (_35993_, _35991_, _35989_);
  or _85893_ (_35994_, _35993_, _35858_);
  nand _85894_ (_35995_, _35994_, _05886_);
  and _85895_ (_35996_, _11400_, _03601_);
  nor _85896_ (_35997_, _35996_, _08363_);
  and _85897_ (_35998_, _35997_, _35995_);
  and _85898_ (_35999_, _11533_, _08363_);
  or _85899_ (_36000_, _35999_, _35998_);
  nand _85900_ (_36001_, _36000_, _11348_);
  nor _85901_ (_36002_, _11806_, \oc8051_golden_model_1.DPH [3]);
  not _85902_ (_36004_, _36002_);
  nor _85903_ (_36005_, _11807_, _11348_);
  and _85904_ (_36006_, _36005_, _36004_);
  nor _85905_ (_36007_, _36006_, _11816_);
  nand _85906_ (_36008_, _36007_, _36001_);
  nor _85907_ (_36009_, _11815_, _11533_);
  nor _85908_ (_36010_, _36009_, _11819_);
  nand _85909_ (_36011_, _36010_, _36008_);
  and _85910_ (_36012_, _11533_, _08786_);
  nor _85911_ (_36013_, _35887_, _08786_);
  or _85912_ (_36015_, _36013_, _36012_);
  and _85913_ (_36016_, _36015_, _11819_);
  nor _85914_ (_36017_, _36016_, _11824_);
  and _85915_ (_36018_, _36017_, _36011_);
  or _85916_ (_36019_, _36018_, _35857_);
  nand _85917_ (_36020_, _36019_, _11341_);
  nor _85918_ (_36021_, _11533_, _11341_);
  nor _85919_ (_36022_, _36021_, _03600_);
  nand _85920_ (_36023_, _36022_, _36020_);
  not _85921_ (_36024_, _11838_);
  and _85922_ (_36026_, _11399_, _03600_);
  nor _85923_ (_36027_, _36026_, _36024_);
  nand _85924_ (_36028_, _36027_, _36023_);
  nor _85925_ (_36029_, _11838_, _11533_);
  nor _85926_ (_36030_, _36029_, _11841_);
  nand _85927_ (_36031_, _36030_, _36028_);
  nand _85928_ (_36032_, _35887_, _08786_);
  or _85929_ (_36033_, _11533_, _08786_);
  and _85930_ (_36034_, _36033_, _11841_);
  and _85931_ (_36035_, _36034_, _36032_);
  nor _85932_ (_36037_, _36035_, _11853_);
  and _85933_ (_36038_, _36037_, _36031_);
  or _85934_ (_36039_, _36038_, _35856_);
  nand _85935_ (_36040_, _36039_, _08430_);
  nor _85936_ (_36041_, _11533_, _08430_);
  nor _85937_ (_36042_, _36041_, _03622_);
  nand _85938_ (_36043_, _36042_, _36040_);
  and _85939_ (_36044_, _11399_, _03622_);
  nor _85940_ (_36045_, _36044_, _10754_);
  and _85941_ (_36046_, _36045_, _36043_);
  nor _85942_ (_36048_, _11534_, _11337_);
  nor _85943_ (_36049_, _36048_, _24116_);
  or _85944_ (_36050_, _36049_, _36046_);
  and _85945_ (_36051_, _11533_, \oc8051_golden_model_1.PSW [7]);
  nor _85946_ (_36052_, _35887_, \oc8051_golden_model_1.PSW [7]);
  or _85947_ (_36053_, _36052_, _36051_);
  and _85948_ (_36054_, _36053_, _11337_);
  nor _85949_ (_36055_, _36054_, _11864_);
  and _85950_ (_36056_, _36055_, _36050_);
  or _85951_ (_36057_, _36056_, _35855_);
  nand _85952_ (_36059_, _36057_, _08459_);
  nor _85953_ (_36060_, _11533_, _08459_);
  nor _85954_ (_36061_, _36060_, _03624_);
  nand _85955_ (_36062_, _36061_, _36059_);
  not _85956_ (_36063_, _11877_);
  and _85957_ (_36064_, _11399_, _03624_);
  nor _85958_ (_36065_, _36064_, _36063_);
  and _85959_ (_36066_, _36065_, _36062_);
  nor _85960_ (_36067_, _11880_, _11534_);
  nor _85961_ (_36068_, _36067_, _24239_);
  or _85962_ (_36070_, _36068_, _36066_);
  and _85963_ (_36071_, _35887_, \oc8051_golden_model_1.PSW [7]);
  nor _85964_ (_36072_, _11533_, \oc8051_golden_model_1.PSW [7]);
  nor _85965_ (_36073_, _36072_, _11881_);
  not _85966_ (_36074_, _36073_);
  nor _85967_ (_36075_, _36074_, _36071_);
  nor _85968_ (_36076_, _36075_, _11885_);
  and _85969_ (_36077_, _36076_, _36070_);
  or _85970_ (_36078_, _36077_, _35854_);
  nand _85971_ (_36079_, _36078_, _08507_);
  nor _85972_ (_36081_, _11533_, _08507_);
  nor _85973_ (_36082_, _36081_, _08587_);
  and _85974_ (_36083_, _36082_, _36079_);
  and _85975_ (_36084_, _35852_, _08587_);
  or _85976_ (_36085_, _36084_, _03798_);
  nor _85977_ (_36086_, _36085_, _36083_);
  and _85978_ (_36087_, _05005_, _03798_);
  or _85979_ (_36088_, _36087_, _36086_);
  nand _85980_ (_36089_, _36088_, _06399_);
  and _85981_ (_36090_, _11534_, _03188_);
  nor _85982_ (_36092_, _36090_, _03621_);
  nand _85983_ (_36093_, _36092_, _36089_);
  and _85984_ (_36094_, _35865_, _09854_);
  nor _85985_ (_36095_, _11399_, _09854_);
  or _85986_ (_36096_, _36095_, _11903_);
  nor _85987_ (_36097_, _36096_, _36094_);
  nor _85988_ (_36098_, _36097_, _11907_);
  and _85989_ (_36099_, _36098_, _36093_);
  or _85990_ (_36100_, _36099_, _35853_);
  nand _85991_ (_36101_, _36100_, _08702_);
  nor _85992_ (_36103_, _11533_, _08702_);
  nor _85993_ (_36104_, _36103_, _08732_);
  and _85994_ (_36105_, _36104_, _36101_);
  and _85995_ (_36106_, _35852_, _08732_);
  or _85996_ (_36107_, _36106_, _03515_);
  nor _85997_ (_36108_, _36107_, _36105_);
  and _85998_ (_36109_, _05005_, _03515_);
  or _85999_ (_36110_, _36109_, _36108_);
  nand _86000_ (_36111_, _36110_, _32165_);
  and _86001_ (_36112_, _11534_, _03203_);
  nor _86002_ (_36114_, _36112_, _03628_);
  nand _86003_ (_36115_, _36114_, _36111_);
  nor _86004_ (_36116_, _35870_, _09854_);
  and _86005_ (_36117_, _11400_, _09854_);
  nor _86006_ (_36118_, _36117_, _36116_);
  and _86007_ (_36119_, _36118_, _03628_);
  nor _86008_ (_36120_, _36119_, _11934_);
  nand _86009_ (_36121_, _36120_, _36115_);
  nor _86010_ (_36122_, _35852_, _11933_);
  nor _86011_ (_36123_, _36122_, _03815_);
  nand _86012_ (_36125_, _36123_, _36121_);
  and _86013_ (_36126_, _11533_, _03815_);
  nor _86014_ (_36127_, _36126_, _32765_);
  nand _86015_ (_36128_, _36127_, _36125_);
  nor _86016_ (_36129_, _35852_, _11940_);
  nor _86017_ (_36130_, _36129_, _03629_);
  nand _86018_ (_36131_, _36130_, _36128_);
  nor _86019_ (_36132_, _11944_, _03581_);
  nor _86020_ (_36133_, _36132_, _03198_);
  nand _86021_ (_36134_, _36133_, _36131_);
  and _86022_ (_36136_, _11534_, _03198_);
  nor _86023_ (_36137_, _36136_, _03453_);
  nand _86024_ (_36138_, _36137_, _36134_);
  and _86025_ (_36139_, _36118_, _03453_);
  nor _86026_ (_36140_, _36139_, _11958_);
  nand _86027_ (_36141_, _36140_, _36138_);
  nor _86028_ (_36142_, _35852_, _11957_);
  nor _86029_ (_36143_, _36142_, _03447_);
  nand _86030_ (_36144_, _36143_, _36141_);
  and _86031_ (_36145_, _11533_, _03447_);
  nor _86032_ (_36147_, _36145_, _33825_);
  nand _86033_ (_36148_, _36147_, _36144_);
  nor _86034_ (_36149_, _35852_, _11964_);
  nor _86035_ (_36150_, _36149_, _03631_);
  nand _86036_ (_36151_, _36150_, _36148_);
  nor _86037_ (_36152_, _11968_, _03581_);
  nor _86038_ (_36153_, _36152_, _03196_);
  and _86039_ (_36154_, _36153_, _36151_);
  and _86040_ (_36155_, _11534_, _03196_);
  nor _86041_ (_36156_, _36155_, _36154_);
  and _86042_ (_36158_, _36156_, _11976_);
  and _86043_ (_36159_, _35852_, _11975_);
  or _86044_ (_36160_, _36159_, _36158_);
  or _86045_ (_36161_, _36160_, _43004_);
  or _86046_ (_36162_, _43000_, \oc8051_golden_model_1.PC [11]);
  and _86047_ (_36163_, _36162_, _41806_);
  and _86048_ (_43682_, _36163_, _36161_);
  and _86049_ (_36164_, _11525_, _08786_);
  and _86050_ (_36165_, _11611_, _11608_);
  nor _86051_ (_36166_, _36165_, _11612_);
  and _86052_ (_36168_, _36166_, _11826_);
  or _86053_ (_36169_, _36168_, _36164_);
  and _86054_ (_36170_, _36169_, _11819_);
  and _86055_ (_36171_, _11390_, _03222_);
  and _86056_ (_36172_, _11390_, _11685_);
  and _86057_ (_36173_, _11484_, _11481_);
  nor _86058_ (_36174_, _36173_, _11485_);
  and _86059_ (_36175_, _36174_, _10018_);
  or _86060_ (_36176_, _36175_, _36172_);
  nor _86061_ (_36177_, _36176_, _09920_);
  nor _86062_ (_36179_, _11321_, \oc8051_golden_model_1.PC [12]);
  nor _86063_ (_36180_, _36179_, _11322_);
  nor _86064_ (_36181_, _36180_, _11653_);
  not _86065_ (_36182_, _36180_);
  nor _86066_ (_36183_, _36182_, _11643_);
  not _86067_ (_36184_, _36183_);
  and _86068_ (_36185_, _11525_, _04409_);
  and _86069_ (_36186_, _09029_, \oc8051_golden_model_1.PC [12]);
  and _86070_ (_36187_, _36186_, _33169_);
  nor _86071_ (_36188_, _36187_, _36185_);
  not _86072_ (_36190_, _36188_);
  and _86073_ (_36191_, _36190_, _32816_);
  and _86074_ (_36192_, _11525_, _03980_);
  nor _86075_ (_36193_, _36192_, _06073_);
  not _86076_ (_36194_, _36193_);
  nor _86077_ (_36195_, _36194_, _36191_);
  and _86078_ (_36196_, _36195_, _36184_);
  and _86079_ (_36197_, _11504_, _11525_);
  and _86080_ (_36198_, _36166_, _11624_);
  or _86081_ (_36199_, _36198_, _36197_);
  nor _86082_ (_36201_, _36199_, _06072_);
  nor _86083_ (_36202_, _36201_, _36196_);
  nor _86084_ (_36203_, _36202_, _33523_);
  and _86085_ (_36204_, _11390_, _11369_);
  not _86086_ (_36205_, _36204_);
  and _86087_ (_36206_, _36174_, _11367_);
  nor _86088_ (_36207_, _36206_, _04081_);
  and _86089_ (_36208_, _36207_, _36205_);
  nor _86090_ (_36209_, _36208_, _36203_);
  nor _86091_ (_36210_, _36209_, _35265_);
  nor _86092_ (_36212_, _36210_, _36181_);
  nor _86093_ (_36213_, _36212_, _11652_);
  nor _86094_ (_36214_, _11360_, _11525_);
  nor _86095_ (_36215_, _36214_, _11660_);
  not _86096_ (_36216_, _36215_);
  nor _86097_ (_36217_, _36216_, _36213_);
  nor _86098_ (_36218_, _36182_, _11659_);
  nor _86099_ (_36219_, _36218_, _03729_);
  not _86100_ (_36220_, _36219_);
  nor _86101_ (_36221_, _36220_, _36217_);
  and _86102_ (_36223_, _11526_, _03729_);
  nor _86103_ (_36224_, _36223_, _11668_);
  not _86104_ (_36225_, _36224_);
  or _86105_ (_36226_, _36225_, _36221_);
  nor _86106_ (_36227_, _36182_, _11666_);
  nor _86107_ (_36228_, _36227_, _11673_);
  and _86108_ (_36229_, _36228_, _36226_);
  nor _86109_ (_36230_, _11672_, _11525_);
  or _86110_ (_36231_, _36230_, _09917_);
  or _86111_ (_36232_, _36231_, _36229_);
  and _86112_ (_36234_, _11391_, _09969_);
  nor _86113_ (_36235_, _36174_, _09969_);
  or _86114_ (_36236_, _36235_, _09921_);
  or _86115_ (_36237_, _36236_, _36234_);
  and _86116_ (_36238_, _36237_, _09920_);
  and _86117_ (_36239_, _36238_, _36232_);
  or _86118_ (_36240_, _36239_, _03615_);
  or _86119_ (_36241_, _36240_, _36177_);
  and _86120_ (_36242_, _36174_, _11693_);
  and _86121_ (_36243_, _11390_, _09876_);
  nor _86122_ (_36245_, _36243_, _36242_);
  nor _86123_ (_36246_, _36245_, _04107_);
  nor _86124_ (_36247_, _36246_, _03604_);
  and _86125_ (_36248_, _36247_, _36241_);
  nor _86126_ (_36249_, _36174_, _10061_);
  and _86127_ (_36250_, _11391_, _10061_);
  nor _86128_ (_36251_, _36250_, _36249_);
  nor _86129_ (_36252_, _36251_, _09856_);
  nor _86130_ (_36253_, _36252_, _10025_);
  not _86131_ (_36254_, _36253_);
  or _86132_ (_36256_, _36254_, _36248_);
  and _86133_ (_36257_, _36180_, _10025_);
  not _86134_ (_36258_, _36257_);
  and _86135_ (_36259_, _36258_, _11720_);
  nand _86136_ (_36260_, _36259_, _36256_);
  nor _86137_ (_36261_, _11720_, _11525_);
  nor _86138_ (_36262_, _36261_, _11356_);
  nand _86139_ (_36263_, _36262_, _36260_);
  nor _86140_ (_36264_, _36182_, _11355_);
  nor _86141_ (_36265_, _36264_, _35954_);
  nand _86142_ (_36267_, _36265_, _36263_);
  nor _86143_ (_36268_, _11729_, _11525_);
  not _86144_ (_36269_, _36268_);
  and _86145_ (_36270_, _36269_, _11350_);
  nand _86146_ (_36271_, _36270_, _36267_);
  nor _86147_ (_36272_, _36182_, _11350_);
  nor _86148_ (_36273_, _36272_, _08187_);
  nand _86149_ (_36274_, _36273_, _36271_);
  nor _86150_ (_36275_, _11525_, _08186_);
  nor _86151_ (_36276_, _36275_, _07912_);
  nand _86152_ (_36278_, _36276_, _36274_);
  nor _86153_ (_36279_, _36182_, _03248_);
  nor _86154_ (_36280_, _36279_, _11741_);
  nand _86155_ (_36281_, _36280_, _36278_);
  nor _86156_ (_36282_, _11740_, _11525_);
  nor _86157_ (_36283_, _36282_, _03625_);
  nand _86158_ (_36284_, _36283_, _36281_);
  and _86159_ (_36285_, _11390_, _03625_);
  nor _86160_ (_36286_, _36285_, _33299_);
  nand _86161_ (_36287_, _36286_, _36284_);
  nor _86162_ (_36289_, _11749_, _11525_);
  nor _86163_ (_36290_, _36289_, _03222_);
  and _86164_ (_36291_, _36290_, _36287_);
  or _86165_ (_36292_, _36291_, _36171_);
  nand _86166_ (_36293_, _36292_, _11756_);
  nor _86167_ (_36294_, _36182_, _11756_);
  nor _86168_ (_36295_, _36294_, _11761_);
  nand _86169_ (_36296_, _36295_, _36293_);
  nor _86170_ (_36297_, _11760_, _11525_);
  nor _86171_ (_36298_, _36297_, _11764_);
  nand _86172_ (_36300_, _36298_, _36296_);
  and _86173_ (_36301_, _36166_, _11764_);
  nor _86174_ (_36302_, _36301_, _06168_);
  and _86175_ (_36303_, _36302_, _36300_);
  nor _86176_ (_36304_, _11526_, _03601_);
  nor _86177_ (_36305_, _36304_, _05895_);
  or _86178_ (_36306_, _36305_, _36303_);
  and _86179_ (_36307_, _11390_, _03601_);
  nor _86180_ (_36308_, _36307_, _08363_);
  nand _86181_ (_36309_, _36308_, _36306_);
  and _86182_ (_36311_, _11526_, _08363_);
  nor _86183_ (_36312_, _36311_, _11347_);
  nand _86184_ (_36313_, _36312_, _36309_);
  nor _86185_ (_36314_, _11807_, \oc8051_golden_model_1.DPH [4]);
  nor _86186_ (_36315_, _36314_, _11808_);
  and _86187_ (_36316_, _36315_, _11347_);
  nor _86188_ (_36317_, _36316_, _11816_);
  nand _86189_ (_36318_, _36317_, _36313_);
  nor _86190_ (_36319_, _11815_, _11525_);
  nor _86191_ (_36320_, _36319_, _11819_);
  and _86192_ (_36322_, _36320_, _36318_);
  or _86193_ (_36323_, _36322_, _36170_);
  nand _86194_ (_36324_, _36323_, _11345_);
  nor _86195_ (_36325_, _36182_, _11345_);
  nor _86196_ (_36326_, _36325_, _11342_);
  nand _86197_ (_36327_, _36326_, _36324_);
  nor _86198_ (_36328_, _11525_, _11341_);
  nor _86199_ (_36329_, _36328_, _03600_);
  nand _86200_ (_36330_, _36329_, _36327_);
  and _86201_ (_36331_, _11390_, _03600_);
  nor _86202_ (_36333_, _36331_, _36024_);
  nand _86203_ (_36334_, _36333_, _36330_);
  nor _86204_ (_36335_, _11838_, _11525_);
  nor _86205_ (_36336_, _36335_, _11841_);
  nand _86206_ (_36337_, _36336_, _36334_);
  nand _86207_ (_36338_, _11525_, _11826_);
  nand _86208_ (_36339_, _36166_, _08786_);
  and _86209_ (_36340_, _36339_, _36338_);
  or _86210_ (_36341_, _36340_, _11842_);
  nand _86211_ (_36342_, _36341_, _36337_);
  nand _86212_ (_36344_, _36342_, _11851_);
  nor _86213_ (_36345_, _36182_, _11851_);
  nor _86214_ (_36346_, _36345_, _08431_);
  nand _86215_ (_36347_, _36346_, _36344_);
  nor _86216_ (_36348_, _11525_, _08430_);
  nor _86217_ (_36349_, _36348_, _03622_);
  nand _86218_ (_36350_, _36349_, _36347_);
  and _86219_ (_36351_, _11390_, _03622_);
  nor _86220_ (_36352_, _36351_, _10754_);
  and _86221_ (_36353_, _36352_, _36350_);
  nor _86222_ (_36355_, _11526_, _11337_);
  nor _86223_ (_36356_, _36355_, _24116_);
  nor _86224_ (_36357_, _36356_, _36353_);
  and _86225_ (_36358_, _11525_, \oc8051_golden_model_1.PSW [7]);
  and _86226_ (_36359_, _36166_, _07871_);
  or _86227_ (_36360_, _36359_, _36358_);
  and _86228_ (_36361_, _36360_, _11337_);
  or _86229_ (_36362_, _36361_, _36357_);
  nand _86230_ (_36363_, _36362_, _11335_);
  nor _86231_ (_36364_, _36182_, _11335_);
  nor _86232_ (_36366_, _36364_, _08460_);
  nand _86233_ (_36367_, _36366_, _36363_);
  nor _86234_ (_36368_, _11525_, _08459_);
  nor _86235_ (_36369_, _36368_, _03624_);
  nand _86236_ (_36370_, _36369_, _36367_);
  and _86237_ (_36371_, _11390_, _03624_);
  nor _86238_ (_36372_, _36371_, _36063_);
  and _86239_ (_36373_, _36372_, _36370_);
  nor _86240_ (_36374_, _11880_, _11526_);
  nor _86241_ (_36375_, _36374_, _24239_);
  or _86242_ (_36377_, _36375_, _36373_);
  nand _86243_ (_36378_, _11525_, _07871_);
  nand _86244_ (_36379_, _36166_, \oc8051_golden_model_1.PSW [7]);
  and _86245_ (_36380_, _36379_, _36378_);
  or _86246_ (_36381_, _36380_, _11881_);
  nand _86247_ (_36382_, _36381_, _36377_);
  nand _86248_ (_36383_, _36382_, _11330_);
  nor _86249_ (_36384_, _36182_, _11330_);
  nor _86250_ (_36385_, _36384_, _08508_);
  nand _86251_ (_36386_, _36385_, _36383_);
  nor _86252_ (_36388_, _11525_, _08507_);
  nor _86253_ (_36389_, _36388_, _08587_);
  and _86254_ (_36390_, _36389_, _36386_);
  and _86255_ (_36391_, _36180_, _08587_);
  or _86256_ (_36392_, _36391_, _03798_);
  nor _86257_ (_36393_, _36392_, _36390_);
  and _86258_ (_36394_, _05777_, _03798_);
  or _86259_ (_36395_, _36394_, _36393_);
  nand _86260_ (_36396_, _36395_, _06399_);
  and _86261_ (_36397_, _11526_, _03188_);
  nor _86262_ (_36399_, _36397_, _03621_);
  and _86263_ (_36400_, _36399_, _36396_);
  and _86264_ (_36401_, _36174_, _09854_);
  nor _86265_ (_36402_, _11391_, _09854_);
  nor _86266_ (_36403_, _36402_, _36401_);
  nor _86267_ (_36404_, _36403_, _11903_);
  or _86268_ (_36405_, _36404_, _36400_);
  nand _86269_ (_36406_, _36405_, _11328_);
  nor _86270_ (_36407_, _36182_, _11328_);
  nor _86271_ (_36408_, _36407_, _08703_);
  nand _86272_ (_36410_, _36408_, _36406_);
  nor _86273_ (_36411_, _11525_, _08702_);
  nor _86274_ (_36412_, _36411_, _08732_);
  nand _86275_ (_36413_, _36412_, _36410_);
  and _86276_ (_36414_, _36180_, _08732_);
  nor _86277_ (_36415_, _36414_, _03515_);
  nand _86278_ (_36416_, _36415_, _36413_);
  and _86279_ (_36417_, _05777_, _03515_);
  nor _86280_ (_36418_, _36417_, _03203_);
  and _86281_ (_36419_, _36418_, _36416_);
  and _86282_ (_36421_, _11525_, _03203_);
  or _86283_ (_36422_, _36421_, _03628_);
  or _86284_ (_36423_, _36422_, _36419_);
  nor _86285_ (_36424_, _36174_, _09854_);
  and _86286_ (_36425_, _11391_, _09854_);
  nor _86287_ (_36426_, _36425_, _36424_);
  nor _86288_ (_36427_, _36426_, _03816_);
  nor _86289_ (_36428_, _36427_, _11934_);
  nand _86290_ (_36429_, _36428_, _36423_);
  nor _86291_ (_36430_, _36182_, _11933_);
  nor _86292_ (_36432_, _36430_, _03815_);
  nand _86293_ (_36433_, _36432_, _36429_);
  and _86294_ (_36434_, _11526_, _03815_);
  nor _86295_ (_36435_, _36434_, _32765_);
  nand _86296_ (_36436_, _36435_, _36433_);
  nor _86297_ (_36437_, _36182_, _11940_);
  nor _86298_ (_36438_, _36437_, _03629_);
  nand _86299_ (_36439_, _36438_, _36436_);
  and _86300_ (_36440_, _03486_, _03629_);
  nor _86301_ (_36441_, _36440_, _03198_);
  and _86302_ (_36443_, _36441_, _36439_);
  and _86303_ (_36444_, _11525_, _03198_);
  or _86304_ (_36445_, _36444_, _03453_);
  or _86305_ (_36446_, _36445_, _36443_);
  nor _86306_ (_36447_, _36426_, _03823_);
  nor _86307_ (_36448_, _36447_, _11958_);
  nand _86308_ (_36449_, _36448_, _36446_);
  nor _86309_ (_36450_, _36182_, _11957_);
  nor _86310_ (_36451_, _36450_, _03447_);
  nand _86311_ (_36452_, _36451_, _36449_);
  and _86312_ (_36454_, _11526_, _03447_);
  nor _86313_ (_36455_, _36454_, _33825_);
  nand _86314_ (_36456_, _36455_, _36452_);
  nor _86315_ (_36457_, _36182_, _11964_);
  nor _86316_ (_36458_, _36457_, _03631_);
  nand _86317_ (_36459_, _36458_, _36456_);
  and _86318_ (_36460_, _03486_, _03631_);
  nor _86319_ (_36461_, _36460_, _03196_);
  nand _86320_ (_36462_, _36461_, _36459_);
  and _86321_ (_36463_, _11525_, _03196_);
  nor _86322_ (_36465_, _36463_, _11975_);
  and _86323_ (_36466_, _36465_, _36462_);
  and _86324_ (_36467_, _36182_, _11975_);
  nor _86325_ (_36468_, _36467_, _36466_);
  or _86326_ (_36469_, _36468_, _43004_);
  or _86327_ (_36470_, _43000_, \oc8051_golden_model_1.PC [12]);
  and _86328_ (_36471_, _36470_, _41806_);
  and _86329_ (_43683_, _36471_, _36469_);
  nor _86330_ (_36472_, _11322_, \oc8051_golden_model_1.PC [13]);
  nor _86331_ (_36473_, _36472_, _11323_);
  or _86332_ (_36475_, _36473_, _11328_);
  or _86333_ (_36476_, _36473_, _11330_);
  or _86334_ (_36477_, _36473_, _11335_);
  or _86335_ (_36478_, _11523_, _11522_);
  not _86336_ (_36479_, _36478_);
  nor _86337_ (_36480_, _36479_, _11613_);
  and _86338_ (_36481_, _36479_, _11613_);
  or _86339_ (_36482_, _36481_, _36480_);
  or _86340_ (_36483_, _36482_, _08786_);
  or _86341_ (_36484_, _11521_, _11826_);
  and _86342_ (_36486_, _36484_, _11819_);
  and _86343_ (_36487_, _36486_, _36483_);
  or _86344_ (_36488_, _11521_, _05894_);
  and _86345_ (_36489_, _11385_, _03222_);
  or _86346_ (_36490_, _36473_, _11350_);
  and _86347_ (_36491_, _36473_, _11356_);
  or _86348_ (_36492_, _11388_, _11387_);
  not _86349_ (_36493_, _36492_);
  nor _86350_ (_36494_, _36493_, _11486_);
  and _86351_ (_36495_, _36493_, _11486_);
  or _86352_ (_36497_, _36495_, _36494_);
  or _86353_ (_36498_, _36497_, _10061_);
  nand _86354_ (_36499_, _11386_, _10061_);
  and _86355_ (_36500_, _36499_, _03604_);
  and _86356_ (_36501_, _36500_, _36498_);
  and _86357_ (_36502_, _36497_, _10018_);
  and _86358_ (_36503_, _11385_, _11685_);
  or _86359_ (_36504_, _36503_, _36502_);
  or _86360_ (_36505_, _36504_, _09920_);
  and _86361_ (_36506_, _11521_, _03729_);
  or _86362_ (_36508_, _11360_, _11521_);
  or _86363_ (_36509_, _36497_, _11369_);
  or _86364_ (_36510_, _11385_, _11367_);
  and _86365_ (_36511_, _36510_, _03610_);
  and _86366_ (_36512_, _36511_, _36509_);
  and _86367_ (_36513_, _36482_, _11624_);
  and _86368_ (_36514_, _11504_, _11521_);
  or _86369_ (_36515_, _36514_, _06072_);
  or _86370_ (_36516_, _36515_, _36513_);
  or _86371_ (_36517_, _36473_, _11643_);
  or _86372_ (_36519_, _11521_, _04763_);
  or _86373_ (_36520_, _11521_, _35582_);
  or _86374_ (_36521_, _04409_, \oc8051_golden_model_1.PC [13]);
  or _86375_ (_36522_, _36521_, _04729_);
  nand _86376_ (_36523_, _36522_, _36520_);
  nand _86377_ (_36524_, _36523_, _32816_);
  and _86378_ (_36525_, _36524_, _36519_);
  and _86379_ (_36526_, _36525_, _36517_);
  or _86380_ (_36527_, _36526_, _06073_);
  and _86381_ (_36528_, _36527_, _11647_);
  and _86382_ (_36530_, _36528_, _36516_);
  or _86383_ (_36531_, _36530_, _36512_);
  and _86384_ (_36532_, _36531_, _11362_);
  and _86385_ (_36533_, _36473_, _11654_);
  or _86386_ (_36534_, _36533_, _11652_);
  or _86387_ (_36535_, _36534_, _36532_);
  and _86388_ (_36536_, _36535_, _36508_);
  or _86389_ (_36537_, _36536_, _11660_);
  or _86390_ (_36538_, _36473_, _11659_);
  and _86391_ (_36539_, _36538_, _03737_);
  and _86392_ (_36541_, _36539_, _36537_);
  or _86393_ (_36542_, _36541_, _36506_);
  and _86394_ (_36543_, _36542_, _11666_);
  and _86395_ (_36544_, _36473_, _11668_);
  or _86396_ (_36545_, _36544_, _11673_);
  or _86397_ (_36546_, _36545_, _36543_);
  or _86398_ (_36547_, _11672_, _11521_);
  and _86399_ (_36548_, _36547_, _09921_);
  and _86400_ (_36549_, _36548_, _36546_);
  or _86401_ (_36550_, _36497_, _09969_);
  nand _86402_ (_36552_, _11386_, _09969_);
  and _86403_ (_36553_, _36552_, _09917_);
  and _86404_ (_36554_, _36553_, _36550_);
  or _86405_ (_36555_, _36554_, _09919_);
  or _86406_ (_36556_, _36555_, _36549_);
  and _86407_ (_36557_, _36556_, _36505_);
  or _86408_ (_36558_, _36557_, _03615_);
  and _86409_ (_36559_, _36497_, _11693_);
  and _86410_ (_36560_, _11385_, _09876_);
  or _86411_ (_36561_, _36560_, _04107_);
  or _86412_ (_36563_, _36561_, _36559_);
  and _86413_ (_36564_, _36563_, _09856_);
  and _86414_ (_36565_, _36564_, _36558_);
  or _86415_ (_36566_, _36565_, _36501_);
  and _86416_ (_36567_, _36566_, _11358_);
  nand _86417_ (_36568_, _36473_, _10025_);
  nand _86418_ (_36569_, _36568_, _11720_);
  or _86419_ (_36570_, _36569_, _36567_);
  or _86420_ (_36571_, _11720_, _11521_);
  and _86421_ (_36572_, _36571_, _11355_);
  and _86422_ (_36574_, _36572_, _36570_);
  or _86423_ (_36575_, _36574_, _36491_);
  and _86424_ (_36576_, _36575_, _11729_);
  nand _86425_ (_36577_, _35954_, _11521_);
  nand _86426_ (_36578_, _36577_, _11350_);
  or _86427_ (_36579_, _36578_, _36576_);
  and _86428_ (_36580_, _36579_, _36490_);
  or _86429_ (_36581_, _36580_, _08187_);
  or _86430_ (_36582_, _11521_, _08186_);
  and _86431_ (_36583_, _36582_, _03248_);
  and _86432_ (_36585_, _36583_, _36581_);
  nand _86433_ (_36586_, _36473_, _07912_);
  nand _86434_ (_36587_, _36586_, _11740_);
  or _86435_ (_36588_, _36587_, _36585_);
  or _86436_ (_36589_, _11740_, _11521_);
  and _86437_ (_36590_, _36589_, _08832_);
  and _86438_ (_36591_, _36590_, _36588_);
  nand _86439_ (_36592_, _11385_, _03625_);
  nand _86440_ (_36593_, _36592_, _11749_);
  or _86441_ (_36594_, _36593_, _36591_);
  or _86442_ (_36596_, _11749_, _11521_);
  and _86443_ (_36597_, _36596_, _03589_);
  and _86444_ (_36598_, _36597_, _36594_);
  or _86445_ (_36599_, _36598_, _36489_);
  and _86446_ (_36600_, _36599_, _11756_);
  and _86447_ (_36601_, _36473_, _11758_);
  or _86448_ (_36602_, _36601_, _11761_);
  or _86449_ (_36603_, _36602_, _36600_);
  or _86450_ (_36604_, _11760_, _11521_);
  and _86451_ (_36605_, _36604_, _11765_);
  and _86452_ (_36607_, _36605_, _36603_);
  and _86453_ (_36608_, _36482_, _11764_);
  or _86454_ (_36609_, _36608_, _06168_);
  or _86455_ (_36610_, _36609_, _36607_);
  and _86456_ (_36611_, _36610_, _36488_);
  or _86457_ (_36612_, _36611_, _03601_);
  or _86458_ (_36613_, _11385_, _05886_);
  and _86459_ (_36614_, _36613_, _08364_);
  and _86460_ (_36615_, _36614_, _36612_);
  and _86461_ (_36616_, _11521_, _08363_);
  or _86462_ (_36618_, _36616_, _36615_);
  and _86463_ (_36619_, _36618_, _11348_);
  or _86464_ (_36620_, _11808_, \oc8051_golden_model_1.DPH [5]);
  nor _86465_ (_36621_, _11809_, _11348_);
  and _86466_ (_36622_, _36621_, _36620_);
  or _86467_ (_36623_, _36622_, _11816_);
  or _86468_ (_36624_, _36623_, _36619_);
  or _86469_ (_36625_, _11815_, _11521_);
  and _86470_ (_36626_, _36625_, _11820_);
  and _86471_ (_36627_, _36626_, _36624_);
  or _86472_ (_36629_, _36627_, _36487_);
  and _86473_ (_36630_, _36629_, _11345_);
  and _86474_ (_36631_, _36473_, _11824_);
  or _86475_ (_36632_, _36631_, _11342_);
  or _86476_ (_36633_, _36632_, _36630_);
  or _86477_ (_36634_, _11521_, _11341_);
  and _86478_ (_36635_, _36634_, _07766_);
  and _86479_ (_36636_, _36635_, _36633_);
  nand _86480_ (_36637_, _11385_, _03600_);
  nand _86481_ (_36638_, _36637_, _11838_);
  or _86482_ (_36640_, _36638_, _36636_);
  or _86483_ (_36641_, _11838_, _11521_);
  and _86484_ (_36642_, _36641_, _11842_);
  and _86485_ (_36643_, _36642_, _36640_);
  or _86486_ (_36644_, _36482_, _11826_);
  or _86487_ (_36645_, _11521_, _08786_);
  and _86488_ (_36646_, _36645_, _11841_);
  and _86489_ (_36647_, _36646_, _36644_);
  or _86490_ (_36648_, _36647_, _36643_);
  and _86491_ (_36649_, _36648_, _11851_);
  and _86492_ (_36651_, _36473_, _11853_);
  or _86493_ (_36652_, _36651_, _08431_);
  or _86494_ (_36653_, _36652_, _36649_);
  or _86495_ (_36654_, _11521_, _08430_);
  and _86496_ (_36655_, _36654_, _07777_);
  and _86497_ (_36656_, _36655_, _36653_);
  nand _86498_ (_36657_, _11385_, _03622_);
  nand _86499_ (_36658_, _36657_, _10753_);
  or _86500_ (_36659_, _36658_, _36656_);
  and _86501_ (_36660_, _11521_, _11338_);
  or _86502_ (_36662_, _36660_, _24116_);
  and _86503_ (_36663_, _36662_, _36659_);
  or _86504_ (_36664_, _36482_, \oc8051_golden_model_1.PSW [7]);
  or _86505_ (_36665_, _11521_, _07871_);
  and _86506_ (_36666_, _36665_, _11337_);
  and _86507_ (_36667_, _36666_, _36664_);
  or _86508_ (_36668_, _36667_, _11864_);
  or _86509_ (_36669_, _36668_, _36663_);
  and _86510_ (_36670_, _36669_, _36477_);
  or _86511_ (_36671_, _36670_, _08460_);
  or _86512_ (_36673_, _11521_, _08459_);
  and _86513_ (_36674_, _36673_, _07795_);
  and _86514_ (_36675_, _36674_, _36671_);
  nand _86515_ (_36676_, _11385_, _03624_);
  nand _86516_ (_36677_, _36676_, _11877_);
  or _86517_ (_36678_, _36677_, _36675_);
  and _86518_ (_36679_, _11881_, _11521_);
  or _86519_ (_36680_, _36679_, _24239_);
  and _86520_ (_36681_, _36680_, _36678_);
  or _86521_ (_36682_, _36482_, _07871_);
  or _86522_ (_36684_, _11521_, \oc8051_golden_model_1.PSW [7]);
  and _86523_ (_36685_, _36684_, _11880_);
  and _86524_ (_36686_, _36685_, _36682_);
  or _86525_ (_36687_, _36686_, _11885_);
  or _86526_ (_36688_, _36687_, _36681_);
  and _86527_ (_36689_, _36688_, _36476_);
  or _86528_ (_36690_, _36689_, _08508_);
  or _86529_ (_36691_, _11521_, _08507_);
  and _86530_ (_36692_, _36691_, _08588_);
  and _86531_ (_36693_, _36692_, _36690_);
  and _86532_ (_36695_, _36473_, _08587_);
  or _86533_ (_36696_, _36695_, _03798_);
  or _86534_ (_36697_, _36696_, _36693_);
  nand _86535_ (_36698_, _05469_, _03798_);
  and _86536_ (_36699_, _36698_, _36697_);
  or _86537_ (_36700_, _36699_, _03188_);
  or _86538_ (_36701_, _11521_, _06399_);
  and _86539_ (_36702_, _36701_, _11903_);
  and _86540_ (_36703_, _36702_, _36700_);
  or _86541_ (_36704_, _36497_, _11908_);
  or _86542_ (_36706_, _11385_, _09854_);
  and _86543_ (_36707_, _36706_, _03621_);
  and _86544_ (_36708_, _36707_, _36704_);
  or _86545_ (_36709_, _36708_, _11907_);
  or _86546_ (_36710_, _36709_, _36703_);
  and _86547_ (_36711_, _36710_, _36475_);
  or _86548_ (_36712_, _36711_, _08703_);
  or _86549_ (_36713_, _11521_, _08702_);
  and _86550_ (_36714_, _36713_, _08733_);
  and _86551_ (_36715_, _36714_, _36712_);
  and _86552_ (_36717_, _36473_, _08732_);
  or _86553_ (_36718_, _36717_, _03515_);
  or _86554_ (_36719_, _36718_, _36715_);
  nand _86555_ (_36720_, _05469_, _03515_);
  and _86556_ (_36721_, _36720_, _36719_);
  or _86557_ (_36722_, _36721_, _03203_);
  or _86558_ (_36723_, _11521_, _32165_);
  and _86559_ (_36724_, _36723_, _03816_);
  and _86560_ (_36725_, _36724_, _36722_);
  nand _86561_ (_36726_, _11386_, _09854_);
  or _86562_ (_36728_, _36497_, _09854_);
  and _86563_ (_36729_, _36728_, _36726_);
  and _86564_ (_36730_, _36729_, _03628_);
  or _86565_ (_36731_, _36730_, _11934_);
  or _86566_ (_36732_, _36731_, _36725_);
  or _86567_ (_36733_, _36473_, _11933_);
  and _86568_ (_36734_, _36733_, _04246_);
  and _86569_ (_36735_, _36734_, _36732_);
  nand _86570_ (_36736_, _11521_, _03815_);
  nand _86571_ (_36737_, _36736_, _11940_);
  or _86572_ (_36739_, _36737_, _36735_);
  or _86573_ (_36740_, _36473_, _11940_);
  and _86574_ (_36741_, _36740_, _11944_);
  and _86575_ (_36742_, _36741_, _36739_);
  nor _86576_ (_36743_, _03860_, _11944_);
  or _86577_ (_36744_, _36743_, _03198_);
  or _86578_ (_36745_, _36744_, _36742_);
  or _86579_ (_36746_, _11521_, _12371_);
  and _86580_ (_36747_, _36746_, _03823_);
  and _86581_ (_36748_, _36747_, _36745_);
  and _86582_ (_36750_, _36729_, _03453_);
  or _86583_ (_36751_, _36750_, _11958_);
  or _86584_ (_36752_, _36751_, _36748_);
  or _86585_ (_36753_, _36473_, _11957_);
  and _86586_ (_36754_, _36753_, _03514_);
  and _86587_ (_36755_, _36754_, _36752_);
  nand _86588_ (_36756_, _11521_, _03447_);
  nand _86589_ (_36757_, _36756_, _11964_);
  or _86590_ (_36758_, _36757_, _36755_);
  or _86591_ (_36759_, _36473_, _11964_);
  and _86592_ (_36761_, _36759_, _11968_);
  and _86593_ (_36762_, _36761_, _36758_);
  nor _86594_ (_36763_, _03860_, _11968_);
  or _86595_ (_36764_, _36763_, _03196_);
  or _86596_ (_36765_, _36764_, _36762_);
  not _86597_ (_36766_, _11521_);
  nand _86598_ (_36767_, _36766_, _03196_);
  and _86599_ (_36768_, _36767_, _11976_);
  and _86600_ (_36769_, _36768_, _36765_);
  and _86601_ (_36770_, _36473_, _11975_);
  or _86602_ (_36772_, _36770_, _36769_);
  or _86603_ (_36773_, _36772_, _43004_);
  or _86604_ (_36774_, _43000_, \oc8051_golden_model_1.PC [13]);
  and _86605_ (_36775_, _36774_, _41806_);
  and _86606_ (_43684_, _36775_, _36773_);
  nor _86607_ (_36776_, _11323_, \oc8051_golden_model_1.PC [14]);
  nor _86608_ (_36777_, _36776_, _11324_);
  nor _86609_ (_36778_, _36777_, _08733_);
  nor _86610_ (_36779_, _11877_, _11515_);
  nor _86611_ (_36780_, _11515_, _10753_);
  nor _86612_ (_36782_, _11838_, _11515_);
  nor _86613_ (_36783_, _11815_, _11515_);
  and _86614_ (_36784_, _11488_, _11383_);
  nor _86615_ (_36785_, _36784_, _11489_);
  or _86616_ (_36786_, _36785_, _11685_);
  or _86617_ (_36787_, _11378_, _10018_);
  and _86618_ (_36788_, _36787_, _09919_);
  and _86619_ (_36789_, _36788_, _36786_);
  and _86620_ (_36790_, _36777_, _11668_);
  nor _86621_ (_36791_, _36777_, _11659_);
  or _86622_ (_36793_, _36785_, _11369_);
  or _86623_ (_36794_, _11378_, _11367_);
  and _86624_ (_36795_, _36794_, _36793_);
  nor _86625_ (_36796_, _36795_, _04081_);
  and _86626_ (_36797_, _11615_, _11519_);
  nor _86627_ (_36798_, _36797_, _11616_);
  nand _86628_ (_36799_, _36798_, _11624_);
  or _86629_ (_36800_, _11624_, _11515_);
  and _86630_ (_36801_, _36800_, _06073_);
  nand _86631_ (_36802_, _36801_, _36799_);
  nor _86632_ (_36804_, _36777_, _11642_);
  nor _86633_ (_36805_, _11632_, \oc8051_golden_model_1.PC [14]);
  and _86634_ (_36806_, _36805_, _09029_);
  and _86635_ (_36807_, _36806_, _33169_);
  nor _86636_ (_36808_, _36807_, _36804_);
  nor _86637_ (_36809_, _36808_, _03980_);
  not _86638_ (_36810_, _36809_);
  nor _86639_ (_36811_, _03980_, _04409_);
  nor _86640_ (_36812_, _36811_, _11514_);
  nor _86641_ (_36813_, _36812_, _11631_);
  and _86642_ (_36815_, _36813_, _36810_);
  not _86643_ (_36816_, _36777_);
  nor _86644_ (_36817_, _36816_, _11630_);
  nor _86645_ (_36818_, _36817_, _06073_);
  not _86646_ (_36819_, _36818_);
  nor _86647_ (_36820_, _36819_, _36815_);
  nor _86648_ (_36821_, _36820_, _04422_);
  nand _86649_ (_36822_, _36821_, _36802_);
  and _86650_ (_36823_, _36777_, _04422_);
  nor _86651_ (_36824_, _36823_, _03610_);
  and _86652_ (_36826_, _36824_, _36822_);
  or _86653_ (_36827_, _36826_, _36796_);
  nand _86654_ (_36828_, _36827_, _11362_);
  nor _86655_ (_36829_, _36777_, _11362_);
  nor _86656_ (_36830_, _36829_, _11652_);
  nand _86657_ (_36831_, _36830_, _36828_);
  nor _86658_ (_36832_, _11360_, _11515_);
  nor _86659_ (_36833_, _36832_, _11660_);
  and _86660_ (_36834_, _36833_, _36831_);
  or _86661_ (_36835_, _36834_, _36791_);
  nand _86662_ (_36837_, _36835_, _03737_);
  nor _86663_ (_36838_, _11514_, _03737_);
  nor _86664_ (_36839_, _36838_, _11668_);
  and _86665_ (_36840_, _36839_, _36837_);
  or _86666_ (_36841_, _36840_, _36790_);
  nand _86667_ (_36842_, _36841_, _11672_);
  nor _86668_ (_36843_, _11672_, _11515_);
  nor _86669_ (_36844_, _36843_, _09917_);
  nand _86670_ (_36845_, _36844_, _36842_);
  and _86671_ (_36846_, _11378_, _09969_);
  not _86672_ (_36848_, _36785_);
  nor _86673_ (_36849_, _36848_, _09969_);
  or _86674_ (_36850_, _36849_, _36846_);
  nor _86675_ (_36851_, _36850_, _09921_);
  nor _86676_ (_36852_, _36851_, _09919_);
  and _86677_ (_36853_, _36852_, _36845_);
  or _86678_ (_36854_, _36853_, _03615_);
  or _86679_ (_36855_, _36854_, _36789_);
  and _86680_ (_36856_, _11378_, _09876_);
  nor _86681_ (_36857_, _36848_, _09876_);
  or _86682_ (_36859_, _36857_, _04107_);
  or _86683_ (_36860_, _36859_, _36856_);
  and _86684_ (_36861_, _36860_, _09856_);
  nand _86685_ (_36862_, _36861_, _36855_);
  and _86686_ (_36863_, _11379_, _10061_);
  nor _86687_ (_36864_, _36785_, _10061_);
  or _86688_ (_36865_, _36864_, _09856_);
  or _86689_ (_36866_, _36865_, _36863_);
  and _86690_ (_36867_, _36866_, _11358_);
  and _86691_ (_36868_, _36867_, _36862_);
  nor _86692_ (_36870_, _36777_, _11358_);
  or _86693_ (_36871_, _36870_, _36868_);
  and _86694_ (_36872_, _36871_, _11720_);
  nor _86695_ (_36873_, _11720_, _11514_);
  or _86696_ (_36874_, _36873_, _36872_);
  nand _86697_ (_36875_, _36874_, _11355_);
  nor _86698_ (_36876_, _36777_, _11355_);
  nor _86699_ (_36877_, _36876_, _35954_);
  and _86700_ (_36878_, _36877_, _36875_);
  nor _86701_ (_36879_, _11729_, _11515_);
  nor _86702_ (_36881_, _36879_, _36878_);
  nand _86703_ (_36882_, _36881_, _11350_);
  nor _86704_ (_36883_, _36777_, _11350_);
  nor _86705_ (_36884_, _36883_, _08187_);
  nand _86706_ (_36885_, _36884_, _36882_);
  nor _86707_ (_36886_, _11515_, _08186_);
  nor _86708_ (_36887_, _36886_, _07912_);
  nand _86709_ (_36888_, _36887_, _36885_);
  nor _86710_ (_36889_, _36777_, _03248_);
  nor _86711_ (_36890_, _36889_, _11741_);
  nand _86712_ (_36892_, _36890_, _36888_);
  nor _86713_ (_36893_, _11740_, _11515_);
  nor _86714_ (_36894_, _36893_, _03625_);
  nand _86715_ (_36895_, _36894_, _36892_);
  nor _86716_ (_36896_, _11378_, _08832_);
  nor _86717_ (_36897_, _36896_, _33299_);
  nand _86718_ (_36898_, _36897_, _36895_);
  nor _86719_ (_36899_, _11749_, _11515_);
  nor _86720_ (_36900_, _36899_, _03222_);
  nand _86721_ (_36901_, _36900_, _36898_);
  nor _86722_ (_36903_, _11378_, _03589_);
  nor _86723_ (_36904_, _36903_, _11758_);
  nand _86724_ (_36905_, _36904_, _36901_);
  and _86725_ (_36906_, _36777_, _11758_);
  nor _86726_ (_36907_, _36906_, _11761_);
  nand _86727_ (_36908_, _36907_, _36905_);
  nor _86728_ (_36909_, _11760_, _11514_);
  nor _86729_ (_36910_, _36909_, _11764_);
  and _86730_ (_36911_, _36910_, _36908_);
  and _86731_ (_36912_, _36798_, _11764_);
  nor _86732_ (_36914_, _36912_, _36911_);
  or _86733_ (_36915_, _36914_, _06168_);
  or _86734_ (_36916_, _11515_, _05894_);
  and _86735_ (_36917_, _36916_, _05886_);
  nand _86736_ (_36918_, _36917_, _36915_);
  nor _86737_ (_36919_, _11378_, _05886_);
  nor _86738_ (_36920_, _36919_, _08363_);
  nand _86739_ (_36921_, _36920_, _36918_);
  and _86740_ (_36922_, _11514_, _08363_);
  nor _86741_ (_36923_, _36922_, _11347_);
  nand _86742_ (_36925_, _36923_, _36921_);
  nor _86743_ (_36926_, _11809_, \oc8051_golden_model_1.DPH [6]);
  nor _86744_ (_36927_, _36926_, _11810_);
  nor _86745_ (_36928_, _36927_, _11348_);
  nor _86746_ (_36929_, _36928_, _11816_);
  and _86747_ (_36930_, _36929_, _36925_);
  or _86748_ (_36931_, _36930_, _36783_);
  nand _86749_ (_36932_, _36931_, _11820_);
  and _86750_ (_36933_, _11514_, _08786_);
  and _86751_ (_36934_, _36798_, _11826_);
  or _86752_ (_36936_, _36934_, _36933_);
  and _86753_ (_36937_, _36936_, _11819_);
  nor _86754_ (_36938_, _36937_, _11824_);
  nand _86755_ (_36939_, _36938_, _36932_);
  nor _86756_ (_36940_, _36777_, _11345_);
  nor _86757_ (_36941_, _36940_, _11342_);
  nand _86758_ (_36942_, _36941_, _36939_);
  nor _86759_ (_36943_, _11515_, _11341_);
  nor _86760_ (_36944_, _36943_, _03600_);
  nand _86761_ (_36945_, _36944_, _36942_);
  nor _86762_ (_36947_, _11378_, _07766_);
  nor _86763_ (_36948_, _36947_, _36024_);
  and _86764_ (_36949_, _36948_, _36945_);
  or _86765_ (_36950_, _36949_, _36782_);
  nand _86766_ (_36951_, _36950_, _11842_);
  or _86767_ (_36952_, _36798_, _11826_);
  or _86768_ (_36953_, _11514_, _08786_);
  and _86769_ (_36954_, _36953_, _11841_);
  and _86770_ (_36955_, _36954_, _36952_);
  nor _86771_ (_36956_, _36955_, _11853_);
  nand _86772_ (_36958_, _36956_, _36951_);
  nor _86773_ (_36959_, _36777_, _11851_);
  nor _86774_ (_36960_, _36959_, _08431_);
  nand _86775_ (_36961_, _36960_, _36958_);
  nor _86776_ (_36962_, _11515_, _08430_);
  nor _86777_ (_36963_, _36962_, _03622_);
  nand _86778_ (_36964_, _36963_, _36961_);
  nor _86779_ (_36965_, _11378_, _07777_);
  nor _86780_ (_36966_, _36965_, _10754_);
  and _86781_ (_36967_, _36966_, _36964_);
  or _86782_ (_36969_, _36967_, _36780_);
  nand _86783_ (_36970_, _36969_, _11338_);
  and _86784_ (_36971_, _11514_, \oc8051_golden_model_1.PSW [7]);
  and _86785_ (_36972_, _36798_, _07871_);
  or _86786_ (_36973_, _36972_, _36971_);
  and _86787_ (_36974_, _36973_, _11337_);
  nor _86788_ (_36975_, _36974_, _11864_);
  nand _86789_ (_36976_, _36975_, _36970_);
  nor _86790_ (_36977_, _36777_, _11335_);
  nor _86791_ (_36978_, _36977_, _08460_);
  nand _86792_ (_36980_, _36978_, _36976_);
  nor _86793_ (_36981_, _11515_, _08459_);
  nor _86794_ (_36982_, _36981_, _03624_);
  nand _86795_ (_36983_, _36982_, _36980_);
  nor _86796_ (_36984_, _11378_, _07795_);
  nor _86797_ (_36985_, _36984_, _36063_);
  and _86798_ (_36986_, _36985_, _36983_);
  or _86799_ (_36987_, _36986_, _36779_);
  nand _86800_ (_36988_, _36987_, _11881_);
  nor _86801_ (_36989_, _36798_, _07871_);
  nor _86802_ (_36991_, _11514_, \oc8051_golden_model_1.PSW [7]);
  nor _86803_ (_36992_, _36991_, _11881_);
  not _86804_ (_36993_, _36992_);
  nor _86805_ (_36994_, _36993_, _36989_);
  nor _86806_ (_36995_, _36994_, _11885_);
  nand _86807_ (_36996_, _36995_, _36988_);
  nor _86808_ (_36997_, _36777_, _11330_);
  nor _86809_ (_36998_, _36997_, _08508_);
  nand _86810_ (_36999_, _36998_, _36996_);
  nor _86811_ (_37000_, _11515_, _08507_);
  nor _86812_ (_37002_, _37000_, _08587_);
  nand _86813_ (_37003_, _37002_, _36999_);
  nor _86814_ (_37004_, _36777_, _08588_);
  nor _86815_ (_37005_, _37004_, _03798_);
  and _86816_ (_37006_, _37005_, _37003_);
  nor _86817_ (_37007_, _05363_, _10652_);
  or _86818_ (_37008_, _37007_, _03188_);
  or _86819_ (_37009_, _37008_, _37006_);
  nor _86820_ (_37010_, _11514_, _06399_);
  nor _86821_ (_37011_, _37010_, _03621_);
  nand _86822_ (_37013_, _37011_, _37009_);
  nor _86823_ (_37014_, _11378_, _09854_);
  and _86824_ (_37015_, _36848_, _09854_);
  or _86825_ (_37016_, _37015_, _11903_);
  or _86826_ (_37017_, _37016_, _37014_);
  and _86827_ (_37018_, _37017_, _11328_);
  nand _86828_ (_37019_, _37018_, _37013_);
  nor _86829_ (_37020_, _36777_, _11328_);
  nor _86830_ (_37021_, _37020_, _08703_);
  nand _86831_ (_37022_, _37021_, _37019_);
  nor _86832_ (_37024_, _11515_, _08702_);
  nor _86833_ (_37025_, _37024_, _08732_);
  and _86834_ (_37026_, _37025_, _37022_);
  or _86835_ (_37027_, _37026_, _36778_);
  nand _86836_ (_37028_, _37027_, _03516_);
  and _86837_ (_37029_, _05363_, _03515_);
  nor _86838_ (_37030_, _37029_, _03203_);
  and _86839_ (_37031_, _37030_, _37028_);
  and _86840_ (_37032_, _11514_, _03203_);
  or _86841_ (_37033_, _37032_, _03628_);
  nor _86842_ (_37035_, _37033_, _37031_);
  and _86843_ (_37036_, _11379_, _09854_);
  nor _86844_ (_37037_, _36785_, _09854_);
  nor _86845_ (_37038_, _37037_, _37036_);
  nor _86846_ (_37039_, _37038_, _03816_);
  or _86847_ (_37040_, _37039_, _37035_);
  and _86848_ (_37041_, _37040_, _11933_);
  nor _86849_ (_37042_, _36777_, _11933_);
  or _86850_ (_37043_, _37042_, _37041_);
  nand _86851_ (_37044_, _37043_, _04246_);
  nor _86852_ (_37046_, _11514_, _04246_);
  nor _86853_ (_37047_, _37046_, _32765_);
  nand _86854_ (_37048_, _37047_, _37044_);
  nor _86855_ (_37049_, _36816_, _11940_);
  nor _86856_ (_37050_, _37049_, _03629_);
  nand _86857_ (_37051_, _37050_, _37048_);
  and _86858_ (_37052_, _03629_, _03549_);
  nor _86859_ (_37053_, _37052_, _03198_);
  nand _86860_ (_37054_, _37053_, _37051_);
  and _86861_ (_37055_, _11514_, _03198_);
  nor _86862_ (_37057_, _37055_, _03453_);
  nand _86863_ (_37058_, _37057_, _37054_);
  nor _86864_ (_37059_, _37038_, _03823_);
  nor _86865_ (_37060_, _37059_, _11958_);
  nand _86866_ (_37061_, _37060_, _37058_);
  nor _86867_ (_37062_, _36816_, _11957_);
  nor _86868_ (_37063_, _37062_, _03447_);
  nand _86869_ (_37064_, _37063_, _37061_);
  nor _86870_ (_37065_, _11514_, _03514_);
  nor _86871_ (_37066_, _37065_, _33825_);
  nand _86872_ (_37068_, _37066_, _37064_);
  nor _86873_ (_37069_, _36816_, _11964_);
  nor _86874_ (_37070_, _37069_, _03631_);
  nand _86875_ (_37071_, _37070_, _37068_);
  and _86876_ (_37072_, _03631_, _03549_);
  nor _86877_ (_37073_, _37072_, _03196_);
  nand _86878_ (_37074_, _37073_, _37071_);
  and _86879_ (_37075_, _11514_, _03196_);
  nor _86880_ (_37076_, _37075_, _11975_);
  and _86881_ (_37077_, _37076_, _37074_);
  nor _86882_ (_37079_, _36777_, _11976_);
  nor _86883_ (_37080_, _37079_, _37077_);
  or _86884_ (_37081_, _37080_, _43004_);
  or _86885_ (_37082_, _43000_, \oc8051_golden_model_1.PC [14]);
  and _86886_ (_37083_, _37082_, _41806_);
  and _86887_ (_43685_, _37083_, _37081_);
  and _86888_ (_37084_, _43004_, \oc8051_golden_model_1.P0INREG [0]);
  or _86889_ (_37085_, _37084_, _01169_);
  and _86890_ (_43686_, _37085_, _41806_);
  and _86891_ (_37086_, _43004_, \oc8051_golden_model_1.P0INREG [1]);
  or _86892_ (_37088_, _37086_, _01153_);
  and _86893_ (_43687_, _37088_, _41806_);
  and _86894_ (_37089_, _43004_, \oc8051_golden_model_1.P0INREG [2]);
  or _86895_ (_37090_, _37089_, _01186_);
  and _86896_ (_43688_, _37090_, _41806_);
  and _86897_ (_37091_, _43004_, \oc8051_golden_model_1.P0INREG [3]);
  or _86898_ (_37092_, _37091_, _01202_);
  and _86899_ (_43689_, _37092_, _41806_);
  and _86900_ (_37093_, _43004_, \oc8051_golden_model_1.P0INREG [4]);
  or _86901_ (_37094_, _37093_, _01162_);
  and _86902_ (_43690_, _37094_, _41806_);
  and _86903_ (_37096_, _43004_, \oc8051_golden_model_1.P0INREG [5]);
  or _86904_ (_37097_, _37096_, _01146_);
  and _86905_ (_43691_, _37097_, _41806_);
  and _86906_ (_37098_, _43004_, \oc8051_golden_model_1.P0INREG [6]);
  or _86907_ (_37099_, _37098_, _01179_);
  and _86908_ (_43692_, _37099_, _41806_);
  and _86909_ (_37100_, _43004_, \oc8051_golden_model_1.P1INREG [0]);
  or _86910_ (_37101_, _37100_, _01133_);
  and _86911_ (_43695_, _37101_, _41806_);
  and _86912_ (_37103_, _43004_, \oc8051_golden_model_1.P1INREG [1]);
  or _86913_ (_37104_, _37103_, _01083_);
  and _86914_ (_43696_, _37104_, _41806_);
  and _86915_ (_37105_, _43004_, \oc8051_golden_model_1.P1INREG [2]);
  or _86916_ (_37106_, _37105_, _01117_);
  and _86917_ (_43697_, _37106_, _41806_);
  and _86918_ (_37107_, _43004_, \oc8051_golden_model_1.P1INREG [3]);
  or _86919_ (_37108_, _37107_, _01099_);
  and _86920_ (_43698_, _37108_, _41806_);
  and _86921_ (_37109_, _43004_, \oc8051_golden_model_1.P1INREG [4]);
  or _86922_ (_37111_, _37109_, _01126_);
  and _86923_ (_43699_, _37111_, _41806_);
  and _86924_ (_37112_, _43004_, \oc8051_golden_model_1.P1INREG [5]);
  or _86925_ (_37113_, _37112_, _01076_);
  and _86926_ (_43702_, _37113_, _41806_);
  and _86927_ (_37114_, _43004_, \oc8051_golden_model_1.P1INREG [6]);
  or _86928_ (_37115_, _37114_, _01110_);
  and _86929_ (_43703_, _37115_, _41806_);
  and _86930_ (_37116_, _43004_, \oc8051_golden_model_1.P2INREG [0]);
  or _86931_ (_37117_, _37116_, _00899_);
  and _86932_ (_43704_, _37117_, _41806_);
  and _86933_ (_37119_, _43004_, \oc8051_golden_model_1.P2INREG [1]);
  or _86934_ (_37120_, _37119_, _00926_);
  and _86935_ (_43705_, _37120_, _41806_);
  and _86936_ (_37121_, _43004_, \oc8051_golden_model_1.P2INREG [2]);
  or _86937_ (_37122_, _37121_, _00874_);
  and _86938_ (_43706_, _37122_, _41806_);
  and _86939_ (_37123_, _43004_, \oc8051_golden_model_1.P2INREG [3]);
  or _86940_ (_37124_, _37123_, _00916_);
  and _86941_ (_43707_, _37124_, _41806_);
  and _86942_ (_37126_, _43004_, \oc8051_golden_model_1.P2INREG [4]);
  or _86943_ (_37127_, _37126_, _00891_);
  and _86944_ (_43708_, _37127_, _41806_);
  and _86945_ (_37128_, _43004_, \oc8051_golden_model_1.P2INREG [5]);
  or _86946_ (_37129_, _37128_, _00933_);
  and _86947_ (_43709_, _37129_, _41806_);
  and _86948_ (_37130_, _43004_, \oc8051_golden_model_1.P2INREG [6]);
  or _86949_ (_37131_, _37130_, _00881_);
  and _86950_ (_43710_, _37131_, _41806_);
  and _86951_ (_37132_, _43004_, \oc8051_golden_model_1.P3INREG [0]);
  or _86952_ (_37134_, _37132_, _01019_);
  and _86953_ (_43713_, _37134_, _41806_);
  and _86954_ (_37135_, _43004_, \oc8051_golden_model_1.P3INREG [1]);
  or _86955_ (_37136_, _37135_, _01045_);
  and _86956_ (_43714_, _37136_, _41806_);
  and _86957_ (_37137_, _43004_, \oc8051_golden_model_1.P3INREG [2]);
  or _86958_ (_37138_, _37137_, _00996_);
  and _86959_ (_43715_, _37138_, _41806_);
  and _86960_ (_37139_, _43004_, \oc8051_golden_model_1.P3INREG [3]);
  or _86961_ (_37140_, _37139_, _01035_);
  and _86962_ (_43716_, _37140_, _41806_);
  and _86963_ (_37142_, _43004_, \oc8051_golden_model_1.P3INREG [4]);
  or _86964_ (_37143_, _37142_, _01012_);
  and _86965_ (_43717_, _37143_, _41806_);
  and _86966_ (_37144_, _43004_, \oc8051_golden_model_1.P3INREG [5]);
  or _86967_ (_37145_, _37144_, _01052_);
  and _86968_ (_43718_, _37145_, _41806_);
  and _86969_ (_37146_, _43004_, \oc8051_golden_model_1.P3INREG [6]);
  or _86970_ (_37147_, _37146_, _01003_);
  and _86971_ (_43719_, _37147_, _41806_);
  nor _86972_ (_00005_[6], _01004_, rst);
  nor _86973_ (_00005_[5], _01053_, rst);
  nor _86974_ (_00005_[4], _01013_, rst);
  nor _86975_ (_00005_[3], _01036_, rst);
  nor _86976_ (_00005_[2], _00997_, rst);
  nor _86977_ (_00005_[1], _01046_, rst);
  nor _86978_ (_00005_[0], _01020_, rst);
  nor _86979_ (_00004_[6], _00882_, rst);
  nor _86980_ (_00004_[5], _00934_, rst);
  nor _86981_ (_00004_[4], _00892_, rst);
  nor _86982_ (_00004_[3], _00917_, rst);
  nor _86983_ (_00004_[2], _00875_, rst);
  nor _86984_ (_00004_[1], _00927_, rst);
  nor _86985_ (_00004_[0], _00900_, rst);
  nor _86986_ (_00003_[6], _01111_, rst);
  nor _86987_ (_00003_[5], _01077_, rst);
  nor _86988_ (_00003_[4], _01127_, rst);
  nor _86989_ (_00003_[3], _01100_, rst);
  nor _86990_ (_00003_[2], _01118_, rst);
  nor _86991_ (_00003_[1], _01084_, rst);
  nor _86992_ (_00003_[0], _01134_, rst);
  nor _86993_ (_00002_[6], _01180_, rst);
  nor _86994_ (_00002_[5], _01147_, rst);
  nor _86995_ (_00002_[4], _01163_, rst);
  nor _86996_ (_00002_[3], _01203_, rst);
  nor _86997_ (_00002_[2], _01187_, rst);
  nor _86998_ (_00002_[1], _01154_, rst);
  nor _86999_ (_00002_[0], _01170_, rst);
  or _87000_ (_37151_, _10641_, _09230_);
  nor _87001_ (_37152_, _37151_, _10903_);
  not _87002_ (_37154_, _28767_);
  and _87003_ (_37155_, _37154_, _28534_);
  nor _87004_ (_37156_, _29111_, _28997_);
  and _87005_ (_37157_, _37156_, _37155_);
  nor _87006_ (_37158_, _27118_, _27001_);
  nor _87007_ (_37159_, _27463_, _27349_);
  and _87008_ (_37160_, _37159_, _37158_);
  nor _87009_ (_37161_, _19863_, _19634_);
  nor _87010_ (_37162_, _26885_, _19976_);
  and _87011_ (_37163_, _37162_, _37161_);
  and _87012_ (_37165_, _37163_, _37160_);
  and _87013_ (_37166_, _37165_, _37157_);
  nor _87014_ (_37167_, _11230_, _11148_);
  nor _87015_ (_37168_, _18722_, _11311_);
  and _87016_ (_37169_, _37168_, _37167_);
  nor _87017_ (_37170_, _10533_, _10452_);
  nor _87018_ (_37171_, _11066_, _10985_);
  and _87019_ (_37172_, _37171_, _37170_);
  and _87020_ (_37173_, _37172_, _37169_);
  not _87021_ (_37174_, _26774_);
  nor _87022_ (_37176_, _37174_, _19517_);
  not _87023_ (_37177_, _28423_);
  nor _87024_ (_37178_, _28650_, _37177_);
  nand _87025_ (_37179_, _37178_, _37176_);
  nor _87026_ (_37180_, _37179_, _18954_);
  and _87027_ (_37181_, _37180_, _37173_);
  nor _87028_ (_37182_, _19068_, _18839_);
  nor _87029_ (_37183_, _19400_, _19182_);
  and _87030_ (_37184_, _37183_, _37182_);
  or _87031_ (_37185_, _31193_, _29972_);
  nor _87032_ (_37187_, _37185_, _31800_);
  or _87033_ (_37188_, _11764_, _03165_);
  nor _87034_ (_37189_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor _87035_ (_37190_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor _87036_ (_37191_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and _87037_ (_37192_, _37191_, _37190_);
  and _87038_ (_37193_, _37192_, _37189_);
  nor _87039_ (_37194_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor _87040_ (_37195_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and _87041_ (_37196_, _37195_, _37194_);
  nor _87042_ (_37198_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor _87043_ (_37199_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and _87044_ (_37200_, _37199_, _37198_);
  and _87045_ (_37201_, _37200_, _37196_);
  and _87046_ (_37202_, _37201_, _37193_);
  nor _87047_ (_37203_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor _87048_ (_37204_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and _87049_ (_37205_, _37204_, _37203_);
  nor _87050_ (_37206_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor _87051_ (_37207_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and _87052_ (_37209_, _37207_, _37206_);
  and _87053_ (_37210_, _37209_, _37205_);
  nor _87054_ (_37211_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor _87055_ (_37212_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and _87056_ (_37213_, _37212_, _37211_);
  nor _87057_ (_37214_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor _87058_ (_37215_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and _87059_ (_37216_, _37215_, _37214_);
  and _87060_ (_37217_, _37216_, _37213_);
  and _87061_ (_37218_, _37217_, _37210_);
  and _87062_ (_37220_, _37218_, _37202_);
  nor _87063_ (_37221_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor _87064_ (_37222_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and _87065_ (_37223_, _37222_, _37221_);
  nor _87066_ (_37224_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor _87067_ (_37225_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and _87068_ (_37226_, _37225_, _37224_);
  and _87069_ (_37227_, _37226_, _37223_);
  nor _87070_ (_37228_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  nor _87071_ (_37229_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  and _87072_ (_37231_, _37229_, _37228_);
  nor _87073_ (_37232_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor _87074_ (_37233_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and _87075_ (_37234_, _37233_, _37232_);
  and _87076_ (_37235_, _37234_, _37231_);
  and _87077_ (_37236_, _37235_, _37227_);
  nor _87078_ (_37237_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor _87079_ (_37238_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and _87080_ (_37239_, _37238_, _37237_);
  nor _87081_ (_37240_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  nor _87082_ (_37242_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  and _87083_ (_37243_, _37242_, _37240_);
  and _87084_ (_37244_, _37243_, _37239_);
  nor _87085_ (_37245_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor _87086_ (_37246_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and _87087_ (_37247_, _37246_, _37245_);
  nor _87088_ (_37248_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor _87089_ (_37249_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and _87090_ (_37250_, _37249_, _37248_);
  and _87091_ (_37251_, _37250_, _37247_);
  and _87092_ (_37253_, _37251_, _37244_);
  and _87093_ (_37254_, _37253_, _37236_);
  nor _87094_ (_37255_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and _87095_ (_37256_, _37255_, op0_cnst);
  nor _87096_ (_37257_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor _87097_ (_37258_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and _87098_ (_37259_, _37258_, _37257_);
  nor _87099_ (_37260_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor _87100_ (_37261_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and _87101_ (_37262_, _37261_, _37260_);
  and _87102_ (_37264_, _37262_, _37259_);
  and _87103_ (_37265_, _37264_, _37256_);
  nor _87104_ (_37266_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor _87105_ (_37267_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and _87106_ (_37268_, _37267_, _37266_);
  nor _87107_ (_37269_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor _87108_ (_37270_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and _87109_ (_37271_, _37270_, _37269_);
  and _87110_ (_37272_, _37271_, _37268_);
  and _87111_ (_37273_, \oc8051_golden_model_1.TCON [1], _28320_);
  nor _87112_ (_37275_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and _87113_ (_37276_, _37275_, _37273_);
  nor _87114_ (_37277_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor _87115_ (_37278_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and _87116_ (_37279_, _37278_, _37277_);
  and _87117_ (_37280_, _37279_, _37276_);
  and _87118_ (_37281_, _37280_, _37272_);
  and _87119_ (_37282_, _37281_, _37265_);
  and _87120_ (_37283_, _37282_, _37254_);
  and _87121_ (_37284_, _37283_, _37220_);
  nand _87122_ (_37286_, _37284_, _37188_);
  nor _87123_ (_37287_, _37286_, _25536_);
  nor _87124_ (_37288_, _29192_, _26140_);
  and _87125_ (_37289_, _37288_, _37287_);
  nor _87126_ (_37290_, _26316_, _25712_);
  and _87127_ (_37291_, _37290_, _37289_);
  and _87128_ (_37292_, _37291_, _37187_);
  nor _87129_ (_37293_, _26227_, _25623_);
  and _87130_ (_37294_, _37293_, _37292_);
  nor _87131_ (_37295_, _29884_, _29454_);
  nor _87132_ (_37297_, _30586_, _30058_);
  and _87133_ (_37298_, _37297_, _37295_);
  nor _87134_ (_37299_, _30398_, _29799_);
  nor _87135_ (_37300_, _31624_, _31016_);
  nand _87136_ (_37301_, _37300_, _37299_);
  nor _87137_ (_37302_, _37301_, _25798_);
  nor _87138_ (_37303_, _29368_, _26403_);
  and _87139_ (_37304_, _37303_, _37302_);
  and _87140_ (_37305_, _37304_, _37298_);
  and _87141_ (_37306_, _37305_, _37294_);
  nor _87142_ (_37308_, _30497_, _29279_);
  nor _87143_ (_37309_, _31711_, _31104_);
  nand _87144_ (_37310_, _37309_, _37308_);
  nor _87145_ (_37311_, _37310_, _19289_);
  and _87146_ (_37312_, _37311_, _37306_);
  nor _87147_ (_37313_, _29629_, _26666_);
  nor _87148_ (_37314_, _30233_, _29716_);
  and _87149_ (_37315_, _37314_, _37313_);
  or _87150_ (_37316_, _31280_, _30672_);
  or _87151_ (_37317_, _37316_, _31886_);
  nor _87152_ (_37319_, _37317_, _25973_);
  nor _87153_ (_37320_, _26579_, _26059_);
  and _87154_ (_37321_, _37320_, _37319_);
  and _87155_ (_37322_, _37321_, _37315_);
  and _87156_ (_37323_, _37322_, _37312_);
  or _87157_ (_37324_, _31369_, _30760_);
  nor _87158_ (_37325_, _37324_, _31975_);
  nor _87159_ (_37326_, _26492_, _25886_);
  nor _87160_ (_37327_, _30146_, _29543_);
  and _87161_ (_37328_, _37327_, _37326_);
  and _87162_ (_37330_, _37328_, _37325_);
  and _87163_ (_37331_, _37330_, _37323_);
  or _87164_ (_37332_, _32061_, _31542_);
  nor _87165_ (_37333_, _37332_, _32147_);
  nor _87166_ (_37334_, _30846_, _30319_);
  nor _87167_ (_37335_, _31456_, _30933_);
  and _87168_ (_37336_, _37335_, _37334_);
  nand _87169_ (_37337_, _37336_, _37333_);
  or _87170_ (_37338_, _37337_, _18494_);
  nor _87171_ (_37339_, _37338_, _18606_);
  and _87172_ (_37341_, _37339_, _37331_);
  and _87173_ (_37342_, _37341_, _37184_);
  and _87174_ (_37343_, _37342_, _37181_);
  or _87175_ (_37344_, _27234_, _19749_);
  or _87176_ (_37345_, _37344_, _28882_);
  nor _87177_ (_37346_, _37345_, _09123_);
  and _87178_ (_37347_, _37346_, _37343_);
  and _87179_ (_37348_, _37347_, _37166_);
  and _87180_ (_37349_, _37348_, _37152_);
  and _87181_ (_37350_, _37349_, _43000_);
  and _87182_ (_37352_, _37350_, _41806_);
  nor _87183_ (_37353_, _10796_, _38443_);
  and _87184_ (_37354_, _10796_, _38443_);
  or _87185_ (_37355_, _37354_, _37353_);
  and _87186_ (_37356_, _28315_, _38487_);
  nor _87187_ (_37357_, _28315_, _38487_);
  or _87188_ (_37358_, _37357_, _37356_);
  and _87189_ (_37359_, _28181_, _38481_);
  or _87190_ (_37360_, _27548_, _40411_);
  nand _87191_ (_37361_, _27548_, _40411_);
  and _87192_ (_37363_, _37361_, _37360_);
  or _87193_ (_37364_, _27668_, _38457_);
  nand _87194_ (_37365_, _27668_, _38457_);
  and _87195_ (_37366_, _37365_, _37364_);
  or _87196_ (_37367_, _37366_, _37363_);
  and _87197_ (_37368_, _27790_, _38463_);
  nor _87198_ (_37369_, _27790_, _38463_);
  or _87199_ (_37370_, _37369_, _37368_);
  or _87200_ (_37371_, _37370_, _37367_);
  or _87201_ (_37372_, _37371_, _37359_);
  nor _87202_ (_37374_, _27912_, _38469_);
  and _87203_ (_37375_, _27912_, _38469_);
  or _87204_ (_37376_, _37375_, _37374_);
  or _87205_ (_37377_, _28046_, _40511_);
  nand _87206_ (_37378_, _28046_, _40511_);
  and _87207_ (_37379_, _37378_, _37377_);
  nor _87208_ (_37380_, _28181_, _38481_);
  or _87209_ (_37381_, _37380_, _37379_);
  or _87210_ (_37382_, _37381_, _37376_);
  or _87211_ (_37383_, _37382_, _37372_);
  or _87212_ (_37385_, _37383_, _37358_);
  or _87213_ (_37386_, _37385_, _37355_);
  and _87214_ (_00007_, _37386_, _37352_);
  nor _87215_ (_37387_, _25047_, _40277_);
  and _87216_ (_37388_, _25047_, _40277_);
  or _87217_ (_37389_, _37388_, _37387_);
  and _87218_ (_37390_, _25164_, _38949_);
  nor _87219_ (_37391_, _25164_, _38949_);
  or _87220_ (_37392_, _37391_, _37390_);
  or _87221_ (_37393_, _37392_, _37389_);
  nor _87222_ (_37395_, _24693_, _38864_);
  and _87223_ (_37396_, _24693_, _38864_);
  or _87224_ (_37397_, _37396_, _37395_);
  not _87225_ (_37398_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor _87226_ (_37399_, _25279_, _37398_);
  and _87227_ (_37400_, _25279_, _37398_);
  or _87228_ (_37401_, _37400_, _37399_);
  or _87229_ (_37402_, _37401_, _37397_);
  or _87230_ (_37403_, _37402_, _37393_);
  and _87231_ (_37404_, _25455_, _31066_);
  nor _87232_ (_37406_, _25455_, _31066_);
  or _87233_ (_37407_, _37406_, _37404_);
  or _87234_ (_37408_, _37407_, _37403_);
  and _87235_ (_37409_, _24932_, _38901_);
  nor _87236_ (_37410_, _24932_, _38901_);
  or _87237_ (_37411_, _37410_, _37409_);
  or _87238_ (_37412_, _37411_, _37408_);
  and _87239_ (_37413_, _10371_, _38839_);
  nor _87240_ (_37414_, _10371_, _38839_);
  or _87241_ (_37415_, _37414_, _37413_);
  or _87242_ (_37417_, _37415_, _37412_);
  and _87243_ (_00006_, _37417_, _37352_);
  or _87244_ (_00001_, _37349_, rst);
  nor _87245_ (_00005_[7], _01029_, rst);
  nor _87246_ (_00004_[7], _00909_, rst);
  nor _87247_ (_00003_[7], _01093_, rst);
  nor _87248_ (_00002_[7], _01196_, rst);
  and _87249_ (_37418_, _37349_, inst_finished_r);
  nor _87250_ (_37419_, _38443_, \oc8051_golden_model_1.SP [7]);
  and _87251_ (_37420_, _38443_, \oc8051_golden_model_1.SP [7]);
  or _87252_ (_37422_, _37420_, _37419_);
  nor _87253_ (_37423_, _38487_, \oc8051_golden_model_1.SP [6]);
  and _87254_ (_37424_, _38487_, \oc8051_golden_model_1.SP [6]);
  or _87255_ (_37425_, _37424_, _37423_);
  nor _87256_ (_37426_, _38481_, \oc8051_golden_model_1.SP [5]);
  and _87257_ (_37427_, _38481_, \oc8051_golden_model_1.SP [5]);
  or _87258_ (_37428_, _37427_, _37426_);
  nor _87259_ (_37429_, _38469_, \oc8051_golden_model_1.SP [3]);
  and _87260_ (_37430_, _38469_, \oc8051_golden_model_1.SP [3]);
  or _87261_ (_37431_, _37430_, _37429_);
  and _87262_ (_37433_, _38457_, \oc8051_golden_model_1.SP [1]);
  nor _87263_ (_37434_, _38451_, \oc8051_golden_model_1.SP [0]);
  and _87264_ (_37435_, _38451_, \oc8051_golden_model_1.SP [0]);
  or _87265_ (_37436_, _37435_, _37434_);
  nor _87266_ (_37437_, _38457_, \oc8051_golden_model_1.SP [1]);
  or _87267_ (_37438_, _37437_, _37436_);
  or _87268_ (_37439_, _37438_, _37433_);
  nor _87269_ (_37440_, _38463_, \oc8051_golden_model_1.SP [2]);
  and _87270_ (_37441_, _38463_, \oc8051_golden_model_1.SP [2]);
  or _87271_ (_37442_, _37441_, _37440_);
  or _87272_ (_37444_, _37442_, _37439_);
  or _87273_ (_37445_, _37444_, _37431_);
  nor _87274_ (_37446_, _38475_, \oc8051_golden_model_1.SP [4]);
  and _87275_ (_37447_, _38475_, \oc8051_golden_model_1.SP [4]);
  or _87276_ (_37448_, _37447_, _37446_);
  or _87277_ (_37449_, _37448_, _37445_);
  or _87278_ (_37450_, _37449_, _37428_);
  or _87279_ (_37451_, _37450_, _37425_);
  or _87280_ (_37452_, _37451_, _37422_);
  and _87281_ (_37453_, _37452_, property_invalid_sp_1_r);
  and _87282_ (property_invalid_sp, _37453_, _37418_);
  and _87283_ (_37455_, _25052_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _87284_ (_37456_, \oc8051_golden_model_1.PSW [4], _38949_);
  or _87285_ (_37457_, _37456_, _37455_);
  and _87286_ (_37458_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _87287_ (_37459_, \oc8051_golden_model_1.PSW [3], _40277_);
  or _87288_ (_37460_, _37459_, _37458_);
  or _87289_ (_37461_, _37460_, _37457_);
  and _87290_ (_37462_, _24593_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _87291_ (_37463_, \oc8051_golden_model_1.PSW [1], _38864_);
  or _87292_ (_37465_, _37463_, _37462_);
  nand _87293_ (_37466_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _87294_ (_37467_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _87295_ (_37468_, _37467_, _37466_);
  or _87296_ (_37469_, _37468_, _37465_);
  or _87297_ (_37470_, _37469_, _37461_);
  and _87298_ (_37471_, _07871_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _87299_ (_37472_, \oc8051_golden_model_1.PSW [7], _38839_);
  or _87300_ (_37473_, _37472_, _37471_);
  and _87301_ (_37474_, _25169_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _87302_ (_37476_, \oc8051_golden_model_1.PSW [5], _37398_);
  or _87303_ (_37477_, _37476_, _37474_);
  nand _87304_ (_37478_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _87305_ (_37479_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _87306_ (_37480_, _37479_, _37478_);
  or _87307_ (_37481_, _37480_, _37477_);
  or _87308_ (_37482_, _37481_, _37473_);
  or _87309_ (_37483_, _37482_, _37470_);
  and _87310_ (_37484_, _37483_, property_invalid_psw_1_r);
  and _87311_ (property_invalid_psw, _37484_, _37418_);
  nand _87312_ (_37486_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _87313_ (_37487_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _87314_ (_37488_, _37487_, _37486_);
  and _87315_ (_37489_, _22590_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _87316_ (_37490_, \oc8051_golden_model_1.P3 [2], _39721_);
  or _87317_ (_37491_, _37490_, _37489_);
  or _87318_ (_37492_, _37491_, _37488_);
  and _87319_ (_37493_, \oc8051_golden_model_1.P3 [0], _39688_);
  and _87320_ (_37494_, _22373_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _87321_ (_37495_, _37494_, _37493_);
  and _87322_ (_37497_, _22487_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _87323_ (_37498_, \oc8051_golden_model_1.P3 [1], _39701_);
  or _87324_ (_37499_, _37498_, _37497_);
  or _87325_ (_37500_, _37499_, _37495_);
  or _87326_ (_37501_, _37500_, _37492_);
  or _87327_ (_37502_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand _87328_ (_37503_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _87329_ (_37504_, _37503_, _37502_);
  or _87330_ (_37505_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand _87331_ (_37506_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _87332_ (_37508_, _37506_, _37505_);
  or _87333_ (_37509_, _37508_, _37504_);
  and _87334_ (_37510_, _09553_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _87335_ (_37511_, \oc8051_golden_model_1.P3 [7], _39241_);
  or _87336_ (_37512_, _37511_, _37510_);
  nand _87337_ (_37513_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _87338_ (_37514_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _87339_ (_37515_, _37514_, _37513_);
  or _87340_ (_37516_, _37515_, _37512_);
  or _87341_ (_37517_, _37516_, _37509_);
  or _87342_ (_37519_, _37517_, _37501_);
  and _87343_ (property_invalid_p3, _37519_, _37418_);
  nand _87344_ (_37520_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _87345_ (_37521_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _87346_ (_37522_, _37521_, _37520_);
  and _87347_ (_37523_, _21818_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _87348_ (_37524_, \oc8051_golden_model_1.P2 [2], _39619_);
  or _87349_ (_37525_, _37524_, _37523_);
  or _87350_ (_37526_, _37525_, _37522_);
  and _87351_ (_37527_, \oc8051_golden_model_1.P2 [0], _39592_);
  and _87352_ (_37529_, _21602_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _87353_ (_37530_, _37529_, _37527_);
  and _87354_ (_37531_, _21716_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _87355_ (_37532_, \oc8051_golden_model_1.P2 [1], _39605_);
  or _87356_ (_37533_, _37532_, _37531_);
  or _87357_ (_37534_, _37533_, _37530_);
  or _87358_ (_37535_, _37534_, _37526_);
  or _87359_ (_37536_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand _87360_ (_37537_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _87361_ (_37538_, _37537_, _37536_);
  or _87362_ (_37540_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand _87363_ (_37541_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _87364_ (_37542_, _37541_, _37540_);
  or _87365_ (_37543_, _37542_, _37538_);
  and _87366_ (_37544_, _09450_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _87367_ (_37545_, \oc8051_golden_model_1.P2 [7], _39183_);
  or _87368_ (_37546_, _37545_, _37544_);
  nand _87369_ (_37547_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _87370_ (_37548_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _87371_ (_37549_, _37548_, _37547_);
  or _87372_ (_37551_, _37549_, _37546_);
  or _87373_ (_37552_, _37551_, _37543_);
  or _87374_ (_37553_, _37552_, _37535_);
  and _87375_ (property_invalid_p2, _37553_, _37418_);
  nand _87376_ (_37554_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _87377_ (_37555_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _87378_ (_37556_, _37555_, _37554_);
  and _87379_ (_37557_, _21045_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _87380_ (_37558_, \oc8051_golden_model_1.P1 [2], _39528_);
  or _87381_ (_37559_, _37558_, _37557_);
  or _87382_ (_37561_, _37559_, _37556_);
  and _87383_ (_37562_, \oc8051_golden_model_1.P1 [0], _39502_);
  and _87384_ (_37563_, _20834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _87385_ (_37564_, _37563_, _37562_);
  and _87386_ (_37565_, _20944_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _87387_ (_37566_, \oc8051_golden_model_1.P1 [1], _39515_);
  or _87388_ (_37567_, _37566_, _37565_);
  or _87389_ (_37568_, _37567_, _37564_);
  or _87390_ (_37569_, _37568_, _37561_);
  or _87391_ (_37570_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand _87392_ (_37572_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _87393_ (_37573_, _37572_, _37570_);
  or _87394_ (_37574_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand _87395_ (_37575_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _87396_ (_37576_, _37575_, _37574_);
  or _87397_ (_37577_, _37576_, _37573_);
  and _87398_ (_37578_, _09348_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _87399_ (_37579_, \oc8051_golden_model_1.P1 [7], _39165_);
  or _87400_ (_37580_, _37579_, _37578_);
  nand _87401_ (_37581_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _87402_ (_37583_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _87403_ (_37584_, _37583_, _37581_);
  or _87404_ (_37585_, _37584_, _37580_);
  or _87405_ (_37586_, _37585_, _37577_);
  or _87406_ (_37587_, _37586_, _37569_);
  and _87407_ (property_invalid_p1, _37587_, _37418_);
  nand _87408_ (_37588_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _87409_ (_37589_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _87410_ (_37590_, _37589_, _37588_);
  and _87411_ (_37591_, _20223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _87412_ (_37593_, \oc8051_golden_model_1.P0 [2], _39438_);
  or _87413_ (_37594_, _37593_, _37591_);
  or _87414_ (_37595_, _37594_, _37590_);
  and _87415_ (_37596_, \oc8051_golden_model_1.P0 [0], _39327_);
  and _87416_ (_37597_, _19980_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or _87417_ (_37598_, _37597_, _37596_);
  and _87418_ (_37599_, _20107_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _87419_ (_37600_, \oc8051_golden_model_1.P0 [1], _39422_);
  or _87420_ (_37601_, _37600_, _37599_);
  or _87421_ (_37602_, _37601_, _37598_);
  or _87422_ (_37604_, _37602_, _37595_);
  or _87423_ (_37605_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand _87424_ (_37606_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _87425_ (_37607_, _37606_, _37605_);
  or _87426_ (_37608_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand _87427_ (_37609_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _87428_ (_37610_, _37609_, _37608_);
  or _87429_ (_37611_, _37610_, _37607_);
  and _87430_ (_37612_, _09234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _87431_ (_37613_, \oc8051_golden_model_1.P0 [7], _39151_);
  or _87432_ (_37615_, _37613_, _37612_);
  nand _87433_ (_37616_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _87434_ (_37617_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _87435_ (_37618_, _37617_, _37616_);
  or _87436_ (_37619_, _37618_, _37615_);
  or _87437_ (_37620_, _37619_, _37611_);
  or _87438_ (_37621_, _37620_, _37604_);
  and _87439_ (property_invalid_p0, _37621_, _37418_);
  or _87440_ (_37622_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nand _87441_ (_37623_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _87442_ (_37625_, _37623_, _37622_);
  or _87443_ (_37626_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand _87444_ (_37627_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _87445_ (_37628_, _37627_, _37626_);
  or _87446_ (_37629_, _37628_, _37625_);
  and _87447_ (_37630_, \oc8051_golden_model_1.IRAM[0] [0], _40890_);
  and _87448_ (_37631_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _87449_ (_37632_, _37631_, _37630_);
  and _87450_ (_37633_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _87451_ (_37634_, \oc8051_golden_model_1.IRAM[0] [1], _40903_);
  or _87452_ (_37636_, _37634_, _37633_);
  or _87453_ (_37637_, _37636_, _37632_);
  or _87454_ (_37638_, _37637_, _37629_);
  or _87455_ (_37639_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand _87456_ (_37640_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and _87457_ (_37641_, _37640_, _37639_);
  or _87458_ (_37642_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand _87459_ (_37643_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _87460_ (_37644_, _37643_, _37642_);
  or _87461_ (_37645_, _37644_, _37641_);
  or _87462_ (_37647_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand _87463_ (_37648_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and _87464_ (_37649_, _37648_, _37647_);
  or _87465_ (_37650_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand _87466_ (_37651_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _87467_ (_37652_, _37651_, _37650_);
  or _87468_ (_37653_, _37652_, _37649_);
  or _87469_ (_37654_, _37653_, _37645_);
  or _87470_ (_37655_, _37654_, _37638_);
  or _87471_ (_37656_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand _87472_ (_37658_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and _87473_ (_37659_, _37658_, _37656_);
  or _87474_ (_37660_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand _87475_ (_37661_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _87476_ (_37662_, _37661_, _37660_);
  or _87477_ (_37663_, _37662_, _37659_);
  or _87478_ (_37664_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand _87479_ (_37665_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _87480_ (_37666_, _37665_, _37664_);
  or _87481_ (_37667_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nand _87482_ (_37669_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and _87483_ (_37670_, _37669_, _37667_);
  or _87484_ (_37671_, _37670_, _37666_);
  or _87485_ (_37672_, _37671_, _37663_);
  and _87486_ (_37673_, _05723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _87487_ (_37674_, \oc8051_golden_model_1.IRAM[1] [4], _40974_);
  or _87488_ (_37675_, _37674_, _37673_);
  and _87489_ (_37676_, \oc8051_golden_model_1.IRAM[1] [5], _40978_);
  and _87490_ (_37677_, _05415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _87491_ (_37678_, _37677_, _37676_);
  or _87492_ (_37680_, _37678_, _37675_);
  or _87493_ (_37681_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand _87494_ (_37682_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and _87495_ (_37683_, _37682_, _37681_);
  or _87496_ (_37684_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nand _87497_ (_37685_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _87498_ (_37686_, _37685_, _37684_);
  or _87499_ (_37687_, _37686_, _37683_);
  or _87500_ (_37688_, _37687_, _37680_);
  or _87501_ (_37689_, _37688_, _37672_);
  or _87502_ (_37691_, _37689_, _37655_);
  or _87503_ (_37692_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand _87504_ (_37693_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and _87505_ (_37694_, _37693_, _37692_);
  or _87506_ (_37695_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand _87507_ (_37696_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _87508_ (_37697_, _37696_, _37695_);
  or _87509_ (_37698_, _37697_, _37694_);
  or _87510_ (_37699_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nand _87511_ (_37700_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and _87512_ (_37702_, _37700_, _37699_);
  and _87513_ (_37703_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _87514_ (_37704_, \oc8051_golden_model_1.IRAM[2] [2], _40993_);
  or _87515_ (_37705_, _37704_, _37703_);
  or _87516_ (_37706_, _37705_, _37702_);
  or _87517_ (_37707_, _37706_, _37698_);
  and _87518_ (_37708_, _05729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _87519_ (_37709_, \oc8051_golden_model_1.IRAM[2] [4], _40998_);
  or _87520_ (_37710_, _37709_, _37708_);
  and _87521_ (_37711_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _87522_ (_37713_, \oc8051_golden_model_1.IRAM[2] [5], _41001_);
  or _87523_ (_37714_, _37713_, _37711_);
  or _87524_ (_37715_, _37714_, _37710_);
  or _87525_ (_37716_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nand _87526_ (_37717_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _87527_ (_37718_, _37717_, _37716_);
  and _87528_ (_37719_, \oc8051_golden_model_1.IRAM[2] [7], _41006_);
  and _87529_ (_37720_, _05152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _87530_ (_37721_, _37720_, _37719_);
  or _87531_ (_37722_, _37721_, _37718_);
  or _87532_ (_37724_, _37722_, _37715_);
  or _87533_ (_37725_, _37724_, _37707_);
  and _87534_ (_37726_, \oc8051_golden_model_1.IRAM[3] [2], _41016_);
  and _87535_ (_37727_, _04825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _87536_ (_37728_, _37727_, _37726_);
  nand _87537_ (_37729_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _87538_ (_37730_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and _87539_ (_37731_, _37730_, _37729_);
  or _87540_ (_37732_, _37731_, _37728_);
  and _87541_ (_37733_, _04569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and _87542_ (_37735_, \oc8051_golden_model_1.IRAM[3] [0], _41010_);
  or _87543_ (_37736_, _37735_, _37733_);
  and _87544_ (_37737_, \oc8051_golden_model_1.IRAM[3] [1], _41013_);
  and _87545_ (_37738_, _04352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _87546_ (_37739_, _37738_, _37737_);
  or _87547_ (_37740_, _37739_, _37736_);
  or _87548_ (_37741_, _37740_, _37732_);
  or _87549_ (_37742_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand _87550_ (_37743_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and _87551_ (_37744_, _37743_, _37742_);
  and _87552_ (_37746_, _05150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and _87553_ (_37747_, \oc8051_golden_model_1.IRAM[3] [7], _40758_);
  or _87554_ (_37748_, _37747_, _37746_);
  or _87555_ (_37749_, _37748_, _37744_);
  or _87556_ (_37750_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand _87557_ (_37751_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and _87558_ (_37752_, _37751_, _37750_);
  or _87559_ (_37753_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand _87560_ (_37754_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and _87561_ (_37755_, _37754_, _37753_);
  or _87562_ (_37757_, _37755_, _37752_);
  or _87563_ (_37758_, _37757_, _37749_);
  or _87564_ (_37759_, _37758_, _37741_);
  or _87565_ (_37760_, _37759_, _37725_);
  or _87566_ (_37761_, _37760_, _37691_);
  and _87567_ (_37762_, _04584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and _87568_ (_37763_, \oc8051_golden_model_1.IRAM[4] [0], _41033_);
  or _87569_ (_37764_, _37763_, _37762_);
  and _87570_ (_37765_, \oc8051_golden_model_1.IRAM[4] [1], _41036_);
  and _87571_ (_37766_, _04368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _87572_ (_37768_, _37766_, _37765_);
  or _87573_ (_37769_, _37768_, _37764_);
  or _87574_ (_37770_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand _87575_ (_37771_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and _87576_ (_37772_, _37771_, _37770_);
  nand _87577_ (_37773_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _87578_ (_37774_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and _87579_ (_37775_, _37774_, _37773_);
  or _87580_ (_37776_, _37775_, _37772_);
  or _87581_ (_37777_, _37776_, _37769_);
  or _87582_ (_37779_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand _87583_ (_37780_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and _87584_ (_37781_, _37780_, _37779_);
  or _87585_ (_37782_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand _87586_ (_37783_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and _87587_ (_37784_, _37783_, _37782_);
  or _87588_ (_37785_, _37784_, _37781_);
  or _87589_ (_37786_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand _87590_ (_37787_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and _87591_ (_37788_, _37787_, _37786_);
  nand _87592_ (_37790_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _87593_ (_37791_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and _87594_ (_37792_, _37791_, _37790_);
  or _87595_ (_37793_, _37792_, _37788_);
  or _87596_ (_37794_, _37793_, _37785_);
  or _87597_ (_37795_, _37794_, _37777_);
  or _87598_ (_37796_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand _87599_ (_37797_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _87600_ (_37798_, _37797_, _37796_);
  nand _87601_ (_37799_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _87602_ (_37801_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and _87603_ (_37802_, _37801_, _37799_);
  or _87604_ (_37803_, _37802_, _37798_);
  or _87605_ (_37804_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand _87606_ (_37805_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _87607_ (_37806_, _37805_, _37804_);
  or _87608_ (_37807_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand _87609_ (_37808_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and _87610_ (_37809_, _37808_, _37807_);
  or _87611_ (_37810_, _37809_, _37806_);
  or _87612_ (_37812_, _37810_, _37803_);
  or _87613_ (_37813_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand _87614_ (_37814_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _87615_ (_37815_, _37814_, _37813_);
  nand _87616_ (_37816_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or _87617_ (_37817_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _87618_ (_37818_, _37817_, _37816_);
  or _87619_ (_37819_, _37818_, _37815_);
  and _87620_ (_37820_, _05743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _87621_ (_37821_, \oc8051_golden_model_1.IRAM[5] [4], _41063_);
  or _87622_ (_37823_, _37821_, _37820_);
  and _87623_ (_37824_, _05435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _87624_ (_37825_, \oc8051_golden_model_1.IRAM[5] [5], _41066_);
  or _87625_ (_37826_, _37825_, _37824_);
  or _87626_ (_37827_, _37826_, _37823_);
  or _87627_ (_37828_, _37827_, _37819_);
  or _87628_ (_37829_, _37828_, _37812_);
  or _87629_ (_37830_, _37829_, _37795_);
  nand _87630_ (_37831_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _87631_ (_37832_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _87632_ (_37834_, _37832_, _37831_);
  and _87633_ (_37835_, \oc8051_golden_model_1.IRAM[6] [2], _41080_);
  and _87634_ (_37836_, _04835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _87635_ (_37837_, _37836_, _37835_);
  or _87636_ (_37838_, _37837_, _37834_);
  or _87637_ (_37839_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand _87638_ (_37840_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _87639_ (_37841_, _37840_, _37839_);
  or _87640_ (_37842_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand _87641_ (_37843_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and _87642_ (_37845_, _37843_, _37842_);
  or _87643_ (_37846_, _37845_, _37841_);
  or _87644_ (_37847_, _37846_, _37838_);
  and _87645_ (_37848_, _05160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and _87646_ (_37849_, \oc8051_golden_model_1.IRAM[6] [7], _41094_);
  or _87647_ (_37850_, _37849_, _37848_);
  nand _87648_ (_37851_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _87649_ (_37852_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _87650_ (_37853_, _37852_, _37851_);
  or _87651_ (_37854_, _37853_, _37850_);
  and _87652_ (_37856_, _05737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _87653_ (_37857_, \oc8051_golden_model_1.IRAM[6] [4], _41085_);
  or _87654_ (_37858_, _37857_, _37856_);
  and _87655_ (_37859_, \oc8051_golden_model_1.IRAM[6] [5], _41088_);
  and _87656_ (_37860_, _05429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _87657_ (_37861_, _37860_, _37859_);
  or _87658_ (_37862_, _37861_, _37858_);
  or _87659_ (_37863_, _37862_, _37854_);
  or _87660_ (_37864_, _37863_, _37847_);
  and _87661_ (_37865_, _04362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _87662_ (_37867_, \oc8051_golden_model_1.IRAM[7] [1], _41101_);
  or _87663_ (_37868_, _37867_, _37865_);
  and _87664_ (_37869_, _04578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and _87665_ (_37870_, \oc8051_golden_model_1.IRAM[7] [0], _41098_);
  or _87666_ (_37871_, _37870_, _37869_);
  or _87667_ (_37872_, _37871_, _37868_);
  and _87668_ (_37873_, _04833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and _87669_ (_37874_, \oc8051_golden_model_1.IRAM[7] [2], _41104_);
  or _87670_ (_37875_, _37874_, _37873_);
  nand _87671_ (_37876_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _87672_ (_37878_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _87673_ (_37879_, _37878_, _37876_);
  or _87674_ (_37880_, _37879_, _37875_);
  or _87675_ (_37881_, _37880_, _37872_);
  or _87676_ (_37882_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand _87677_ (_37883_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and _87678_ (_37884_, _37883_, _37882_);
  or _87679_ (_37885_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand _87680_ (_37886_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and _87681_ (_37887_, _37886_, _37885_);
  or _87682_ (_37889_, _37887_, _37884_);
  nand _87683_ (_37890_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _87684_ (_37891_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and _87685_ (_37892_, _37891_, _37890_);
  and _87686_ (_37893_, _05158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and _87687_ (_37894_, \oc8051_golden_model_1.IRAM[7] [7], _40794_);
  or _87688_ (_37895_, _37894_, _37893_);
  or _87689_ (_37896_, _37895_, _37892_);
  or _87690_ (_37897_, _37896_, _37889_);
  or _87691_ (_37898_, _37897_, _37881_);
  or _87692_ (_37900_, _37898_, _37864_);
  or _87693_ (_37901_, _37900_, _37830_);
  or _87694_ (_37902_, _37901_, _37761_);
  and _87695_ (_37903_, _04599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _87696_ (_37904_, \oc8051_golden_model_1.IRAM[8] [0], _41121_);
  or _87697_ (_37905_, _37904_, _37903_);
  and _87698_ (_37906_, \oc8051_golden_model_1.IRAM[8] [1], _41124_);
  and _87699_ (_37907_, _04385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _87700_ (_37908_, _37907_, _37906_);
  or _87701_ (_37909_, _37908_, _37905_);
  or _87702_ (_37911_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand _87703_ (_37912_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _87704_ (_37913_, _37912_, _37911_);
  nand _87705_ (_37914_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _87706_ (_37915_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _87707_ (_37916_, _37915_, _37914_);
  or _87708_ (_37917_, _37916_, _37913_);
  or _87709_ (_37918_, _37917_, _37909_);
  or _87710_ (_37919_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand _87711_ (_37920_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _87712_ (_37922_, _37920_, _37919_);
  or _87713_ (_37923_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand _87714_ (_37924_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _87715_ (_37925_, _37924_, _37923_);
  or _87716_ (_37926_, _37925_, _37922_);
  or _87717_ (_37927_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand _87718_ (_37928_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _87719_ (_37929_, _37928_, _37927_);
  nand _87720_ (_37930_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or _87721_ (_37931_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _87722_ (_37933_, _37931_, _37930_);
  or _87723_ (_37934_, _37933_, _37929_);
  or _87724_ (_37935_, _37934_, _37926_);
  or _87725_ (_37936_, _37935_, _37918_);
  or _87726_ (_37937_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand _87727_ (_37938_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _87728_ (_37939_, _37938_, _37937_);
  nand _87729_ (_37940_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _87730_ (_37941_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _87731_ (_37942_, _37941_, _37940_);
  or _87732_ (_37944_, _37942_, _37939_);
  or _87733_ (_37945_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand _87734_ (_37946_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _87735_ (_37947_, _37946_, _37945_);
  or _87736_ (_37948_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand _87737_ (_37949_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _87738_ (_37950_, _37949_, _37948_);
  or _87739_ (_37951_, _37950_, _37947_);
  or _87740_ (_37952_, _37951_, _37944_);
  and _87741_ (_37953_, _05449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _87742_ (_37955_, \oc8051_golden_model_1.IRAM[9] [5], _41155_);
  or _87743_ (_37956_, _37955_, _37953_);
  and _87744_ (_37957_, _05757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and _87745_ (_37958_, \oc8051_golden_model_1.IRAM[9] [4], _41152_);
  or _87746_ (_37959_, _37958_, _37957_);
  or _87747_ (_37960_, _37959_, _37956_);
  or _87748_ (_37961_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand _87749_ (_37962_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _87750_ (_37963_, _37962_, _37961_);
  nand _87751_ (_37964_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _87752_ (_37966_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _87753_ (_37967_, _37966_, _37964_);
  or _87754_ (_37968_, _37967_, _37963_);
  or _87755_ (_37969_, _37968_, _37960_);
  or _87756_ (_37970_, _37969_, _37952_);
  or _87757_ (_37971_, _37970_, _37936_);
  and _87758_ (_37972_, _04851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and _87759_ (_37973_, \oc8051_golden_model_1.IRAM[10] [2], _41168_);
  or _87760_ (_37974_, _37973_, _37972_);
  nand _87761_ (_37975_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _87762_ (_37976_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and _87763_ (_37977_, _37976_, _37975_);
  or _87764_ (_37978_, _37977_, _37974_);
  or _87765_ (_37979_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nand _87766_ (_37980_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _87767_ (_37981_, _37980_, _37979_);
  or _87768_ (_37982_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nand _87769_ (_37983_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and _87770_ (_37984_, _37983_, _37982_);
  or _87771_ (_37985_, _37984_, _37981_);
  or _87772_ (_37987_, _37985_, _37978_);
  and _87773_ (_37988_, \oc8051_golden_model_1.IRAM[10] [7], _40831_);
  and _87774_ (_37989_, _05176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _87775_ (_37990_, _37989_, _37988_);
  nand _87776_ (_37991_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _87777_ (_37992_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and _87778_ (_37993_, _37992_, _37991_);
  or _87779_ (_37994_, _37993_, _37990_);
  and _87780_ (_37995_, _05752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and _87781_ (_37996_, \oc8051_golden_model_1.IRAM[10] [4], _41174_);
  or _87782_ (_37998_, _37996_, _37995_);
  and _87783_ (_37999_, \oc8051_golden_model_1.IRAM[10] [5], _41177_);
  and _87784_ (_38000_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _87785_ (_38001_, _38000_, _37999_);
  or _87786_ (_38002_, _38001_, _37998_);
  or _87787_ (_38003_, _38002_, _37994_);
  or _87788_ (_38004_, _38003_, _37987_);
  and _87789_ (_38005_, _04594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _87790_ (_38006_, \oc8051_golden_model_1.IRAM[11] [0], _41186_);
  or _87791_ (_38007_, _38006_, _38005_);
  and _87792_ (_38009_, \oc8051_golden_model_1.IRAM[11] [1], _41189_);
  and _87793_ (_38010_, _04380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _87794_ (_38011_, _38010_, _38009_);
  or _87795_ (_38012_, _38011_, _38007_);
  and _87796_ (_38013_, \oc8051_golden_model_1.IRAM[11] [2], _41192_);
  and _87797_ (_38014_, _04849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _87798_ (_38015_, _38014_, _38013_);
  nand _87799_ (_38016_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _87800_ (_38017_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _87801_ (_38018_, _38017_, _38016_);
  or _87802_ (_38020_, _38018_, _38015_);
  or _87803_ (_38021_, _38020_, _38012_);
  or _87804_ (_38022_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand _87805_ (_38023_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _87806_ (_38024_, _38023_, _38022_);
  or _87807_ (_38025_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand _87808_ (_38026_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _87809_ (_38027_, _38026_, _38025_);
  or _87810_ (_38028_, _38027_, _38024_);
  and _87811_ (_38029_, _05174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _87812_ (_38031_, \oc8051_golden_model_1.IRAM[11] [7], _41204_);
  or _87813_ (_38032_, _38031_, _38029_);
  nand _87814_ (_38033_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _87815_ (_38034_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _87816_ (_38035_, _38034_, _38033_);
  or _87817_ (_38036_, _38035_, _38032_);
  or _87818_ (_38037_, _38036_, _38028_);
  or _87819_ (_38038_, _38037_, _38021_);
  or _87820_ (_38039_, _38038_, _38004_);
  or _87821_ (_38040_, _38039_, _37971_);
  or _87822_ (_38042_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand _87823_ (_38043_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _87824_ (_38044_, _38043_, _38042_);
  nand _87825_ (_38045_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or _87826_ (_38046_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _87827_ (_38047_, _38046_, _38045_);
  or _87828_ (_38048_, _38047_, _38044_);
  and _87829_ (_38049_, \oc8051_golden_model_1.IRAM[12] [1], _41217_);
  and _87830_ (_38050_, _04397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _87831_ (_38051_, _38050_, _38049_);
  and _87832_ (_38053_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and _87833_ (_38054_, \oc8051_golden_model_1.IRAM[12] [0], _41210_);
  or _87834_ (_38055_, _38054_, _38053_);
  or _87835_ (_38056_, _38055_, _38051_);
  or _87836_ (_38057_, _38056_, _38048_);
  or _87837_ (_38058_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand _87838_ (_38059_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _87839_ (_38060_, _38059_, _38058_);
  nand _87840_ (_38061_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _87841_ (_38062_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and _87842_ (_38064_, _38062_, _38061_);
  or _87843_ (_38065_, _38064_, _38060_);
  or _87844_ (_38066_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand _87845_ (_38067_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _87846_ (_38068_, _38067_, _38066_);
  or _87847_ (_38069_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand _87848_ (_38070_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _87849_ (_38071_, _38070_, _38069_);
  or _87850_ (_38072_, _38071_, _38068_);
  or _87851_ (_38073_, _38072_, _38065_);
  or _87852_ (_38075_, _38073_, _38057_);
  or _87853_ (_38076_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand _87854_ (_38077_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _87855_ (_38078_, _38077_, _38076_);
  or _87856_ (_38079_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand _87857_ (_38080_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _87858_ (_38081_, _38080_, _38079_);
  or _87859_ (_38082_, _38081_, _38078_);
  or _87860_ (_38083_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand _87861_ (_38084_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _87862_ (_38086_, _38084_, _38083_);
  nand _87863_ (_38087_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _87864_ (_38088_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _87865_ (_38089_, _38088_, _38087_);
  or _87866_ (_38090_, _38089_, _38086_);
  or _87867_ (_38091_, _38090_, _38082_);
  and _87868_ (_38092_, _05769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and _87869_ (_38093_, \oc8051_golden_model_1.IRAM[13] [4], _41267_);
  or _87870_ (_38094_, _38093_, _38092_);
  and _87871_ (_38095_, \oc8051_golden_model_1.IRAM[13] [5], _41270_);
  and _87872_ (_38097_, _05461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _87873_ (_38098_, _38097_, _38095_);
  or _87874_ (_38099_, _38098_, _38094_);
  or _87875_ (_38100_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand _87876_ (_38101_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _87877_ (_38102_, _38101_, _38100_);
  nand _87878_ (_38103_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _87879_ (_38104_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _87880_ (_38105_, _38104_, _38103_);
  or _87881_ (_38106_, _38105_, _38102_);
  or _87882_ (_38108_, _38106_, _38099_);
  or _87883_ (_38109_, _38108_, _38091_);
  or _87884_ (_38110_, _38109_, _38075_);
  or _87885_ (_38111_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nand _87886_ (_38112_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _87887_ (_38113_, _38112_, _38111_);
  or _87888_ (_38114_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nand _87889_ (_38115_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and _87890_ (_38116_, _38115_, _38114_);
  or _87891_ (_38117_, _38116_, _38113_);
  and _87892_ (_38119_, \oc8051_golden_model_1.IRAM[14] [2], _41283_);
  and _87893_ (_38120_, _04863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _87894_ (_38121_, _38120_, _38119_);
  nand _87895_ (_38122_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _87896_ (_38123_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and _87897_ (_38124_, _38123_, _38122_);
  or _87898_ (_38125_, _38124_, _38121_);
  or _87899_ (_38126_, _38125_, _38117_);
  and _87900_ (_38127_, \oc8051_golden_model_1.IRAM[14] [5], _41292_);
  and _87901_ (_38128_, _05456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _87902_ (_38130_, _38128_, _38127_);
  and _87903_ (_38131_, _05764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and _87904_ (_38132_, \oc8051_golden_model_1.IRAM[14] [4], _41289_);
  or _87905_ (_38133_, _38132_, _38131_);
  or _87906_ (_38134_, _38133_, _38130_);
  and _87907_ (_38135_, _05190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _87908_ (_38136_, \oc8051_golden_model_1.IRAM[14] [7], _40842_);
  or _87909_ (_38137_, _38136_, _38135_);
  nand _87910_ (_38138_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _87911_ (_38139_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and _87912_ (_38141_, _38139_, _38138_);
  or _87913_ (_38142_, _38141_, _38137_);
  or _87914_ (_38143_, _38142_, _38134_);
  or _87915_ (_38144_, _38143_, _38126_);
  and _87916_ (_38145_, _04861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _87917_ (_38146_, \oc8051_golden_model_1.IRAM[15] [2], _41306_);
  or _87918_ (_38147_, _38146_, _38145_);
  nand _87919_ (_38148_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _87920_ (_38149_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _87921_ (_38150_, _38149_, _38148_);
  or _87922_ (_38152_, _38150_, _38147_);
  and _87923_ (_38153_, _04606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _87924_ (_38154_, \oc8051_golden_model_1.IRAM[15] [0], _41300_);
  or _87925_ (_38155_, _38154_, _38153_);
  and _87926_ (_38156_, _04392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _87927_ (_38157_, \oc8051_golden_model_1.IRAM[15] [1], _41303_);
  or _87928_ (_38158_, _38157_, _38156_);
  or _87929_ (_38159_, _38158_, _38155_);
  or _87930_ (_38160_, _38159_, _38152_);
  and _87931_ (_38161_, \oc8051_golden_model_1.IRAM[15] [7], _40873_);
  and _87932_ (_38163_, _05188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _87933_ (_38164_, _38163_, _38161_);
  nand _87934_ (_38165_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _87935_ (_38166_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _87936_ (_38167_, _38166_, _38165_);
  or _87937_ (_38168_, _38167_, _38164_);
  or _87938_ (_38169_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand _87939_ (_38170_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _87940_ (_38171_, _38170_, _38169_);
  or _87941_ (_38172_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand _87942_ (_38174_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _87943_ (_38175_, _38174_, _38172_);
  or _87944_ (_38176_, _38175_, _38171_);
  or _87945_ (_38177_, _38176_, _38168_);
  or _87946_ (_38178_, _38177_, _38160_);
  or _87947_ (_38179_, _38178_, _38144_);
  or _87948_ (_38180_, _38179_, _38110_);
  or _87949_ (_38181_, _38180_, _38040_);
  or _87950_ (_38182_, _38181_, _37902_);
  and _87951_ (property_invalid_iram, _38182_, _37418_);
  nand _87952_ (_38184_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _87953_ (_38185_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _87954_ (_38186_, _38185_, _38184_);
  and _87955_ (_38187_, _17923_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor _87956_ (_38188_, _17923_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _87957_ (_38189_, _38188_, _38187_);
  or _87958_ (_38190_, _38189_, _38186_);
  nor _87959_ (_38191_, _17740_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _87960_ (_38192_, _17740_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _87961_ (_38193_, _38192_, _38191_);
  and _87962_ (_38195_, _17829_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor _87963_ (_38196_, _17829_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _87964_ (_38197_, _38196_, _38195_);
  or _87965_ (_38198_, _38197_, _38193_);
  or _87966_ (_38199_, _38198_, _38190_);
  or _87967_ (_38200_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand _87968_ (_38201_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _87969_ (_38202_, _38201_, _38200_);
  or _87970_ (_38203_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand _87971_ (_38204_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _87972_ (_38206_, _38204_, _38203_);
  or _87973_ (_38207_, _38206_, _38202_);
  and _87974_ (_38208_, _08918_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor _87975_ (_38209_, _08918_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _87976_ (_38210_, _38209_, _38208_);
  nand _87977_ (_38211_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _87978_ (_38212_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _87979_ (_38213_, _38212_, _38211_);
  or _87980_ (_38214_, _38213_, _38210_);
  or _87981_ (_38215_, _38214_, _38207_);
  or _87982_ (_38217_, _38215_, _38199_);
  and _87983_ (property_invalid_dph, _38217_, _37418_);
  nand _87984_ (_38218_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or _87985_ (_38219_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _87986_ (_38220_, _38219_, _38218_);
  and _87987_ (_38221_, _17271_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _87988_ (_38222_, \oc8051_golden_model_1.DPL [2], _38799_);
  or _87989_ (_38223_, _38222_, _38221_);
  or _87990_ (_38224_, _38223_, _38220_);
  and _87991_ (_38225_, \oc8051_golden_model_1.DPL [0], _38791_);
  and _87992_ (_38227_, _17089_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or _87993_ (_38228_, _38227_, _38225_);
  and _87994_ (_38229_, _17177_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _87995_ (_38230_, \oc8051_golden_model_1.DPL [1], _38795_);
  or _87996_ (_38231_, _38230_, _38229_);
  or _87997_ (_38232_, _38231_, _38228_);
  or _87998_ (_38233_, _38232_, _38224_);
  or _87999_ (_38234_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand _88000_ (_38235_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _88001_ (_38236_, _38235_, _38234_);
  or _88002_ (_38238_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand _88003_ (_38239_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _88004_ (_38240_, _38239_, _38238_);
  or _88005_ (_38241_, _38240_, _38236_);
  and _88006_ (_38242_, _08821_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _88007_ (_38243_, \oc8051_golden_model_1.DPL [7], _38590_);
  or _88008_ (_38244_, _38243_, _38242_);
  nand _88009_ (_38245_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or _88010_ (_38246_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _88011_ (_38247_, _38246_, _38245_);
  or _88012_ (_38249_, _38247_, _38244_);
  or _88013_ (_38250_, _38249_, _38241_);
  or _88014_ (_38251_, _38250_, _38233_);
  and _88015_ (property_invalid_dpl, _38251_, _37418_);
  nand _88016_ (_38252_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _88017_ (_38253_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _88018_ (_38254_, _38253_, _38252_);
  and _88019_ (_38255_, _07426_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _88020_ (_38256_, \oc8051_golden_model_1.B [2], _30599_);
  or _88021_ (_38257_, _38256_, _38255_);
  or _88022_ (_38259_, _38257_, _38254_);
  and _88023_ (_38260_, \oc8051_golden_model_1.B [0], _29264_);
  and _88024_ (_38261_, _07418_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _88025_ (_38262_, _38261_, _38260_);
  and _88026_ (_38263_, _07412_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _88027_ (_38264_, \oc8051_golden_model_1.B [1], _29926_);
  or _88028_ (_38265_, _38264_, _38263_);
  or _88029_ (_38266_, _38265_, _38262_);
  or _88030_ (_38267_, _38266_, _38259_);
  or _88031_ (_38268_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _88032_ (_38270_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _88033_ (_38271_, _38270_, _38268_);
  or _88034_ (_38272_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _88035_ (_38273_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _88036_ (_38274_, _38273_, _38272_);
  or _88037_ (_38275_, _38274_, _38271_);
  and _88038_ (_38276_, _06826_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _88039_ (_38277_, \oc8051_golden_model_1.B [7], _28098_);
  or _88040_ (_38278_, _38277_, _38276_);
  nand _88041_ (_38279_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _88042_ (_38281_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _88043_ (_38282_, _38281_, _38279_);
  or _88044_ (_38283_, _38282_, _38278_);
  or _88045_ (_38284_, _38283_, _38275_);
  or _88046_ (_38285_, _38284_, _38267_);
  and _88047_ (property_invalid_b_reg, _38285_, _37418_);
  nand _88048_ (_38286_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _88049_ (_38287_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _88050_ (_38288_, _38287_, _38286_);
  and _88051_ (_38289_, _07584_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _88052_ (_38291_, \oc8051_golden_model_1.ACC [2], _39082_);
  or _88053_ (_38292_, _38291_, _38289_);
  or _88054_ (_38293_, _38292_, _38288_);
  nor _88055_ (_38294_, _03274_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _88056_ (_38295_, _03274_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _88057_ (_38296_, _38295_, _38294_);
  and _88058_ (_38297_, _03335_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _88059_ (_38298_, _03335_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _88060_ (_38299_, _38298_, _38297_);
  or _88061_ (_38300_, _38299_, _38296_);
  or _88062_ (_38302_, _38300_, _38293_);
  or _88063_ (_38303_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _88064_ (_38304_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _88065_ (_38305_, _38304_, _38303_);
  or _88066_ (_38306_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _88067_ (_38307_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _88068_ (_38308_, _38307_, _38306_);
  or _88069_ (_38309_, _38308_, _38305_);
  and _88070_ (_38310_, _07433_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _88071_ (_38311_, _07433_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _88072_ (_38313_, _38311_, _38310_);
  nand _88073_ (_38314_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _88074_ (_38315_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _88075_ (_38316_, _38315_, _38314_);
  or _88076_ (_38317_, _38316_, _38313_);
  or _88077_ (_38318_, _38317_, _38309_);
  or _88078_ (_38319_, _38318_, _38302_);
  and _88079_ (property_invalid_acc, _38319_, _37418_);
  and _88080_ (_38320_, _32793_, _43931_);
  nor _88081_ (_38321_, _32793_, _43931_);
  and _88082_ (_38323_, _33139_, _43935_);
  nor _88083_ (_38324_, _33139_, _43935_);
  and _88084_ (_38325_, _33488_, _43939_);
  and _88085_ (_38326_, _35539_, _38549_);
  nor _88086_ (_38327_, _35539_, _38549_);
  nor _88087_ (_38328_, _11981_, _38571_);
  nor _88088_ (_38329_, _36772_, _38535_);
  and _88089_ (_38330_, _11981_, _38571_);
  or _88090_ (_38331_, _38330_, _38329_);
  or _88091_ (_38332_, _38331_, _38328_);
  nand _88092_ (_38334_, _35205_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _88093_ (_38335_, _35205_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _88094_ (_38336_, _38335_, _38334_);
  nor _88095_ (_38337_, _36160_, _38539_);
  and _88096_ (_38338_, _35846_, _38554_);
  nor _88097_ (_38339_, _35846_, _38554_);
  and _88098_ (_38340_, _36468_, _38560_);
  nand _88099_ (_38341_, _32414_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _88100_ (_38342_, _32414_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _88101_ (_38343_, _38342_, _38341_);
  nor _88102_ (_38345_, _36468_, _38560_);
  or _88103_ (_38346_, _38345_, _38343_);
  or _88104_ (_38347_, _38346_, _38340_);
  and _88105_ (_38348_, _37080_, _38566_);
  nor _88106_ (_38349_, _37080_, _38566_);
  or _88107_ (_38350_, _38349_, _38348_);
  or _88108_ (_38351_, _38350_, _38347_);
  or _88109_ (_38352_, _38351_, _38339_);
  or _88110_ (_38353_, _38352_, _38338_);
  or _88111_ (_38354_, _38353_, _38337_);
  and _88112_ (_38356_, _36160_, _38539_);
  and _88113_ (_38357_, _36772_, _38535_);
  or _88114_ (_38358_, _38357_, _38356_);
  or _88115_ (_38359_, _38358_, _38354_);
  or _88116_ (_38360_, _38359_, _38336_);
  or _88117_ (_38361_, _38360_, _38332_);
  or _88118_ (_38362_, _38361_, _38327_);
  or _88119_ (_38363_, _38362_, _38326_);
  or _88120_ (_38364_, _38363_, _38325_);
  or _88121_ (_38365_, _38364_, _38324_);
  or _88122_ (_38367_, _38365_, _38323_);
  nor _88123_ (_38368_, _34187_, _43947_);
  nor _88124_ (_38369_, _34887_, _43955_);
  and _88125_ (_38370_, _34187_, _43947_);
  or _88126_ (_38371_, _38370_, _38369_);
  or _88127_ (_38372_, _38371_, _38368_);
  nor _88128_ (_38373_, _33488_, _43939_);
  and _88129_ (_38374_, _33837_, _43943_);
  or _88130_ (_38375_, _38374_, _38373_);
  nor _88131_ (_38376_, _33837_, _43943_);
  and _88132_ (_38378_, _34887_, _43955_);
  or _88133_ (_38379_, _38378_, _38376_);
  or _88134_ (_38380_, _38379_, _38375_);
  or _88135_ (_38381_, _38380_, _38372_);
  or _88136_ (_38382_, _38381_, _38367_);
  nor _88137_ (_38383_, _34533_, _43951_);
  and _88138_ (_38384_, _34533_, _43951_);
  or _88139_ (_38385_, _38384_, _38383_);
  or _88140_ (_38386_, _38385_, _38382_);
  or _88141_ (_38387_, _38386_, _38321_);
  or _88142_ (_38389_, _38387_, _38320_);
  and _88143_ (property_invalid_pc, _38389_, _37350_);
  buf _88144_ (_01429_, _41806_);
  buf _88145_ (_01480_, _41806_);
  buf _88146_ (_01532_, _41806_);
  buf _88147_ (_01584_, _41806_);
  buf _88148_ (_01629_, _41806_);
  buf _88149_ (_01675_, _41806_);
  buf _88150_ (_01728_, _41806_);
  buf _88151_ (_01779_, _41806_);
  buf _88152_ (_01831_, _41806_);
  buf _88153_ (_01883_, _41806_);
  buf _88154_ (_01935_, _41806_);
  buf _88155_ (_01987_, _41806_);
  buf _88156_ (_02039_, _41806_);
  buf _88157_ (_02091_, _41806_);
  buf _88158_ (_02143_, _41806_);
  buf _88159_ (_02195_, _41806_);
  buf _88160_ (_38916_, _38813_);
  buf _88161_ (_38917_, _38814_);
  buf _88162_ (_38930_, _38813_);
  buf _88163_ (_38931_, _38814_);
  buf _88164_ (_39244_, _38832_);
  buf _88165_ (_39245_, _38834_);
  buf _88166_ (_39246_, _38835_);
  buf _88167_ (_39247_, _38836_);
  buf _88168_ (_39248_, _38837_);
  buf _88169_ (_39249_, _38838_);
  buf _88170_ (_39250_, _38840_);
  buf _88171_ (_39252_, _38841_);
  buf _88172_ (_39253_, _38842_);
  buf _88173_ (_39254_, _38843_);
  buf _88174_ (_39255_, _38844_);
  buf _88175_ (_39256_, _38846_);
  buf _88176_ (_39257_, _38847_);
  buf _88177_ (_39258_, _38848_);
  buf _88178_ (_39310_, _38832_);
  buf _88179_ (_39311_, _38834_);
  buf _88180_ (_39312_, _38835_);
  buf _88181_ (_39313_, _38836_);
  buf _88182_ (_39314_, _38837_);
  buf _88183_ (_39315_, _38838_);
  buf _88184_ (_39316_, _38840_);
  buf _88185_ (_39317_, _38841_);
  buf _88186_ (_39318_, _38842_);
  buf _88187_ (_39319_, _38843_);
  buf _88188_ (_39320_, _38844_);
  buf _88189_ (_39321_, _38846_);
  buf _88190_ (_39322_, _38847_);
  buf _88191_ (_39323_, _38848_);
  buf _88192_ (_39651_, _39617_);
  buf _88193_ (_39766_, _39617_);
  dff _88194_ (p0in_reg[0], _00002_[0], clk);
  dff _88195_ (p0in_reg[1], _00002_[1], clk);
  dff _88196_ (p0in_reg[2], _00002_[2], clk);
  dff _88197_ (p0in_reg[3], _00002_[3], clk);
  dff _88198_ (p0in_reg[4], _00002_[4], clk);
  dff _88199_ (p0in_reg[5], _00002_[5], clk);
  dff _88200_ (p0in_reg[6], _00002_[6], clk);
  dff _88201_ (p0in_reg[7], _00002_[7], clk);
  dff _88202_ (p1in_reg[0], _00003_[0], clk);
  dff _88203_ (p1in_reg[1], _00003_[1], clk);
  dff _88204_ (p1in_reg[2], _00003_[2], clk);
  dff _88205_ (p1in_reg[3], _00003_[3], clk);
  dff _88206_ (p1in_reg[4], _00003_[4], clk);
  dff _88207_ (p1in_reg[5], _00003_[5], clk);
  dff _88208_ (p1in_reg[6], _00003_[6], clk);
  dff _88209_ (p1in_reg[7], _00003_[7], clk);
  dff _88210_ (p2in_reg[0], _00004_[0], clk);
  dff _88211_ (p2in_reg[1], _00004_[1], clk);
  dff _88212_ (p2in_reg[2], _00004_[2], clk);
  dff _88213_ (p2in_reg[3], _00004_[3], clk);
  dff _88214_ (p2in_reg[4], _00004_[4], clk);
  dff _88215_ (p2in_reg[5], _00004_[5], clk);
  dff _88216_ (p2in_reg[6], _00004_[6], clk);
  dff _88217_ (p2in_reg[7], _00004_[7], clk);
  dff _88218_ (p3in_reg[0], _00005_[0], clk);
  dff _88219_ (p3in_reg[1], _00005_[1], clk);
  dff _88220_ (p3in_reg[2], _00005_[2], clk);
  dff _88221_ (p3in_reg[3], _00005_[3], clk);
  dff _88222_ (p3in_reg[4], _00005_[4], clk);
  dff _88223_ (p3in_reg[5], _00005_[5], clk);
  dff _88224_ (p3in_reg[6], _00005_[6], clk);
  dff _88225_ (p3in_reg[7], _00005_[7], clk);
  dff _88226_ (op0_cnst, _00001_, clk);
  dff _88227_ (inst_finished_r, _00000_, clk);
  dff _88228_ (property_invalid_psw_1_r, _00006_, clk);
  dff _88229_ (property_invalid_sp_1_r, _00007_, clk);
  dff _88230_ (\oc8051_gm_cxrom_1.cell0.data [0], _01433_, clk);
  dff _88231_ (\oc8051_gm_cxrom_1.cell0.data [1], _01437_, clk);
  dff _88232_ (\oc8051_gm_cxrom_1.cell0.data [2], _01441_, clk);
  dff _88233_ (\oc8051_gm_cxrom_1.cell0.data [3], _01444_, clk);
  dff _88234_ (\oc8051_gm_cxrom_1.cell0.data [4], _01448_, clk);
  dff _88235_ (\oc8051_gm_cxrom_1.cell0.data [5], _01452_, clk);
  dff _88236_ (\oc8051_gm_cxrom_1.cell0.data [6], _01456_, clk);
  dff _88237_ (\oc8051_gm_cxrom_1.cell0.data [7], _01426_, clk);
  dff _88238_ (\oc8051_gm_cxrom_1.cell0.valid , _01429_, clk);
  dff _88239_ (\oc8051_gm_cxrom_1.cell1.data [0], _01484_, clk);
  dff _88240_ (\oc8051_gm_cxrom_1.cell1.data [1], _01488_, clk);
  dff _88241_ (\oc8051_gm_cxrom_1.cell1.data [2], _01492_, clk);
  dff _88242_ (\oc8051_gm_cxrom_1.cell1.data [3], _01496_, clk);
  dff _88243_ (\oc8051_gm_cxrom_1.cell1.data [4], _01500_, clk);
  dff _88244_ (\oc8051_gm_cxrom_1.cell1.data [5], _01504_, clk);
  dff _88245_ (\oc8051_gm_cxrom_1.cell1.data [6], _01508_, clk);
  dff _88246_ (\oc8051_gm_cxrom_1.cell1.data [7], _01477_, clk);
  dff _88247_ (\oc8051_gm_cxrom_1.cell1.valid , _01480_, clk);
  dff _88248_ (\oc8051_gm_cxrom_1.cell10.data [0], _01939_, clk);
  dff _88249_ (\oc8051_gm_cxrom_1.cell10.data [1], _01943_, clk);
  dff _88250_ (\oc8051_gm_cxrom_1.cell10.data [2], _01947_, clk);
  dff _88251_ (\oc8051_gm_cxrom_1.cell10.data [3], _01951_, clk);
  dff _88252_ (\oc8051_gm_cxrom_1.cell10.data [4], _01955_, clk);
  dff _88253_ (\oc8051_gm_cxrom_1.cell10.data [5], _01959_, clk);
  dff _88254_ (\oc8051_gm_cxrom_1.cell10.data [6], _01963_, clk);
  dff _88255_ (\oc8051_gm_cxrom_1.cell10.data [7], _01932_, clk);
  dff _88256_ (\oc8051_gm_cxrom_1.cell10.valid , _01935_, clk);
  dff _88257_ (\oc8051_gm_cxrom_1.cell11.data [0], _01991_, clk);
  dff _88258_ (\oc8051_gm_cxrom_1.cell11.data [1], _01995_, clk);
  dff _88259_ (\oc8051_gm_cxrom_1.cell11.data [2], _01999_, clk);
  dff _88260_ (\oc8051_gm_cxrom_1.cell11.data [3], _02003_, clk);
  dff _88261_ (\oc8051_gm_cxrom_1.cell11.data [4], _02007_, clk);
  dff _88262_ (\oc8051_gm_cxrom_1.cell11.data [5], _02011_, clk);
  dff _88263_ (\oc8051_gm_cxrom_1.cell11.data [6], _02015_, clk);
  dff _88264_ (\oc8051_gm_cxrom_1.cell11.data [7], _01984_, clk);
  dff _88265_ (\oc8051_gm_cxrom_1.cell11.valid , _01987_, clk);
  dff _88266_ (\oc8051_gm_cxrom_1.cell12.data [0], _02043_, clk);
  dff _88267_ (\oc8051_gm_cxrom_1.cell12.data [1], _02047_, clk);
  dff _88268_ (\oc8051_gm_cxrom_1.cell12.data [2], _02051_, clk);
  dff _88269_ (\oc8051_gm_cxrom_1.cell12.data [3], _02055_, clk);
  dff _88270_ (\oc8051_gm_cxrom_1.cell12.data [4], _02059_, clk);
  dff _88271_ (\oc8051_gm_cxrom_1.cell12.data [5], _02063_, clk);
  dff _88272_ (\oc8051_gm_cxrom_1.cell12.data [6], _02067_, clk);
  dff _88273_ (\oc8051_gm_cxrom_1.cell12.data [7], _02036_, clk);
  dff _88274_ (\oc8051_gm_cxrom_1.cell12.valid , _02039_, clk);
  dff _88275_ (\oc8051_gm_cxrom_1.cell13.data [0], _02095_, clk);
  dff _88276_ (\oc8051_gm_cxrom_1.cell13.data [1], _02099_, clk);
  dff _88277_ (\oc8051_gm_cxrom_1.cell13.data [2], _02103_, clk);
  dff _88278_ (\oc8051_gm_cxrom_1.cell13.data [3], _02107_, clk);
  dff _88279_ (\oc8051_gm_cxrom_1.cell13.data [4], _02111_, clk);
  dff _88280_ (\oc8051_gm_cxrom_1.cell13.data [5], _02115_, clk);
  dff _88281_ (\oc8051_gm_cxrom_1.cell13.data [6], _02119_, clk);
  dff _88282_ (\oc8051_gm_cxrom_1.cell13.data [7], _02088_, clk);
  dff _88283_ (\oc8051_gm_cxrom_1.cell13.valid , _02091_, clk);
  dff _88284_ (\oc8051_gm_cxrom_1.cell14.data [0], _02147_, clk);
  dff _88285_ (\oc8051_gm_cxrom_1.cell14.data [1], _02151_, clk);
  dff _88286_ (\oc8051_gm_cxrom_1.cell14.data [2], _02155_, clk);
  dff _88287_ (\oc8051_gm_cxrom_1.cell14.data [3], _02159_, clk);
  dff _88288_ (\oc8051_gm_cxrom_1.cell14.data [4], _02163_, clk);
  dff _88289_ (\oc8051_gm_cxrom_1.cell14.data [5], _02167_, clk);
  dff _88290_ (\oc8051_gm_cxrom_1.cell14.data [6], _02171_, clk);
  dff _88291_ (\oc8051_gm_cxrom_1.cell14.data [7], _02140_, clk);
  dff _88292_ (\oc8051_gm_cxrom_1.cell14.valid , _02143_, clk);
  dff _88293_ (\oc8051_gm_cxrom_1.cell15.data [0], _02199_, clk);
  dff _88294_ (\oc8051_gm_cxrom_1.cell15.data [1], _02203_, clk);
  dff _88295_ (\oc8051_gm_cxrom_1.cell15.data [2], _02207_, clk);
  dff _88296_ (\oc8051_gm_cxrom_1.cell15.data [3], _02211_, clk);
  dff _88297_ (\oc8051_gm_cxrom_1.cell15.data [4], _02215_, clk);
  dff _88298_ (\oc8051_gm_cxrom_1.cell15.data [5], _02219_, clk);
  dff _88299_ (\oc8051_gm_cxrom_1.cell15.data [6], _02223_, clk);
  dff _88300_ (\oc8051_gm_cxrom_1.cell15.data [7], _02192_, clk);
  dff _88301_ (\oc8051_gm_cxrom_1.cell15.valid , _02195_, clk);
  dff _88302_ (\oc8051_gm_cxrom_1.cell2.data [0], _01536_, clk);
  dff _88303_ (\oc8051_gm_cxrom_1.cell2.data [1], _01540_, clk);
  dff _88304_ (\oc8051_gm_cxrom_1.cell2.data [2], _01544_, clk);
  dff _88305_ (\oc8051_gm_cxrom_1.cell2.data [3], _01548_, clk);
  dff _88306_ (\oc8051_gm_cxrom_1.cell2.data [4], _01552_, clk);
  dff _88307_ (\oc8051_gm_cxrom_1.cell2.data [5], _01555_, clk);
  dff _88308_ (\oc8051_gm_cxrom_1.cell2.data [6], _01559_, clk);
  dff _88309_ (\oc8051_gm_cxrom_1.cell2.data [7], _01529_, clk);
  dff _88310_ (\oc8051_gm_cxrom_1.cell2.valid , _01532_, clk);
  dff _88311_ (\oc8051_gm_cxrom_1.cell3.data [0], _01588_, clk);
  dff _88312_ (\oc8051_gm_cxrom_1.cell3.data [1], _01591_, clk);
  dff _88313_ (\oc8051_gm_cxrom_1.cell3.data [2], _01595_, clk);
  dff _88314_ (\oc8051_gm_cxrom_1.cell3.data [3], _01599_, clk);
  dff _88315_ (\oc8051_gm_cxrom_1.cell3.data [4], _01603_, clk);
  dff _88316_ (\oc8051_gm_cxrom_1.cell3.data [5], _01607_, clk);
  dff _88317_ (\oc8051_gm_cxrom_1.cell3.data [6], _01611_, clk);
  dff _88318_ (\oc8051_gm_cxrom_1.cell3.data [7], _01581_, clk);
  dff _88319_ (\oc8051_gm_cxrom_1.cell3.valid , _01584_, clk);
  dff _88320_ (\oc8051_gm_cxrom_1.cell4.data [0], _01630_, clk);
  dff _88321_ (\oc8051_gm_cxrom_1.cell4.data [1], _01631_, clk);
  dff _88322_ (\oc8051_gm_cxrom_1.cell4.data [2], _01634_, clk);
  dff _88323_ (\oc8051_gm_cxrom_1.cell4.data [3], _01638_, clk);
  dff _88324_ (\oc8051_gm_cxrom_1.cell4.data [4], _01642_, clk);
  dff _88325_ (\oc8051_gm_cxrom_1.cell4.data [5], _01646_, clk);
  dff _88326_ (\oc8051_gm_cxrom_1.cell4.data [6], _01650_, clk);
  dff _88327_ (\oc8051_gm_cxrom_1.cell4.data [7], _01628_, clk);
  dff _88328_ (\oc8051_gm_cxrom_1.cell4.valid , _01629_, clk);
  dff _88329_ (\oc8051_gm_cxrom_1.cell5.data [0], _01679_, clk);
  dff _88330_ (\oc8051_gm_cxrom_1.cell5.data [1], _01683_, clk);
  dff _88331_ (\oc8051_gm_cxrom_1.cell5.data [2], _01687_, clk);
  dff _88332_ (\oc8051_gm_cxrom_1.cell5.data [3], _01691_, clk);
  dff _88333_ (\oc8051_gm_cxrom_1.cell5.data [4], _01695_, clk);
  dff _88334_ (\oc8051_gm_cxrom_1.cell5.data [5], _01699_, clk);
  dff _88335_ (\oc8051_gm_cxrom_1.cell5.data [6], _01703_, clk);
  dff _88336_ (\oc8051_gm_cxrom_1.cell5.data [7], _01672_, clk);
  dff _88337_ (\oc8051_gm_cxrom_1.cell5.valid , _01675_, clk);
  dff _88338_ (\oc8051_gm_cxrom_1.cell6.data [0], _01732_, clk);
  dff _88339_ (\oc8051_gm_cxrom_1.cell6.data [1], _01736_, clk);
  dff _88340_ (\oc8051_gm_cxrom_1.cell6.data [2], _01740_, clk);
  dff _88341_ (\oc8051_gm_cxrom_1.cell6.data [3], _01743_, clk);
  dff _88342_ (\oc8051_gm_cxrom_1.cell6.data [4], _01747_, clk);
  dff _88343_ (\oc8051_gm_cxrom_1.cell6.data [5], _01751_, clk);
  dff _88344_ (\oc8051_gm_cxrom_1.cell6.data [6], _01755_, clk);
  dff _88345_ (\oc8051_gm_cxrom_1.cell6.data [7], _01725_, clk);
  dff _88346_ (\oc8051_gm_cxrom_1.cell6.valid , _01728_, clk);
  dff _88347_ (\oc8051_gm_cxrom_1.cell7.data [0], _01783_, clk);
  dff _88348_ (\oc8051_gm_cxrom_1.cell7.data [1], _01787_, clk);
  dff _88349_ (\oc8051_gm_cxrom_1.cell7.data [2], _01791_, clk);
  dff _88350_ (\oc8051_gm_cxrom_1.cell7.data [3], _01795_, clk);
  dff _88351_ (\oc8051_gm_cxrom_1.cell7.data [4], _01799_, clk);
  dff _88352_ (\oc8051_gm_cxrom_1.cell7.data [5], _01803_, clk);
  dff _88353_ (\oc8051_gm_cxrom_1.cell7.data [6], _01807_, clk);
  dff _88354_ (\oc8051_gm_cxrom_1.cell7.data [7], _01777_, clk);
  dff _88355_ (\oc8051_gm_cxrom_1.cell7.valid , _01779_, clk);
  dff _88356_ (\oc8051_gm_cxrom_1.cell8.data [0], _01835_, clk);
  dff _88357_ (\oc8051_gm_cxrom_1.cell8.data [1], _01839_, clk);
  dff _88358_ (\oc8051_gm_cxrom_1.cell8.data [2], _01843_, clk);
  dff _88359_ (\oc8051_gm_cxrom_1.cell8.data [3], _01847_, clk);
  dff _88360_ (\oc8051_gm_cxrom_1.cell8.data [4], _01851_, clk);
  dff _88361_ (\oc8051_gm_cxrom_1.cell8.data [5], _01854_, clk);
  dff _88362_ (\oc8051_gm_cxrom_1.cell8.data [6], _01858_, clk);
  dff _88363_ (\oc8051_gm_cxrom_1.cell8.data [7], _01828_, clk);
  dff _88364_ (\oc8051_gm_cxrom_1.cell8.valid , _01831_, clk);
  dff _88365_ (\oc8051_gm_cxrom_1.cell9.data [0], _01887_, clk);
  dff _88366_ (\oc8051_gm_cxrom_1.cell9.data [1], _01891_, clk);
  dff _88367_ (\oc8051_gm_cxrom_1.cell9.data [2], _01895_, clk);
  dff _88368_ (\oc8051_gm_cxrom_1.cell9.data [3], _01899_, clk);
  dff _88369_ (\oc8051_gm_cxrom_1.cell9.data [4], _01903_, clk);
  dff _88370_ (\oc8051_gm_cxrom_1.cell9.data [5], _01907_, clk);
  dff _88371_ (\oc8051_gm_cxrom_1.cell9.data [6], _01910_, clk);
  dff _88372_ (\oc8051_gm_cxrom_1.cell9.data [7], _01880_, clk);
  dff _88373_ (\oc8051_gm_cxrom_1.cell9.valid , _01883_, clk);
  dff _88374_ (\oc8051_golden_model_1.IRAM[15] [0], _40819_, clk);
  dff _88375_ (\oc8051_golden_model_1.IRAM[15] [1], _40821_, clk);
  dff _88376_ (\oc8051_golden_model_1.IRAM[15] [2], _40822_, clk);
  dff _88377_ (\oc8051_golden_model_1.IRAM[15] [3], _40823_, clk);
  dff _88378_ (\oc8051_golden_model_1.IRAM[15] [4], _40824_, clk);
  dff _88379_ (\oc8051_golden_model_1.IRAM[15] [5], _40825_, clk);
  dff _88380_ (\oc8051_golden_model_1.IRAM[15] [6], _40827_, clk);
  dff _88381_ (\oc8051_golden_model_1.IRAM[15] [7], _40565_, clk);
  dff _88382_ (\oc8051_golden_model_1.IRAM[14] [0], _40807_, clk);
  dff _88383_ (\oc8051_golden_model_1.IRAM[14] [1], _40809_, clk);
  dff _88384_ (\oc8051_golden_model_1.IRAM[14] [2], _40810_, clk);
  dff _88385_ (\oc8051_golden_model_1.IRAM[14] [3], _40811_, clk);
  dff _88386_ (\oc8051_golden_model_1.IRAM[14] [4], _40812_, clk);
  dff _88387_ (\oc8051_golden_model_1.IRAM[14] [5], _40813_, clk);
  dff _88388_ (\oc8051_golden_model_1.IRAM[14] [6], _40815_, clk);
  dff _88389_ (\oc8051_golden_model_1.IRAM[14] [7], _40816_, clk);
  dff _88390_ (\oc8051_golden_model_1.IRAM[13] [0], _40795_, clk);
  dff _88391_ (\oc8051_golden_model_1.IRAM[13] [1], _40796_, clk);
  dff _88392_ (\oc8051_golden_model_1.IRAM[13] [2], _40798_, clk);
  dff _88393_ (\oc8051_golden_model_1.IRAM[13] [3], _40799_, clk);
  dff _88394_ (\oc8051_golden_model_1.IRAM[13] [4], _40800_, clk);
  dff _88395_ (\oc8051_golden_model_1.IRAM[13] [5], _40801_, clk);
  dff _88396_ (\oc8051_golden_model_1.IRAM[13] [6], _40802_, clk);
  dff _88397_ (\oc8051_golden_model_1.IRAM[13] [7], _40804_, clk);
  dff _88398_ (\oc8051_golden_model_1.IRAM[12] [0], _40783_, clk);
  dff _88399_ (\oc8051_golden_model_1.IRAM[12] [1], _40784_, clk);
  dff _88400_ (\oc8051_golden_model_1.IRAM[12] [2], _40786_, clk);
  dff _88401_ (\oc8051_golden_model_1.IRAM[12] [3], _40787_, clk);
  dff _88402_ (\oc8051_golden_model_1.IRAM[12] [4], _40788_, clk);
  dff _88403_ (\oc8051_golden_model_1.IRAM[12] [5], _40789_, clk);
  dff _88404_ (\oc8051_golden_model_1.IRAM[12] [6], _40790_, clk);
  dff _88405_ (\oc8051_golden_model_1.IRAM[12] [7], _40792_, clk);
  dff _88406_ (\oc8051_golden_model_1.IRAM[11] [0], _40771_, clk);
  dff _88407_ (\oc8051_golden_model_1.IRAM[11] [1], _40772_, clk);
  dff _88408_ (\oc8051_golden_model_1.IRAM[11] [2], _40773_, clk);
  dff _88409_ (\oc8051_golden_model_1.IRAM[11] [3], _40774_, clk);
  dff _88410_ (\oc8051_golden_model_1.IRAM[11] [4], _40776_, clk);
  dff _88411_ (\oc8051_golden_model_1.IRAM[11] [5], _40777_, clk);
  dff _88412_ (\oc8051_golden_model_1.IRAM[11] [6], _40778_, clk);
  dff _88413_ (\oc8051_golden_model_1.IRAM[11] [7], _40779_, clk);
  dff _88414_ (\oc8051_golden_model_1.IRAM[10] [0], _40759_, clk);
  dff _88415_ (\oc8051_golden_model_1.IRAM[10] [1], _40760_, clk);
  dff _88416_ (\oc8051_golden_model_1.IRAM[10] [2], _40761_, clk);
  dff _88417_ (\oc8051_golden_model_1.IRAM[10] [3], _40762_, clk);
  dff _88418_ (\oc8051_golden_model_1.IRAM[10] [4], _40764_, clk);
  dff _88419_ (\oc8051_golden_model_1.IRAM[10] [5], _40765_, clk);
  dff _88420_ (\oc8051_golden_model_1.IRAM[10] [6], _40766_, clk);
  dff _88421_ (\oc8051_golden_model_1.IRAM[10] [7], _40767_, clk);
  dff _88422_ (\oc8051_golden_model_1.IRAM[9] [0], _40747_, clk);
  dff _88423_ (\oc8051_golden_model_1.IRAM[9] [1], _40748_, clk);
  dff _88424_ (\oc8051_golden_model_1.IRAM[9] [2], _40749_, clk);
  dff _88425_ (\oc8051_golden_model_1.IRAM[9] [3], _40750_, clk);
  dff _88426_ (\oc8051_golden_model_1.IRAM[9] [4], _40751_, clk);
  dff _88427_ (\oc8051_golden_model_1.IRAM[9] [5], _40753_, clk);
  dff _88428_ (\oc8051_golden_model_1.IRAM[9] [6], _40754_, clk);
  dff _88429_ (\oc8051_golden_model_1.IRAM[9] [7], _40755_, clk);
  dff _88430_ (\oc8051_golden_model_1.IRAM[8] [0], _40735_, clk);
  dff _88431_ (\oc8051_golden_model_1.IRAM[8] [1], _40736_, clk);
  dff _88432_ (\oc8051_golden_model_1.IRAM[8] [2], _40737_, clk);
  dff _88433_ (\oc8051_golden_model_1.IRAM[8] [3], _40738_, clk);
  dff _88434_ (\oc8051_golden_model_1.IRAM[8] [4], _40739_, clk);
  dff _88435_ (\oc8051_golden_model_1.IRAM[8] [5], _40741_, clk);
  dff _88436_ (\oc8051_golden_model_1.IRAM[8] [6], _40742_, clk);
  dff _88437_ (\oc8051_golden_model_1.IRAM[8] [7], _40743_, clk);
  dff _88438_ (\oc8051_golden_model_1.IRAM[7] [0], _40722_, clk);
  dff _88439_ (\oc8051_golden_model_1.IRAM[7] [1], _40723_, clk);
  dff _88440_ (\oc8051_golden_model_1.IRAM[7] [2], _40724_, clk);
  dff _88441_ (\oc8051_golden_model_1.IRAM[7] [3], _40725_, clk);
  dff _88442_ (\oc8051_golden_model_1.IRAM[7] [4], _40727_, clk);
  dff _88443_ (\oc8051_golden_model_1.IRAM[7] [5], _40728_, clk);
  dff _88444_ (\oc8051_golden_model_1.IRAM[7] [6], _40729_, clk);
  dff _88445_ (\oc8051_golden_model_1.IRAM[7] [7], _40730_, clk);
  dff _88446_ (\oc8051_golden_model_1.IRAM[6] [0], _40710_, clk);
  dff _88447_ (\oc8051_golden_model_1.IRAM[6] [1], _40711_, clk);
  dff _88448_ (\oc8051_golden_model_1.IRAM[6] [2], _40712_, clk);
  dff _88449_ (\oc8051_golden_model_1.IRAM[6] [3], _40713_, clk);
  dff _88450_ (\oc8051_golden_model_1.IRAM[6] [4], _40715_, clk);
  dff _88451_ (\oc8051_golden_model_1.IRAM[6] [5], _40716_, clk);
  dff _88452_ (\oc8051_golden_model_1.IRAM[6] [6], _40717_, clk);
  dff _88453_ (\oc8051_golden_model_1.IRAM[6] [7], _40718_, clk);
  dff _88454_ (\oc8051_golden_model_1.IRAM[5] [0], _40698_, clk);
  dff _88455_ (\oc8051_golden_model_1.IRAM[5] [1], _40699_, clk);
  dff _88456_ (\oc8051_golden_model_1.IRAM[5] [2], _40700_, clk);
  dff _88457_ (\oc8051_golden_model_1.IRAM[5] [3], _40701_, clk);
  dff _88458_ (\oc8051_golden_model_1.IRAM[5] [4], _40702_, clk);
  dff _88459_ (\oc8051_golden_model_1.IRAM[5] [5], _40704_, clk);
  dff _88460_ (\oc8051_golden_model_1.IRAM[5] [6], _40705_, clk);
  dff _88461_ (\oc8051_golden_model_1.IRAM[5] [7], _40706_, clk);
  dff _88462_ (\oc8051_golden_model_1.IRAM[4] [0], _40686_, clk);
  dff _88463_ (\oc8051_golden_model_1.IRAM[4] [1], _40687_, clk);
  dff _88464_ (\oc8051_golden_model_1.IRAM[4] [2], _40688_, clk);
  dff _88465_ (\oc8051_golden_model_1.IRAM[4] [3], _40689_, clk);
  dff _88466_ (\oc8051_golden_model_1.IRAM[4] [4], _40690_, clk);
  dff _88467_ (\oc8051_golden_model_1.IRAM[4] [5], _40692_, clk);
  dff _88468_ (\oc8051_golden_model_1.IRAM[4] [6], _40693_, clk);
  dff _88469_ (\oc8051_golden_model_1.IRAM[4] [7], _40694_, clk);
  dff _88470_ (\oc8051_golden_model_1.IRAM[3] [0], _40673_, clk);
  dff _88471_ (\oc8051_golden_model_1.IRAM[3] [1], _40674_, clk);
  dff _88472_ (\oc8051_golden_model_1.IRAM[3] [2], _40675_, clk);
  dff _88473_ (\oc8051_golden_model_1.IRAM[3] [3], _40676_, clk);
  dff _88474_ (\oc8051_golden_model_1.IRAM[3] [4], _40678_, clk);
  dff _88475_ (\oc8051_golden_model_1.IRAM[3] [5], _40679_, clk);
  dff _88476_ (\oc8051_golden_model_1.IRAM[3] [6], _40680_, clk);
  dff _88477_ (\oc8051_golden_model_1.IRAM[3] [7], _40681_, clk);
  dff _88478_ (\oc8051_golden_model_1.IRAM[2] [0], _40661_, clk);
  dff _88479_ (\oc8051_golden_model_1.IRAM[2] [1], _40662_, clk);
  dff _88480_ (\oc8051_golden_model_1.IRAM[2] [2], _40663_, clk);
  dff _88481_ (\oc8051_golden_model_1.IRAM[2] [3], _40664_, clk);
  dff _88482_ (\oc8051_golden_model_1.IRAM[2] [4], _40665_, clk);
  dff _88483_ (\oc8051_golden_model_1.IRAM[2] [5], _40667_, clk);
  dff _88484_ (\oc8051_golden_model_1.IRAM[2] [6], _40668_, clk);
  dff _88485_ (\oc8051_golden_model_1.IRAM[2] [7], _40669_, clk);
  dff _88486_ (\oc8051_golden_model_1.IRAM[1] [0], _40648_, clk);
  dff _88487_ (\oc8051_golden_model_1.IRAM[1] [1], _40649_, clk);
  dff _88488_ (\oc8051_golden_model_1.IRAM[1] [2], _40650_, clk);
  dff _88489_ (\oc8051_golden_model_1.IRAM[1] [3], _40651_, clk);
  dff _88490_ (\oc8051_golden_model_1.IRAM[1] [4], _40653_, clk);
  dff _88491_ (\oc8051_golden_model_1.IRAM[1] [5], _40654_, clk);
  dff _88492_ (\oc8051_golden_model_1.IRAM[1] [6], _40655_, clk);
  dff _88493_ (\oc8051_golden_model_1.IRAM[1] [7], _40656_, clk);
  dff _88494_ (\oc8051_golden_model_1.IRAM[0] [0], _40634_, clk);
  dff _88495_ (\oc8051_golden_model_1.IRAM[0] [1], _40635_, clk);
  dff _88496_ (\oc8051_golden_model_1.IRAM[0] [2], _40637_, clk);
  dff _88497_ (\oc8051_golden_model_1.IRAM[0] [3], _40638_, clk);
  dff _88498_ (\oc8051_golden_model_1.IRAM[0] [4], _40640_, clk);
  dff _88499_ (\oc8051_golden_model_1.IRAM[0] [5], _40641_, clk);
  dff _88500_ (\oc8051_golden_model_1.IRAM[0] [6], _40642_, clk);
  dff _88501_ (\oc8051_golden_model_1.IRAM[0] [7], _40644_, clk);
  dff _88502_ (\oc8051_golden_model_1.B [0], _43480_, clk);
  dff _88503_ (\oc8051_golden_model_1.B [1], _43481_, clk);
  dff _88504_ (\oc8051_golden_model_1.B [2], _43482_, clk);
  dff _88505_ (\oc8051_golden_model_1.B [3], _43485_, clk);
  dff _88506_ (\oc8051_golden_model_1.B [4], _43486_, clk);
  dff _88507_ (\oc8051_golden_model_1.B [5], _43487_, clk);
  dff _88508_ (\oc8051_golden_model_1.B [6], _43488_, clk);
  dff _88509_ (\oc8051_golden_model_1.B [7], _40566_, clk);
  dff _88510_ (\oc8051_golden_model_1.ACC [0], _43491_, clk);
  dff _88511_ (\oc8051_golden_model_1.ACC [1], _43492_, clk);
  dff _88512_ (\oc8051_golden_model_1.ACC [2], _43493_, clk);
  dff _88513_ (\oc8051_golden_model_1.ACC [3], _43494_, clk);
  dff _88514_ (\oc8051_golden_model_1.ACC [4], _43495_, clk);
  dff _88515_ (\oc8051_golden_model_1.ACC [5], _43496_, clk);
  dff _88516_ (\oc8051_golden_model_1.ACC [6], _43497_, clk);
  dff _88517_ (\oc8051_golden_model_1.ACC [7], _40567_, clk);
  dff _88518_ (\oc8051_golden_model_1.DPL [0], _43498_, clk);
  dff _88519_ (\oc8051_golden_model_1.DPL [1], _43499_, clk);
  dff _88520_ (\oc8051_golden_model_1.DPL [2], _43500_, clk);
  dff _88521_ (\oc8051_golden_model_1.DPL [3], _43501_, clk);
  dff _88522_ (\oc8051_golden_model_1.DPL [4], _43502_, clk);
  dff _88523_ (\oc8051_golden_model_1.DPL [5], _43505_, clk);
  dff _88524_ (\oc8051_golden_model_1.DPL [6], _43506_, clk);
  dff _88525_ (\oc8051_golden_model_1.DPL [7], _40568_, clk);
  dff _88526_ (\oc8051_golden_model_1.DPH [0], _43507_, clk);
  dff _88527_ (\oc8051_golden_model_1.DPH [1], _43510_, clk);
  dff _88528_ (\oc8051_golden_model_1.DPH [2], _43511_, clk);
  dff _88529_ (\oc8051_golden_model_1.DPH [3], _43512_, clk);
  dff _88530_ (\oc8051_golden_model_1.DPH [4], _43513_, clk);
  dff _88531_ (\oc8051_golden_model_1.DPH [5], _43514_, clk);
  dff _88532_ (\oc8051_golden_model_1.DPH [6], _43515_, clk);
  dff _88533_ (\oc8051_golden_model_1.DPH [7], _40569_, clk);
  dff _88534_ (\oc8051_golden_model_1.IE [0], _43516_, clk);
  dff _88535_ (\oc8051_golden_model_1.IE [1], _43517_, clk);
  dff _88536_ (\oc8051_golden_model_1.IE [2], _43518_, clk);
  dff _88537_ (\oc8051_golden_model_1.IE [3], _43519_, clk);
  dff _88538_ (\oc8051_golden_model_1.IE [4], _43520_, clk);
  dff _88539_ (\oc8051_golden_model_1.IE [5], _43521_, clk);
  dff _88540_ (\oc8051_golden_model_1.IE [6], _43522_, clk);
  dff _88541_ (\oc8051_golden_model_1.IE [7], _40571_, clk);
  dff _88542_ (\oc8051_golden_model_1.IP [0], _43525_, clk);
  dff _88543_ (\oc8051_golden_model_1.IP [1], _43526_, clk);
  dff _88544_ (\oc8051_golden_model_1.IP [2], _43527_, clk);
  dff _88545_ (\oc8051_golden_model_1.IP [3], _43530_, clk);
  dff _88546_ (\oc8051_golden_model_1.IP [4], _43531_, clk);
  dff _88547_ (\oc8051_golden_model_1.IP [5], _43532_, clk);
  dff _88548_ (\oc8051_golden_model_1.IP [6], _43533_, clk);
  dff _88549_ (\oc8051_golden_model_1.IP [7], _40572_, clk);
  dff _88550_ (\oc8051_golden_model_1.P0 [0], _43534_, clk);
  dff _88551_ (\oc8051_golden_model_1.P0 [1], _43535_, clk);
  dff _88552_ (\oc8051_golden_model_1.P0 [2], _43536_, clk);
  dff _88553_ (\oc8051_golden_model_1.P0 [3], _43537_, clk);
  dff _88554_ (\oc8051_golden_model_1.P0 [4], _43538_, clk);
  dff _88555_ (\oc8051_golden_model_1.P0 [5], _43539_, clk);
  dff _88556_ (\oc8051_golden_model_1.P0 [6], _43540_, clk);
  dff _88557_ (\oc8051_golden_model_1.P0 [7], _40573_, clk);
  dff _88558_ (\oc8051_golden_model_1.P1 [0], _43543_, clk);
  dff _88559_ (\oc8051_golden_model_1.P1 [1], _43544_, clk);
  dff _88560_ (\oc8051_golden_model_1.P1 [2], _43545_, clk);
  dff _88561_ (\oc8051_golden_model_1.P1 [3], _43546_, clk);
  dff _88562_ (\oc8051_golden_model_1.P1 [4], _43547_, clk);
  dff _88563_ (\oc8051_golden_model_1.P1 [5], _43550_, clk);
  dff _88564_ (\oc8051_golden_model_1.P1 [6], _43551_, clk);
  dff _88565_ (\oc8051_golden_model_1.P1 [7], _40574_, clk);
  dff _88566_ (\oc8051_golden_model_1.P2 [0], _43552_, clk);
  dff _88567_ (\oc8051_golden_model_1.P2 [1], _43553_, clk);
  dff _88568_ (\oc8051_golden_model_1.P2 [2], _43554_, clk);
  dff _88569_ (\oc8051_golden_model_1.P2 [3], _43555_, clk);
  dff _88570_ (\oc8051_golden_model_1.P2 [4], _43556_, clk);
  dff _88571_ (\oc8051_golden_model_1.P2 [5], _43557_, clk);
  dff _88572_ (\oc8051_golden_model_1.P2 [6], _43558_, clk);
  dff _88573_ (\oc8051_golden_model_1.P2 [7], _40575_, clk);
  dff _88574_ (\oc8051_golden_model_1.P3 [0], _43561_, clk);
  dff _88575_ (\oc8051_golden_model_1.P3 [1], _43562_, clk);
  dff _88576_ (\oc8051_golden_model_1.P3 [2], _43563_, clk);
  dff _88577_ (\oc8051_golden_model_1.P3 [3], _43564_, clk);
  dff _88578_ (\oc8051_golden_model_1.P3 [4], _43565_, clk);
  dff _88579_ (\oc8051_golden_model_1.P3 [5], _43566_, clk);
  dff _88580_ (\oc8051_golden_model_1.P3 [6], _43567_, clk);
  dff _88581_ (\oc8051_golden_model_1.P3 [7], _40577_, clk);
  dff _88582_ (\oc8051_golden_model_1.PSW [0], _43570_, clk);
  dff _88583_ (\oc8051_golden_model_1.PSW [1], _43571_, clk);
  dff _88584_ (\oc8051_golden_model_1.PSW [2], _43572_, clk);
  dff _88585_ (\oc8051_golden_model_1.PSW [3], _43573_, clk);
  dff _88586_ (\oc8051_golden_model_1.PSW [4], _43574_, clk);
  dff _88587_ (\oc8051_golden_model_1.PSW [5], _43575_, clk);
  dff _88588_ (\oc8051_golden_model_1.PSW [6], _43576_, clk);
  dff _88589_ (\oc8051_golden_model_1.PSW [7], _40578_, clk);
  dff _88590_ (\oc8051_golden_model_1.PCON [0], _43579_, clk);
  dff _88591_ (\oc8051_golden_model_1.PCON [1], _43580_, clk);
  dff _88592_ (\oc8051_golden_model_1.PCON [2], _43581_, clk);
  dff _88593_ (\oc8051_golden_model_1.PCON [3], _43582_, clk);
  dff _88594_ (\oc8051_golden_model_1.PCON [4], _43583_, clk);
  dff _88595_ (\oc8051_golden_model_1.PCON [5], _43584_, clk);
  dff _88596_ (\oc8051_golden_model_1.PCON [6], _43585_, clk);
  dff _88597_ (\oc8051_golden_model_1.PCON [7], _40579_, clk);
  dff _88598_ (\oc8051_golden_model_1.SBUF [0], _43588_, clk);
  dff _88599_ (\oc8051_golden_model_1.SBUF [1], _43589_, clk);
  dff _88600_ (\oc8051_golden_model_1.SBUF [2], _43590_, clk);
  dff _88601_ (\oc8051_golden_model_1.SBUF [3], _43591_, clk);
  dff _88602_ (\oc8051_golden_model_1.SBUF [4], _43592_, clk);
  dff _88603_ (\oc8051_golden_model_1.SBUF [5], _43594_, clk);
  dff _88604_ (\oc8051_golden_model_1.SBUF [6], _43595_, clk);
  dff _88605_ (\oc8051_golden_model_1.SBUF [7], _40580_, clk);
  dff _88606_ (\oc8051_golden_model_1.SCON [0], _43596_, clk);
  dff _88607_ (\oc8051_golden_model_1.SCON [1], _43599_, clk);
  dff _88608_ (\oc8051_golden_model_1.SCON [2], _43600_, clk);
  dff _88609_ (\oc8051_golden_model_1.SCON [3], _43601_, clk);
  dff _88610_ (\oc8051_golden_model_1.SCON [4], _43602_, clk);
  dff _88611_ (\oc8051_golden_model_1.SCON [5], _43603_, clk);
  dff _88612_ (\oc8051_golden_model_1.SCON [6], _43604_, clk);
  dff _88613_ (\oc8051_golden_model_1.SCON [7], _40581_, clk);
  dff _88614_ (\oc8051_golden_model_1.SP [0], _43606_, clk);
  dff _88615_ (\oc8051_golden_model_1.SP [1], _43607_, clk);
  dff _88616_ (\oc8051_golden_model_1.SP [2], _43608_, clk);
  dff _88617_ (\oc8051_golden_model_1.SP [3], _43609_, clk);
  dff _88618_ (\oc8051_golden_model_1.SP [4], _43610_, clk);
  dff _88619_ (\oc8051_golden_model_1.SP [5], _43611_, clk);
  dff _88620_ (\oc8051_golden_model_1.SP [6], _43612_, clk);
  dff _88621_ (\oc8051_golden_model_1.SP [7], _40583_, clk);
  dff _88622_ (\oc8051_golden_model_1.TCON [0], _43613_, clk);
  dff _88623_ (\oc8051_golden_model_1.TCON [1], _43614_, clk);
  dff _88624_ (\oc8051_golden_model_1.TCON [2], _43615_, clk);
  dff _88625_ (\oc8051_golden_model_1.TCON [3], _43618_, clk);
  dff _88626_ (\oc8051_golden_model_1.TCON [4], _43619_, clk);
  dff _88627_ (\oc8051_golden_model_1.TCON [5], _43620_, clk);
  dff _88628_ (\oc8051_golden_model_1.TCON [6], _43621_, clk);
  dff _88629_ (\oc8051_golden_model_1.TCON [7], _40584_, clk);
  dff _88630_ (\oc8051_golden_model_1.TH0 [0], _43624_, clk);
  dff _88631_ (\oc8051_golden_model_1.TH0 [1], _43625_, clk);
  dff _88632_ (\oc8051_golden_model_1.TH0 [2], _43626_, clk);
  dff _88633_ (\oc8051_golden_model_1.TH0 [3], _43627_, clk);
  dff _88634_ (\oc8051_golden_model_1.TH0 [4], _43628_, clk);
  dff _88635_ (\oc8051_golden_model_1.TH0 [5], _43629_, clk);
  dff _88636_ (\oc8051_golden_model_1.TH0 [6], _43630_, clk);
  dff _88637_ (\oc8051_golden_model_1.TH0 [7], _40585_, clk);
  dff _88638_ (\oc8051_golden_model_1.TH1 [0], _43631_, clk);
  dff _88639_ (\oc8051_golden_model_1.TH1 [1], _43632_, clk);
  dff _88640_ (\oc8051_golden_model_1.TH1 [2], _43633_, clk);
  dff _88641_ (\oc8051_golden_model_1.TH1 [3], _43634_, clk);
  dff _88642_ (\oc8051_golden_model_1.TH1 [4], _43635_, clk);
  dff _88643_ (\oc8051_golden_model_1.TH1 [5], _43638_, clk);
  dff _88644_ (\oc8051_golden_model_1.TH1 [6], _43639_, clk);
  dff _88645_ (\oc8051_golden_model_1.TH1 [7], _40586_, clk);
  dff _88646_ (\oc8051_golden_model_1.TL0 [0], _43640_, clk);
  dff _88647_ (\oc8051_golden_model_1.TL0 [1], _43643_, clk);
  dff _88648_ (\oc8051_golden_model_1.TL0 [2], _43644_, clk);
  dff _88649_ (\oc8051_golden_model_1.TL0 [3], _43645_, clk);
  dff _88650_ (\oc8051_golden_model_1.TL0 [4], _43646_, clk);
  dff _88651_ (\oc8051_golden_model_1.TL0 [5], _43647_, clk);
  dff _88652_ (\oc8051_golden_model_1.TL0 [6], _43648_, clk);
  dff _88653_ (\oc8051_golden_model_1.TL0 [7], _40587_, clk);
  dff _88654_ (\oc8051_golden_model_1.TL1 [0], _43649_, clk);
  dff _88655_ (\oc8051_golden_model_1.TL1 [1], _43650_, clk);
  dff _88656_ (\oc8051_golden_model_1.TL1 [2], _43651_, clk);
  dff _88657_ (\oc8051_golden_model_1.TL1 [3], _43652_, clk);
  dff _88658_ (\oc8051_golden_model_1.TL1 [4], _43653_, clk);
  dff _88659_ (\oc8051_golden_model_1.TL1 [5], _43654_, clk);
  dff _88660_ (\oc8051_golden_model_1.TL1 [6], _43655_, clk);
  dff _88661_ (\oc8051_golden_model_1.TL1 [7], _40589_, clk);
  dff _88662_ (\oc8051_golden_model_1.TMOD [0], _43658_, clk);
  dff _88663_ (\oc8051_golden_model_1.TMOD [1], _43659_, clk);
  dff _88664_ (\oc8051_golden_model_1.TMOD [2], _43660_, clk);
  dff _88665_ (\oc8051_golden_model_1.TMOD [3], _43663_, clk);
  dff _88666_ (\oc8051_golden_model_1.TMOD [4], _43664_, clk);
  dff _88667_ (\oc8051_golden_model_1.TMOD [5], _43665_, clk);
  dff _88668_ (\oc8051_golden_model_1.TMOD [6], _43666_, clk);
  dff _88669_ (\oc8051_golden_model_1.TMOD [7], _40590_, clk);
  dff _88670_ (\oc8051_golden_model_1.PC [0], _43667_, clk);
  dff _88671_ (\oc8051_golden_model_1.PC [1], _43670_, clk);
  dff _88672_ (\oc8051_golden_model_1.PC [2], _43671_, clk);
  dff _88673_ (\oc8051_golden_model_1.PC [3], _43672_, clk);
  dff _88674_ (\oc8051_golden_model_1.PC [4], _43673_, clk);
  dff _88675_ (\oc8051_golden_model_1.PC [5], _43674_, clk);
  dff _88676_ (\oc8051_golden_model_1.PC [6], _43675_, clk);
  dff _88677_ (\oc8051_golden_model_1.PC [7], _43676_, clk);
  dff _88678_ (\oc8051_golden_model_1.PC [8], _43677_, clk);
  dff _88679_ (\oc8051_golden_model_1.PC [9], _43678_, clk);
  dff _88680_ (\oc8051_golden_model_1.PC [10], _43679_, clk);
  dff _88681_ (\oc8051_golden_model_1.PC [11], _43682_, clk);
  dff _88682_ (\oc8051_golden_model_1.PC [12], _43683_, clk);
  dff _88683_ (\oc8051_golden_model_1.PC [13], _43684_, clk);
  dff _88684_ (\oc8051_golden_model_1.PC [14], _43685_, clk);
  dff _88685_ (\oc8051_golden_model_1.PC [15], _40591_, clk);
  dff _88686_ (\oc8051_golden_model_1.P0INREG [0], _43686_, clk);
  dff _88687_ (\oc8051_golden_model_1.P0INREG [1], _43687_, clk);
  dff _88688_ (\oc8051_golden_model_1.P0INREG [2], _43688_, clk);
  dff _88689_ (\oc8051_golden_model_1.P0INREG [3], _43689_, clk);
  dff _88690_ (\oc8051_golden_model_1.P0INREG [4], _43690_, clk);
  dff _88691_ (\oc8051_golden_model_1.P0INREG [5], _43691_, clk);
  dff _88692_ (\oc8051_golden_model_1.P0INREG [6], _43692_, clk);
  dff _88693_ (\oc8051_golden_model_1.P0INREG [7], _40592_, clk);
  dff _88694_ (\oc8051_golden_model_1.P1INREG [0], _43695_, clk);
  dff _88695_ (\oc8051_golden_model_1.P1INREG [1], _43696_, clk);
  dff _88696_ (\oc8051_golden_model_1.P1INREG [2], _43697_, clk);
  dff _88697_ (\oc8051_golden_model_1.P1INREG [3], _43698_, clk);
  dff _88698_ (\oc8051_golden_model_1.P1INREG [4], _43699_, clk);
  dff _88699_ (\oc8051_golden_model_1.P1INREG [5], _43702_, clk);
  dff _88700_ (\oc8051_golden_model_1.P1INREG [6], _43703_, clk);
  dff _88701_ (\oc8051_golden_model_1.P1INREG [7], _40593_, clk);
  dff _88702_ (\oc8051_golden_model_1.P2INREG [0], _43704_, clk);
  dff _88703_ (\oc8051_golden_model_1.P2INREG [1], _43705_, clk);
  dff _88704_ (\oc8051_golden_model_1.P2INREG [2], _43706_, clk);
  dff _88705_ (\oc8051_golden_model_1.P2INREG [3], _43707_, clk);
  dff _88706_ (\oc8051_golden_model_1.P2INREG [4], _43708_, clk);
  dff _88707_ (\oc8051_golden_model_1.P2INREG [5], _43709_, clk);
  dff _88708_ (\oc8051_golden_model_1.P2INREG [6], _43710_, clk);
  dff _88709_ (\oc8051_golden_model_1.P2INREG [7], _40595_, clk);
  dff _88710_ (\oc8051_golden_model_1.P3INREG [0], _43713_, clk);
  dff _88711_ (\oc8051_golden_model_1.P3INREG [1], _43714_, clk);
  dff _88712_ (\oc8051_golden_model_1.P3INREG [2], _43715_, clk);
  dff _88713_ (\oc8051_golden_model_1.P3INREG [3], _43716_, clk);
  dff _88714_ (\oc8051_golden_model_1.P3INREG [4], _43717_, clk);
  dff _88715_ (\oc8051_golden_model_1.P3INREG [5], _43718_, clk);
  dff _88716_ (\oc8051_golden_model_1.P3INREG [6], _43719_, clk);
  dff _88717_ (\oc8051_golden_model_1.P3INREG [7], _40596_, clk);
  dff _88718_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03014_, clk);
  dff _88719_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03025_, clk);
  dff _88720_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03046_, clk);
  dff _88721_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03068_, clk);
  dff _88722_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03089_, clk);
  dff _88723_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00893_, clk);
  dff _88724_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03100_, clk);
  dff _88725_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00862_, clk);
  dff _88726_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03111_, clk);
  dff _88727_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03122_, clk);
  dff _88728_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03133_, clk);
  dff _88729_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03144_, clk);
  dff _88730_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03155_, clk);
  dff _88731_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03166_, clk);
  dff _88732_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03177_, clk);
  dff _88733_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00914_, clk);
  dff _88734_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02465_, clk);
  dff _88735_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22434_, clk);
  dff _88736_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02660_, clk);
  dff _88737_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02854_, clk);
  dff _88738_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03057_, clk);
  dff _88739_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03268_, clk);
  dff _88740_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03469_, clk);
  dff _88741_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03670_, clk);
  dff _88742_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03871_, clk);
  dff _88743_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04072_, clk);
  dff _88744_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04173_, clk);
  dff _88745_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04274_, clk);
  dff _88746_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04375_, clk);
  dff _88747_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04476_, clk);
  dff _88748_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04577_, clk);
  dff _88749_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04678_, clk);
  dff _88750_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04779_, clk);
  dff _88751_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24620_, clk);
  dff _88752_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38825_, clk);
  dff _88753_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38826_, clk);
  dff _88754_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38827_, clk);
  dff _88755_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38828_, clk);
  dff _88756_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38829_, clk);
  dff _88757_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38830_, clk);
  dff _88758_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38831_, clk);
  dff _88759_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38811_, clk);
  dff _88760_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38832_, clk);
  dff _88761_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38834_, clk);
  dff _88762_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38835_, clk);
  dff _88763_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38836_, clk);
  dff _88764_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38837_, clk);
  dff _88765_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38838_, clk);
  dff _88766_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38840_, clk);
  dff _88767_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38813_, clk);
  dff _88768_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38841_, clk);
  dff _88769_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38842_, clk);
  dff _88770_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38843_, clk);
  dff _88771_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38844_, clk);
  dff _88772_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38846_, clk);
  dff _88773_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38847_, clk);
  dff _88774_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38848_, clk);
  dff _88775_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38814_, clk);
  dff _88776_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _30468_, clk);
  dff _88777_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06011_, clk);
  dff _88778_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _30471_, clk);
  dff _88779_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _06014_, clk);
  dff _88780_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _30473_, clk);
  dff _88781_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _30475_, clk);
  dff _88782_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _06017_, clk);
  dff _88783_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _30477_, clk);
  dff _88784_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _30479_, clk);
  dff _88785_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06020_, clk);
  dff _88786_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _30481_, clk);
  dff _88787_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _06023_, clk);
  dff _88788_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _30483_, clk);
  dff _88789_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _30485_, clk);
  dff _88790_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _30487_, clk);
  dff _88791_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _06026_, clk);
  dff _88792_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _30489_, clk);
  dff _88793_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _06029_, clk);
  dff _88794_ (\oc8051_top_1.oc8051_decoder1.wr , _06032_, clk);
  dff _88795_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _06091_, clk);
  dff _88796_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _06093_, clk);
  dff _88797_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _05996_, clk);
  dff _88798_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _06096_, clk);
  dff _88799_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _06099_, clk);
  dff _88800_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05999_, clk);
  dff _88801_ (\oc8051_top_1.oc8051_decoder1.state [0], _06102_, clk);
  dff _88802_ (\oc8051_top_1.oc8051_decoder1.state [1], _06002_, clk);
  dff _88803_ (\oc8051_top_1.oc8051_decoder1.op [0], _06105_, clk);
  dff _88804_ (\oc8051_top_1.oc8051_decoder1.op [1], _06108_, clk);
  dff _88805_ (\oc8051_top_1.oc8051_decoder1.op [2], _06111_, clk);
  dff _88806_ (\oc8051_top_1.oc8051_decoder1.op [3], _06114_, clk);
  dff _88807_ (\oc8051_top_1.oc8051_decoder1.op [4], _06117_, clk);
  dff _88808_ (\oc8051_top_1.oc8051_decoder1.op [5], _06120_, clk);
  dff _88809_ (\oc8051_top_1.oc8051_decoder1.op [6], _06123_, clk);
  dff _88810_ (\oc8051_top_1.oc8051_decoder1.op [7], _06005_, clk);
  dff _88811_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _06008_, clk);
  dff _88812_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39617_, clk);
  dff _88813_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38985_, clk);
  dff _88814_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38986_, clk);
  dff _88815_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38987_, clk);
  dff _88816_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38989_, clk);
  dff _88817_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38990_, clk);
  dff _88818_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38991_, clk);
  dff _88819_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38992_, clk);
  dff _88820_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38993_, clk);
  dff _88821_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38994_, clk);
  dff _88822_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38995_, clk);
  dff _88823_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38996_, clk);
  dff _88824_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38997_, clk);
  dff _88825_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38998_, clk);
  dff _88826_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39000_, clk);
  dff _88827_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39001_, clk);
  dff _88828_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38872_, clk);
  dff _88829_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39005_, clk);
  dff _88830_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39006_, clk);
  dff _88831_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39007_, clk);
  dff _88832_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39008_, clk);
  dff _88833_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39009_, clk);
  dff _88834_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39010_, clk);
  dff _88835_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39011_, clk);
  dff _88836_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39012_, clk);
  dff _88837_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39013_, clk);
  dff _88838_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39014_, clk);
  dff _88839_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39015_, clk);
  dff _88840_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39016_, clk);
  dff _88841_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39017_, clk);
  dff _88842_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39018_, clk);
  dff _88843_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39019_, clk);
  dff _88844_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38874_, clk);
  dff _88845_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39197_, clk);
  dff _88846_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39198_, clk);
  dff _88847_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39199_, clk);
  dff _88848_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39200_, clk);
  dff _88849_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39201_, clk);
  dff _88850_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39202_, clk);
  dff _88851_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39204_, clk);
  dff _88852_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39205_, clk);
  dff _88853_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39206_, clk);
  dff _88854_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39207_, clk);
  dff _88855_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39208_, clk);
  dff _88856_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39209_, clk);
  dff _88857_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39210_, clk);
  dff _88858_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39211_, clk);
  dff _88859_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39212_, clk);
  dff _88860_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39213_, clk);
  dff _88861_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39215_, clk);
  dff _88862_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39216_, clk);
  dff _88863_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39217_, clk);
  dff _88864_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39218_, clk);
  dff _88865_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39219_, clk);
  dff _88866_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39220_, clk);
  dff _88867_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39221_, clk);
  dff _88868_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39222_, clk);
  dff _88869_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39223_, clk);
  dff _88870_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39224_, clk);
  dff _88871_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39226_, clk);
  dff _88872_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39227_, clk);
  dff _88873_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39228_, clk);
  dff _88874_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39229_, clk);
  dff _88875_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39230_, clk);
  dff _88876_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38938_, clk);
  dff _88877_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38911_, clk);
  dff _88878_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _88879_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39231_, clk);
  dff _88880_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39232_, clk);
  dff _88881_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39233_, clk);
  dff _88882_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39234_, clk);
  dff _88883_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38913_, clk);
  dff _88884_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39236_, clk);
  dff _88885_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39237_, clk);
  dff _88886_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39238_, clk);
  dff _88887_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39239_, clk);
  dff _88888_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39240_, clk);
  dff _88889_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39242_, clk);
  dff _88890_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39243_, clk);
  dff _88891_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38914_, clk);
  dff _88892_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39244_, clk);
  dff _88893_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39245_, clk);
  dff _88894_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39246_, clk);
  dff _88895_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39247_, clk);
  dff _88896_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39248_, clk);
  dff _88897_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39249_, clk);
  dff _88898_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39250_, clk);
  dff _88899_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38916_, clk);
  dff _88900_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39252_, clk);
  dff _88901_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39253_, clk);
  dff _88902_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39254_, clk);
  dff _88903_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39255_, clk);
  dff _88904_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39256_, clk);
  dff _88905_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39257_, clk);
  dff _88906_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39258_, clk);
  dff _88907_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38917_, clk);
  dff _88908_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38918_, clk);
  dff _88909_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38919_, clk);
  dff _88910_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39259_, clk);
  dff _88911_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39260_, clk);
  dff _88912_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39261_, clk);
  dff _88913_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39263_, clk);
  dff _88914_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39264_, clk);
  dff _88915_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39265_, clk);
  dff _88916_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39266_, clk);
  dff _88917_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38920_, clk);
  dff _88918_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39267_, clk);
  dff _88919_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39268_, clk);
  dff _88920_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39269_, clk);
  dff _88921_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39270_, clk);
  dff _88922_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39271_, clk);
  dff _88923_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39272_, clk);
  dff _88924_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39274_, clk);
  dff _88925_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39275_, clk);
  dff _88926_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39276_, clk);
  dff _88927_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39277_, clk);
  dff _88928_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39278_, clk);
  dff _88929_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39279_, clk);
  dff _88930_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39280_, clk);
  dff _88931_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39281_, clk);
  dff _88932_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39282_, clk);
  dff _88933_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38922_, clk);
  dff _88934_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39283_, clk);
  dff _88935_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39285_, clk);
  dff _88936_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39286_, clk);
  dff _88937_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39287_, clk);
  dff _88938_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39288_, clk);
  dff _88939_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39289_, clk);
  dff _88940_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39290_, clk);
  dff _88941_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39291_, clk);
  dff _88942_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39292_, clk);
  dff _88943_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39293_, clk);
  dff _88944_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39294_, clk);
  dff _88945_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39296_, clk);
  dff _88946_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39297_, clk);
  dff _88947_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39298_, clk);
  dff _88948_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39299_, clk);
  dff _88949_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38923_, clk);
  dff _88950_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38924_, clk);
  dff _88951_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38927_, clk);
  dff _88952_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38925_, clk);
  dff _88953_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39300_, clk);
  dff _88954_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39301_, clk);
  dff _88955_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39302_, clk);
  dff _88956_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39303_, clk);
  dff _88957_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39304_, clk);
  dff _88958_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39305_, clk);
  dff _88959_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39307_, clk);
  dff _88960_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38928_, clk);
  dff _88961_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39308_, clk);
  dff _88962_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39309_, clk);
  dff _88963_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38929_, clk);
  dff _88964_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39310_, clk);
  dff _88965_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39311_, clk);
  dff _88966_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39312_, clk);
  dff _88967_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39313_, clk);
  dff _88968_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39314_, clk);
  dff _88969_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39315_, clk);
  dff _88970_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39316_, clk);
  dff _88971_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38930_, clk);
  dff _88972_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39317_, clk);
  dff _88973_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39318_, clk);
  dff _88974_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39319_, clk);
  dff _88975_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39320_, clk);
  dff _88976_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39321_, clk);
  dff _88977_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39322_, clk);
  dff _88978_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39323_, clk);
  dff _88979_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38931_, clk);
  dff _88980_ (\oc8051_top_1.oc8051_memory_interface1.reti , _38932_, clk);
  dff _88981_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39324_, clk);
  dff _88982_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39325_, clk);
  dff _88983_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39326_, clk);
  dff _88984_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39328_, clk);
  dff _88985_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39329_, clk);
  dff _88986_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39330_, clk);
  dff _88987_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39331_, clk);
  dff _88988_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38934_, clk);
  dff _88989_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _38935_, clk);
  dff _88990_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38936_, clk);
  dff _88991_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39332_, clk);
  dff _88992_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39333_, clk);
  dff _88993_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39334_, clk);
  dff _88994_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38937_, clk);
  dff _88995_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39335_, clk);
  dff _88996_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39336_, clk);
  dff _88997_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39337_, clk);
  dff _88998_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39339_, clk);
  dff _88999_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39340_, clk);
  dff _89000_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39341_, clk);
  dff _89001_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39342_, clk);
  dff _89002_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39343_, clk);
  dff _89003_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39344_, clk);
  dff _89004_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39345_, clk);
  dff _89005_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39346_, clk);
  dff _89006_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39347_, clk);
  dff _89007_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39348_, clk);
  dff _89008_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39350_, clk);
  dff _89009_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39351_, clk);
  dff _89010_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39352_, clk);
  dff _89011_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39353_, clk);
  dff _89012_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39354_, clk);
  dff _89013_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39355_, clk);
  dff _89014_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39356_, clk);
  dff _89015_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39357_, clk);
  dff _89016_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39358_, clk);
  dff _89017_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39359_, clk);
  dff _89018_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39361_, clk);
  dff _89019_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39362_, clk);
  dff _89020_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39363_, clk);
  dff _89021_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39364_, clk);
  dff _89022_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39365_, clk);
  dff _89023_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39366_, clk);
  dff _89024_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39367_, clk);
  dff _89025_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39368_, clk);
  dff _89026_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38939_, clk);
  dff _89027_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39369_, clk);
  dff _89028_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39370_, clk);
  dff _89029_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39372_, clk);
  dff _89030_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39373_, clk);
  dff _89031_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39374_, clk);
  dff _89032_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39375_, clk);
  dff _89033_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39376_, clk);
  dff _89034_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38940_, clk);
  dff _89035_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38941_, clk);
  dff _89036_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38942_, clk);
  dff _89037_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39377_, clk);
  dff _89038_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39378_, clk);
  dff _89039_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39379_, clk);
  dff _89040_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39380_, clk);
  dff _89041_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39381_, clk);
  dff _89042_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39383_, clk);
  dff _89043_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39384_, clk);
  dff _89044_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39385_, clk);
  dff _89045_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39386_, clk);
  dff _89046_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39387_, clk);
  dff _89047_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39388_, clk);
  dff _89048_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39389_, clk);
  dff _89049_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39390_, clk);
  dff _89050_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39391_, clk);
  dff _89051_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39392_, clk);
  dff _89052_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38943_, clk);
  dff _89053_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38944_, clk);
  dff _89054_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38945_, clk);
  dff _89055_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38946_, clk);
  dff _89056_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39394_, clk);
  dff _89057_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39395_, clk);
  dff _89058_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39396_, clk);
  dff _89059_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39397_, clk);
  dff _89060_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39398_, clk);
  dff _89061_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39399_, clk);
  dff _89062_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39400_, clk);
  dff _89063_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39401_, clk);
  dff _89064_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39402_, clk);
  dff _89065_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39403_, clk);
  dff _89066_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39405_, clk);
  dff _89067_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39406_, clk);
  dff _89068_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39407_, clk);
  dff _89069_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39408_, clk);
  dff _89070_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39409_, clk);
  dff _89071_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38947_, clk);
  dff _89072_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38948_, clk);
  dff _89073_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39764_, clk);
  dff _89074_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39783_, clk);
  dff _89075_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39784_, clk);
  dff _89076_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39785_, clk);
  dff _89077_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39786_, clk);
  dff _89078_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39787_, clk);
  dff _89079_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39788_, clk);
  dff _89080_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39789_, clk);
  dff _89081_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39765_, clk);
  dff _89082_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39766_, clk);
  dff _89083_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39790_, clk);
  dff _89084_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39791_, clk);
  dff _89085_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39767_, clk);
  dff _89086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _43133_, clk);
  dff _89087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _43139_, clk);
  dff _89088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _43145_, clk);
  dff _89089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _43151_, clk);
  dff _89090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _43157_, clk);
  dff _89091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _43163_, clk);
  dff _89092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _43169_, clk);
  dff _89093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _43172_, clk);
  dff _89094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _43413_, clk);
  dff _89095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _43417_, clk);
  dff _89096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _43421_, clk);
  dff _89097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _43425_, clk);
  dff _89098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _43429_, clk);
  dff _89099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _43433_, clk);
  dff _89100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _43437_, clk);
  dff _89101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _43440_, clk);
  dff _89102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _43180_, clk);
  dff _89103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _43184_, clk);
  dff _89104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _43188_, clk);
  dff _89105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _43192_, clk);
  dff _89106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _43196_, clk);
  dff _89107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _43200_, clk);
  dff _89108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _43204_, clk);
  dff _89109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _43207_, clk);
  dff _89110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _43378_, clk);
  dff _89111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _43382_, clk);
  dff _89112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _43386_, clk);
  dff _89113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _43390_, clk);
  dff _89114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _43394_, clk);
  dff _89115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _43398_, clk);
  dff _89116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _43402_, clk);
  dff _89117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _43405_, clk);
  dff _89118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _43346_, clk);
  dff _89119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _43350_, clk);
  dff _89120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _43354_, clk);
  dff _89121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _43358_, clk);
  dff _89122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _43362_, clk);
  dff _89123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _43366_, clk);
  dff _89124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _43370_, clk);
  dff _89125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _43373_, clk);
  dff _89126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _43315_, clk);
  dff _89127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _43319_, clk);
  dff _89128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _43322_, clk);
  dff _89129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _43326_, clk);
  dff _89130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _43330_, clk);
  dff _89131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _43334_, clk);
  dff _89132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _43338_, clk);
  dff _89133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _43341_, clk);
  dff _89134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _43283_, clk);
  dff _89135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _43287_, clk);
  dff _89136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _43291_, clk);
  dff _89137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _43295_, clk);
  dff _89138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _43299_, clk);
  dff _89139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _43303_, clk);
  dff _89140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _43307_, clk);
  dff _89141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _43310_, clk);
  dff _89142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _43248_, clk);
  dff _89143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _43252_, clk);
  dff _89144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _43256_, clk);
  dff _89145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _43260_, clk);
  dff _89146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _43264_, clk);
  dff _89147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _43268_, clk);
  dff _89148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _43272_, clk);
  dff _89149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _43275_, clk);
  dff _89150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _43215_, clk);
  dff _89151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _43219_, clk);
  dff _89152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _43223_, clk);
  dff _89153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _43227_, clk);
  dff _89154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _43231_, clk);
  dff _89155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _43235_, clk);
  dff _89156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _43239_, clk);
  dff _89157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _43242_, clk);
  dff _89158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _43445_, clk);
  dff _89159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _43449_, clk);
  dff _89160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _43453_, clk);
  dff _89161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _43457_, clk);
  dff _89162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _43461_, clk);
  dff _89163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _43465_, clk);
  dff _89164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _43469_, clk);
  dff _89165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _43472_, clk);
  dff _89166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _43796_, clk);
  dff _89167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _43800_, clk);
  dff _89168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _43804_, clk);
  dff _89169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _43808_, clk);
  dff _89170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _43812_, clk);
  dff _89171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _43816_, clk);
  dff _89172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _43820_, clk);
  dff _89173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _43823_, clk);
  dff _89174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _43764_, clk);
  dff _89175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _43768_, clk);
  dff _89176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _43772_, clk);
  dff _89177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _43776_, clk);
  dff _89178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _43780_, clk);
  dff _89179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _43784_, clk);
  dff _89180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _43788_, clk);
  dff _89181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _43791_, clk);
  dff _89182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _43732_, clk);
  dff _89183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _43736_, clk);
  dff _89184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _43740_, clk);
  dff _89185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _43744_, clk);
  dff _89186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _43748_, clk);
  dff _89187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _43752_, clk);
  dff _89188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _43756_, clk);
  dff _89189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _43759_, clk);
  dff _89190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _43617_, clk);
  dff _89191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _43637_, clk);
  dff _89192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _43657_, clk);
  dff _89193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _43669_, clk);
  dff _89194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _43694_, clk);
  dff _89195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _43712_, clk);
  dff _89196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _43723_, clk);
  dff _89197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _43726_, clk);
  dff _89198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _43477_, clk);
  dff _89199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _43484_, clk);
  dff _89200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _43504_, clk);
  dff _89201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _43524_, clk);
  dff _89202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _43542_, clk);
  dff _89203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _43560_, clk);
  dff _89204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _43578_, clk);
  dff _89205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _43593_, clk);
  dff _89206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _43826_, clk);
  dff _89207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _43829_, clk);
  dff _89208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _43833_, clk);
  dff _89209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _43837_, clk);
  dff _89210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _43841_, clk);
  dff _89211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _43844_, clk);
  dff _89212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _43847_, clk);
  dff _89213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _42875_, clk);
  dff _89214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _01406_, clk);
  dff _89215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _01408_, clk);
  dff _89216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _01410_, clk);
  dff _89217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _01412_, clk);
  dff _89218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _01414_, clk);
  dff _89219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _01416_, clk);
  dff _89220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _01418_, clk);
  dff _89221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _42863_, clk);
  dff _89222_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _89223_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _89224_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _89225_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _89226_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _89227_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _89228_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _89229_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _89230_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _89231_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _89232_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _89233_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _89234_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _89235_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _89236_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _89237_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _89238_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _89239_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _89240_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _89241_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _89242_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _89243_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _89244_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _89245_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _89246_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _89247_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _89248_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _89249_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _89250_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _89251_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _89252_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _89253_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _89254_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _89255_ (\oc8051_top_1.oc8051_sfr1.bit_out , _39648_, clk);
  dff _89256_ (\oc8051_top_1.oc8051_sfr1.wait_data , _39649_, clk);
  dff _89257_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39713_, clk);
  dff _89258_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39714_, clk);
  dff _89259_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39715_, clk);
  dff _89260_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39716_, clk);
  dff _89261_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39717_, clk);
  dff _89262_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39718_, clk);
  dff _89263_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39719_, clk);
  dff _89264_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39650_, clk);
  dff _89265_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39651_, clk);
  dff _89266_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24174_, clk);
  dff _89267_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24186_, clk);
  dff _89268_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24198_, clk);
  dff _89269_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24210_, clk);
  dff _89270_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24222_, clk);
  dff _89271_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24234_, clk);
  dff _89272_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24246_, clk);
  dff _89273_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22313_, clk);
  dff _89274_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08932_, clk);
  dff _89275_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08943_, clk);
  dff _89276_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08954_, clk);
  dff _89277_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08965_, clk);
  dff _89278_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08976_, clk);
  dff _89279_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08987_, clk);
  dff _89280_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08998_, clk);
  dff _89281_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06695_, clk);
  dff _89282_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13612_, clk);
  dff _89283_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13621_, clk);
  dff _89284_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13631_, clk);
  dff _89285_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13640_, clk);
  dff _89286_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13650_, clk);
  dff _89287_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13660_, clk);
  dff _89288_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13670_, clk);
  dff _89289_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12702_, clk);
  dff _89290_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13679_, clk);
  dff _89291_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13688_, clk);
  dff _89292_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13698_, clk);
  dff _89293_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13708_, clk);
  dff _89294_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13718_, clk);
  dff _89295_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13727_, clk);
  dff _89296_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13736_, clk);
  dff _89297_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12723_, clk);
  dff _89298_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0, clk);
  dff _89299_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0, clk);
  dff _89300_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _89301_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _41806_, clk);
  dff _89302_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _42729_, clk);
  dff _89303_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _42731_, clk);
  dff _89304_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42733_, clk);
  dff _89305_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _42734_, clk);
  dff _89306_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _42736_, clk);
  dff _89307_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42738_, clk);
  dff _89308_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42740_, clk);
  dff _89309_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41804_, clk);
  dff _89310_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _42742_, clk);
  dff _89311_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _41802_, clk);
  dff _89312_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _41800_, clk);
  dff _89313_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _42744_, clk);
  dff _89314_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _42746_, clk);
  dff _89315_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _41798_, clk);
  dff _89316_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _42748_, clk);
  dff _89317_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _42750_, clk);
  dff _89318_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _41796_, clk);
  dff _89319_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _42752_, clk);
  dff _89320_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41795_, clk);
  dff _89321_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _42754_, clk);
  dff _89322_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41793_, clk);
  dff _89323_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _41761_, clk);
  dff _89324_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _41759_, clk);
  dff _89325_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _41757_, clk);
  dff _89326_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _41755_, clk);
  dff _89327_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _42756_, clk);
  dff _89328_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _42758_, clk);
  dff _89329_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _42760_, clk);
  dff _89330_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _41753_, clk);
  dff _89331_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _42762_, clk);
  dff _89332_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _42764_, clk);
  dff _89333_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _42766_, clk);
  dff _89334_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _42768_, clk);
  dff _89335_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _42770_, clk);
  dff _89336_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _42772_, clk);
  dff _89337_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _42774_, clk);
  dff _89338_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41751_, clk);
  dff _89339_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _42776_, clk);
  dff _89340_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _42778_, clk);
  dff _89341_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _42780_, clk);
  dff _89342_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _42782_, clk);
  dff _89343_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _42784_, clk);
  dff _89344_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _42786_, clk);
  dff _89345_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _42788_, clk);
  dff _89346_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _41748_, clk);
  dff _89347_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41207_, clk);
  dff _89348_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41209_, clk);
  dff _89349_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41211_, clk);
  dff _89350_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41213_, clk);
  dff _89351_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41214_, clk);
  dff _89352_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41216_, clk);
  dff _89353_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41218_, clk);
  dff _89354_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35484_, clk);
  dff _89355_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41220_, clk);
  dff _89356_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41221_, clk);
  dff _89357_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41223_, clk);
  dff _89358_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41225_, clk);
  dff _89359_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41227_, clk);
  dff _89360_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41228_, clk);
  dff _89361_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41230_, clk);
  dff _89362_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35507_, clk);
  dff _89363_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41232_, clk);
  dff _89364_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41234_, clk);
  dff _89365_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41235_, clk);
  dff _89366_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41237_, clk);
  dff _89367_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41239_, clk);
  dff _89368_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41240_, clk);
  dff _89369_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41242_, clk);
  dff _89370_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35530_, clk);
  dff _89371_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41244_, clk);
  dff _89372_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41245_, clk);
  dff _89373_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41247_, clk);
  dff _89374_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41249_, clk);
  dff _89375_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41251_, clk);
  dff _89376_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41252_, clk);
  dff _89377_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41254_, clk);
  dff _89378_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35552_, clk);
  dff _89379_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21479_, clk);
  dff _89380_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21490_, clk);
  dff _89381_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21502_, clk);
  dff _89382_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21514_, clk);
  dff _89383_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21526_, clk);
  dff _89384_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21538_, clk);
  dff _89385_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16545_, clk);
  dff _89386_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09544_, clk);
  dff _89387_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10690_, clk);
  dff _89388_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10701_, clk);
  dff _89389_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10712_, clk);
  dff _89390_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10723_, clk);
  dff _89391_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10734_, clk);
  dff _89392_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10745_, clk);
  dff _89393_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10756_, clk);
  dff _89394_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09564_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0988 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0988 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0988 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0988 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0988 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0988 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0988 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0989 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0990 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0991 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0992 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0993 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0995 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0996 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1011 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1011 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1011 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1011 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1011 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1011 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1011 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1018 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1019 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.n1027 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1027 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1027 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1027 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1027 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1043 , \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.n1044 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1044 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1044 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1044 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1044 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1044 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1044 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1137 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1137 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1137 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1137 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1139 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1141 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1141 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1142 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1142 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1143 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1144 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1144 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1145 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1145 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1146 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1194 , \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n1239 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1240 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1240 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1240 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1240 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1240 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1240 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1240 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1241 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1241 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1241 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1241 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1241 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1241 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1241 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1242 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1242 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1242 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1242 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1242 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1242 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1242 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1242 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1243 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1244 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1244 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1244 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1247 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1247 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1247 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1247 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1247 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1248 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1248 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1248 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1248 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1248 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1248 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1248 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1249 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1251 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1252 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1253 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1254 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1255 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1264 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1280 , \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.n1281 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1281 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1281 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1281 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1281 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1281 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1281 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1323 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1323 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1323 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1323 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1323 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1323 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1323 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1323 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1323 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1323 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1323 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1323 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1323 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1323 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1323 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1323 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1325 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1325 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1325 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1325 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1325 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1325 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1325 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1327 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1328 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1329 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1330 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1331 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1332 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1340 , \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.n1341 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1341 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1341 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1341 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1341 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1341 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1343 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1347 [8], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1349 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1349 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1349 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1349 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1350 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1354 [4], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1356 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1356 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1356 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1356 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1356 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1356 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1356 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1356 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1356 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1364 , \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1365 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1365 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1365 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1365 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1365 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1365 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1366 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1366 [6], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1381 , \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.n1382 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1382 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1382 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1382 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1404 [8], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1405 , \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1410 [4], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1411 , \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1419 , \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1420 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1420 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1420 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1420 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1420 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1420 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1421 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1421 [1], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1421 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1421 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1421 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1421 [5], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1421 [6], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1436 , \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.n1437 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1437 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1437 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1437 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1439 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1439 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1439 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1439 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1439 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1439 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1439 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1439 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1439 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1441 [8], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1442 , \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1443 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1443 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1443 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1443 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1444 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1444 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1444 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1446 [4], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1447 , \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1448 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1448 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1448 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1448 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1448 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1448 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1448 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1448 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1448 [8], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1455 , \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1456 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1456 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1456 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1456 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1456 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1456 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1457 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1457 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1457 [6], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1472 , \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1473 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1473 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1473 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1473 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1476 [8], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1477 , \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1484 , \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1485 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1485 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1485 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1485 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1485 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1485 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1486 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1486 [1], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1486 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1486 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1486 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1486 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1486 [6], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1489 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1489 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1489 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1489 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1489 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1489 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1489 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1489 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1489 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1491 [8], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1493 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1495 [4], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1496 , \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1497 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1497 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1497 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1497 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1497 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1497 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1497 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1497 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1497 [8], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1521 , \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1522 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1524 [4], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1525 , \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1527 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1527 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1527 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1527 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1527 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1527 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1527 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1528 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1528 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1530 [8], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1531 , \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1538 , \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1539 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1539 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1539 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1539 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1539 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1539 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1540 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1540 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1540 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1540 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1540 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1540 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1540 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1541 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1541 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1541 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1541 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1541 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1541 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1541 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1543 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1543 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1543 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1543 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1543 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1543 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1543 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1544 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1544 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1544 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1547 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1547 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1548 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1548 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1548 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1549 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1549 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1549 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1549 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1549 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1549 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1549 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1549 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1550 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1550 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1550 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1550 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1550 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1550 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1550 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1550 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1551 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1552 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1553 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1555 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1557 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1559 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1566 , \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1571 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [8], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1575 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1575 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [4], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1585 , \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1586 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1586 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1586 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1586 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1586 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1586 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1587 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1602 , \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.n1603 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1603 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1603 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1603 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [8], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1608 , \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1610 [4], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1611 , \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1618 , \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1619 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1619 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1619 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1619 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1619 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1619 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1620 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1620 [1], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1620 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1620 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1620 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1620 [5], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1620 [6], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1635 , \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.n1636 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1636 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1636 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1636 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [8], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1641 , \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1643 [4], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1644 , \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1651 , \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1652 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1652 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1652 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1652 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1652 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1652 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1653 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1653 [1], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1653 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1653 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1653 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1653 [5], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1653 [6], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1668 , \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.n1669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [8], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1674 , \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1676 [4], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1677 , \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1684 , \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1685 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1685 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1685 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1685 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1685 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1685 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1686 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1686 [1], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1686 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1686 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1686 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1686 [5], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1686 [6], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1701 , \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.n1702 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1702 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1702 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1702 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1727 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1727 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1727 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1727 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1727 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1727 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1727 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1728 [0], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1728 [1], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1728 [2], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1728 [3], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1728 [4], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1728 [5], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1728 [6], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1729 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1784 , \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.n1785 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1785 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1785 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1785 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1785 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1785 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1785 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1801 , \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.n1802 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1802 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1802 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1802 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1802 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1802 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1802 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1818 , \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.n1819 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1819 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1819 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1819 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1819 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1819 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1819 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1835 , \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.n1836 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1836 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1836 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1836 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1836 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1836 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1836 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1859 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1859 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1859 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1859 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1859 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1859 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1859 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1860 [0], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1860 [1], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1860 [2], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1860 [3], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1860 [4], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1860 [5], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1860 [6], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1861 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1916 , \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.n1917 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1917 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1917 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1917 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1917 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1917 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1917 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1933 , \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.n1934 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1934 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1934 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1934 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1934 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1934 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1934 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1950 , \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.n1951 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1951 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1951 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1951 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1951 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1951 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1951 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1967 , \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.n1968 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1968 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1968 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1968 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1968 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1968 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1968 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2065 , \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.n2066 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2066 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2066 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2066 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2066 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2066 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2066 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2082 , \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.n2083 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2083 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2083 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2083 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2083 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2083 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2083 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2099 , \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.n2100 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2100 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2100 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2100 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2100 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2100 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2116 , \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.n2117 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2117 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2117 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2117 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2117 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2117 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2117 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2121 , \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2122 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2122 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2122 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2122 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2122 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2122 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2122 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2123 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2123 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2123 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2123 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2123 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2123 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2124 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2124 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2124 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2124 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2124 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2124 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2124 [6], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2125 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2125 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2125 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2125 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2125 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2125 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2125 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2140 , \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.n2141 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2141 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2141 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2141 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2141 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2141 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2180 , \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2181 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2181 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2181 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2181 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2181 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2181 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2181 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2181 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2182 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2182 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2182 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2182 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2182 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2182 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2182 [6], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2183 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2183 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2183 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2183 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2183 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2183 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2183 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2190 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2190 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2190 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2190 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2191 , \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2192 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2192 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2192 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2192 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2192 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2192 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2193 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2193 [1], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2193 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2193 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2193 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2193 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2193 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2208 , \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.n2209 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2209 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2209 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2209 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2209 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2209 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2421 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2424 , \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2426 , \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2432 , \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2433 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2433 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2433 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2433 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2433 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2433 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2434 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2434 [1], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2434 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2434 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2434 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2434 [5], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2434 [6], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2449 , \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.n2450 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2450 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2450 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2450 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 , \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2456 , \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2462 , \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2463 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2463 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2463 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2463 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2463 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2463 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2464 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2464 [1], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2464 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2464 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2464 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2464 [5], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2464 [6], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2479 , \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.n2480 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2480 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2480 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2480 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 , \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2486 , \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2492 , \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2493 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2493 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2493 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2494 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2494 [1], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2494 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2494 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2494 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2494 [5], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2494 [6], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2509 , \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.n2510 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2510 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2510 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2510 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 , \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2516 , \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2522 , \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2523 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2523 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2523 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2523 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2523 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2523 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2524 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2524 [1], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2524 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2524 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2524 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2524 [5], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2524 [6], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2539 , \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.n2540 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2540 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2540 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2540 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2545 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2545 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2545 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2545 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2545 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2545 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2545 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2547 [6], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2548 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2548 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2548 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2552 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2552 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2552 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2552 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2552 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2552 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2552 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2552 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2552 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2558 , \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2559 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2559 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2559 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2560 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2575 , \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.n2576 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2576 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2576 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2576 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2576 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2576 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2579 , \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2581 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2581 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2581 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2581 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2581 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2581 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2581 [6], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2582 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2582 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2582 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2582 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2582 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2582 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2582 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2614 , \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2615 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2615 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2615 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2615 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2615 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2615 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2615 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2615 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2616 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2616 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2616 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2616 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2616 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2616 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2616 [6], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2617 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2617 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2617 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2617 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2617 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2617 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2617 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2622 , \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2623 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2623 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2623 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2623 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2624 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2624 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2624 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2624 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2624 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2624 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2624 [6], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2625 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2625 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2625 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2625 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2625 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2625 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2625 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2630 , \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2631 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2631 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2631 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2631 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2631 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2631 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2631 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2631 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2632 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2632 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2632 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2632 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2632 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2632 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2632 [6], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2633 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2633 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2633 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2633 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2633 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2633 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2633 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2638 , \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2639 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2639 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2639 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2640 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2640 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2640 [6], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2641 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2641 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2641 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2641 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2641 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2641 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2641 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2646 , \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2647 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2647 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2647 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2647 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2647 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2647 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2647 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2647 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2648 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2648 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2648 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2648 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2648 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2648 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2648 [6], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2649 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2649 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2649 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2649 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2649 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2649 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2649 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2674 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2674 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2674 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2674 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2674 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2674 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2675 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2675 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2675 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2675 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2675 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2675 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2675 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2676 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2676 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2676 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2676 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2676 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2676 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2676 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2676 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2677 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2677 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2677 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2677 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2678 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2678 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2678 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2678 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2678 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2678 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2679 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2680 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2681 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2682 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2683 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2684 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2685 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2686 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2693 , \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2715 [0], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2715 [1], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2715 [2], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2715 [3], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2715 [4], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2715 [5], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2715 [6], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2731 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2731 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2731 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2731 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2731 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2731 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2731 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2732 , \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2733 , \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2734 , \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2735 , \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2736 , \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2737 , \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2738 , \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2739 , \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2746 , \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.n2747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2747 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2747 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2747 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2762 , \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.n2763 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2763 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2763 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2763 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2763 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2763 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2763 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2795 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2795 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2795 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2795 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2795 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2795 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2795 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2795 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2796 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2796 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2796 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2796 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2796 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2796 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2796 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2797 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2797 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2797 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2797 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2797 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2797 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2797 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2797 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 , \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2818 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2818 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2818 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2818 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2818 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2818 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2818 [6], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2833 , \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.n2834 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2834 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2834 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2834 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2834 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2834 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2838 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2839 [0], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2839 [1], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2839 [2], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2839 [3], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2840 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2840 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2840 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2840 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2841 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2842 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2843 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2844 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2855 , \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.n2856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2874 , \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.n2875 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2875 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2875 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2875 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2875 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2875 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2875 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2891 , \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.n2892 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2892 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2892 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2892 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2892 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2892 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2892 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
