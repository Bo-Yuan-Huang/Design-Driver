
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire [15:0] _26822_;
  wire [7:0] _26823_;
  wire [7:0] _26824_;
  wire [7:0] _26825_;
  wire [7:0] _26826_;
  wire [7:0] _26827_;
  wire [7:0] _26828_;
  wire [7:0] _26829_;
  wire [7:0] _26830_;
  wire [7:0] _26831_;
  wire [7:0] _26832_;
  wire [7:0] _26833_;
  wire [7:0] _26834_;
  wire [7:0] _26835_;
  wire [7:0] _26836_;
  wire [7:0] _26837_;
  wire [7:0] _26838_;
  wire _26839_;
  wire [7:0] _26840_;
  wire [2:0] _26841_;
  wire [2:0] _26842_;
  wire [1:0] _26843_;
  wire [7:0] _26844_;
  wire _26845_;
  wire [1:0] _26846_;
  wire [1:0] _26847_;
  wire [2:0] _26848_;
  wire [2:0] _26849_;
  wire [1:0] _26850_;
  wire [3:0] _26851_;
  wire [1:0] _26852_;
  wire _26853_;
  wire [7:0] _26854_;
  wire [7:0] _26855_;
  wire [7:0] _26856_;
  wire [7:0] _26857_;
  wire [7:0] _26858_;
  wire [7:0] _26859_;
  wire [7:0] _26860_;
  wire [7:0] _26861_;
  wire [15:0] _26862_;
  wire [15:0] _26863_;
  wire _26864_;
  wire [4:0] _26865_;
  wire [7:0] _26866_;
  wire [7:0] _26867_;
  wire _26868_;
  wire _26869_;
  wire [15:0] _26870_;
  wire [15:0] _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire [7:0] _26875_;
  wire [2:0] _26876_;
  wire [7:0] _26877_;
  wire _26878_;
  wire [7:0] _26879_;
  wire _26880_;
  wire _26881_;
  wire [3:0] _26882_;
  wire [31:0] _26883_;
  wire [31:0] _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire [15:0] _26888_;
  wire _26889_;
  wire _26890_;
  wire [7:0] _26891_;
  wire _26892_;
  wire [2:0] _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire [7:0] _27313_;
  wire _27314_;
  wire [3:0] _27315_;
  wire _27316_;
  wire _27317_;
  wire [7:0] _27318_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _27319_ (_22731_, rst);
  not _27320_ (_22732_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor _27321_ (_22733_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _27322_ (_22734_, _22733_, _22732_);
  not _27323_ (_22735_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _27324_ (_22736_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and _27325_ (_22737_, _22736_, _22735_);
  and _27326_ (_22738_, _22737_, _22734_);
  and _27327_ (_22740_, _22738_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _27328_ (_22741_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _27329_ (_22742_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27330_ (_22744_, _22740_, _22742_);
  or _27331_ (_22745_, _22744_, _22741_);
  and _27332_ (_26863_[0], _22745_, _22731_);
  and _27333_ (_22746_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _27334_ (_22747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _27335_ (_22749_, _22740_, _22747_);
  or _27336_ (_22750_, _22749_, _22746_);
  and _27337_ (_26863_[1], _22750_, _22731_);
  and _27338_ (_22751_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _27339_ (_22752_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27340_ (_22753_, _22740_, _22752_);
  or _27341_ (_22755_, _22753_, _22751_);
  and _27342_ (_26863_[2], _22755_, _22731_);
  and _27343_ (_22757_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _27344_ (_22758_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27345_ (_22759_, _22740_, _22758_);
  or _27346_ (_22760_, _22759_, _22757_);
  and _27347_ (_26863_[3], _22760_, _22731_);
  or _27348_ (_22761_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not _27349_ (_22762_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand _27350_ (_22763_, _22740_, _22762_);
  and _27351_ (_22764_, _22763_, _22731_);
  and _27352_ (_26863_[4], _22764_, _22761_);
  or _27353_ (_22766_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not _27354_ (_22767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _27355_ (_22768_, _22740_, _22767_);
  and _27356_ (_22769_, _22768_, _22731_);
  and _27357_ (_26863_[5], _22769_, _22766_);
  or _27358_ (_22771_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not _27359_ (_22772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _27360_ (_22773_, _22740_, _22772_);
  and _27361_ (_22774_, _22773_, _22731_);
  and _27362_ (_26863_[6], _22774_, _22771_);
  and _27363_ (_22775_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _27364_ (_22776_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _27365_ (_22777_, _22740_, _22776_);
  or _27366_ (_22778_, _22777_, _22775_);
  and _27367_ (_26863_[7], _22778_, _22731_);
  or _27368_ (_22779_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not _27369_ (_22780_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _27370_ (_22781_, _22740_, _22780_);
  and _27371_ (_22782_, _22781_, _22731_);
  and _27372_ (_26863_[8], _22782_, _22779_);
  and _27373_ (_22783_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not _27374_ (_22784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _27375_ (_22785_, _22740_, _22784_);
  or _27376_ (_22786_, _22785_, _22783_);
  and _27377_ (_26863_[9], _22786_, _22731_);
  or _27378_ (_22788_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not _27379_ (_22789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _27380_ (_22790_, _22740_, _22789_);
  and _27381_ (_22791_, _22790_, _22731_);
  and _27382_ (_26863_[10], _22791_, _22788_);
  or _27383_ (_22792_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  not _27384_ (_22793_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _27385_ (_22794_, _22740_, _22793_);
  and _27386_ (_22795_, _22794_, _22731_);
  and _27387_ (_26863_[11], _22795_, _22792_);
  or _27388_ (_22796_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _27389_ (_22797_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _27390_ (_22799_, _22740_, _22797_);
  and _27391_ (_22800_, _22799_, _22731_);
  and _27392_ (_26863_[12], _22800_, _22796_);
  and _27393_ (_22801_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _27394_ (_22802_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _27395_ (_22803_, _22740_, _22802_);
  or _27396_ (_22804_, _22803_, _22801_);
  and _27397_ (_26863_[13], _22804_, _22731_);
  or _27398_ (_22805_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not _27399_ (_22806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _27400_ (_22808_, _22740_, _22806_);
  and _27401_ (_22809_, _22808_, _22731_);
  and _27402_ (_26863_[14], _22809_, _22805_);
  and _27403_ (_22810_, \oc8051_top_1.oc8051_decoder1.wr , _22735_);
  not _27404_ (_22811_, _22810_);
  not _27405_ (_22812_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _27406_ (_22813_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _22735_);
  and _27407_ (_22814_, _22813_, _22812_);
  and _27408_ (_22815_, _22814_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _27409_ (_22816_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _27410_ (_22817_, _22816_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _27411_ (_22818_, _22817_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _27412_ (_22820_, _22818_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _27413_ (_22821_, _22820_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _27414_ (_22822_, _22821_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _27415_ (_22823_, _22822_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _27416_ (_22824_, _22822_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _27417_ (_22825_, _22824_, _22823_);
  and _27418_ (_22826_, _22825_, _22815_);
  not _27419_ (_22827_, _22826_);
  and _27420_ (_22828_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _27421_ (_22829_, _22828_, _22813_);
  not _27422_ (_22830_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _27423_ (_22831_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _22735_);
  and _27424_ (_22832_, _22831_, _22830_);
  and _27425_ (_22833_, _22832_, _22812_);
  and _27426_ (_22834_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _27427_ (_22835_, _22834_, _22829_);
  nor _27428_ (_22836_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _27429_ (_22837_, _22836_, _22813_);
  and _27430_ (_22838_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _27431_ (_22839_, _22832_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _27432_ (_22840_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _27433_ (_22841_, _22840_, _22838_);
  and _27434_ (_22843_, _22841_, _22835_);
  nand _27435_ (_22844_, _22843_, _22827_);
  not _27436_ (_22845_, _22844_);
  nor _27437_ (_22846_, _22845_, _22814_);
  nor _27438_ (_22847_, _22846_, _22811_);
  not _27439_ (_22849_, _22847_);
  and _27440_ (_22850_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _27441_ (_22851_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _27442_ (_22852_, _22851_, _22850_);
  not _27443_ (_22853_, _22818_);
  not _27444_ (_22854_, _22815_);
  nor _27445_ (_22855_, _22817_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _27446_ (_22856_, _22855_, _22854_);
  and _27447_ (_22857_, _22856_, _22853_);
  and _27448_ (_22858_, _22836_, _22830_);
  nor _27449_ (_22859_, _22858_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _27450_ (_22861_, _22859_);
  and _27451_ (_22862_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _27452_ (_22863_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _27453_ (_22864_, _22863_, _22862_);
  not _27454_ (_22865_, _22864_);
  nor _27455_ (_22866_, _22865_, _22857_);
  and _27456_ (_22867_, _22866_, _22852_);
  not _27457_ (_22868_, _22867_);
  not _27458_ (_22869_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27459_ (_22871_, _22844_, _22869_);
  and _27460_ (_22872_, _22871_, _22868_);
  not _27461_ (_22874_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _27462_ (_22875_, _22815_, _22874_);
  and _27463_ (_22876_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _27464_ (_22877_, _22876_, _22875_);
  and _27465_ (_22878_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  not _27466_ (_22880_, _22878_);
  and _27467_ (_22881_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _27468_ (_22882_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _27469_ (_22884_, _22882_, _22881_);
  and _27470_ (_22885_, _22884_, _22880_);
  and _27471_ (_22886_, _22885_, _22877_);
  nor _27472_ (_22887_, _22886_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27473_ (_22888_, _22887_, _22872_);
  nor _27474_ (_22890_, _22888_, _22849_);
  nor _27475_ (_22891_, _22818_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _27476_ (_22893_, _22891_);
  nor _27477_ (_22894_, _22854_, _22820_);
  and _27478_ (_22896_, _22894_, _22893_);
  and _27479_ (_22897_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor _27480_ (_22898_, _22897_, _22896_);
  and _27481_ (_22899_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _27482_ (_22900_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _27483_ (_22901_, _22900_, _22899_);
  and _27484_ (_22902_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _27485_ (_22903_, _22902_, _22829_);
  and _27486_ (_22904_, _22903_, _22901_);
  and _27487_ (_22905_, _22904_, _22898_);
  not _27488_ (_22906_, _22905_);
  and _27489_ (_22907_, _22906_, _22871_);
  and _27490_ (_22908_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nor _27491_ (_22909_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _27492_ (_22910_, _22909_, _22816_);
  and _27493_ (_22911_, _22910_, _22815_);
  nor _27494_ (_22912_, _22911_, _22908_);
  and _27495_ (_22913_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and _27496_ (_22914_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _27497_ (_22916_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _27498_ (_22917_, _22916_, _22914_);
  nor _27499_ (_22918_, _22917_, _22913_);
  and _27500_ (_22919_, _22918_, _22912_);
  nor _27501_ (_22920_, _22919_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27502_ (_22921_, _22920_, _22907_);
  nor _27503_ (_22922_, _22921_, _22849_);
  nor _27504_ (_22923_, _22922_, _22890_);
  nor _27505_ (_22924_, _22820_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _27506_ (_22925_, _22924_);
  nor _27507_ (_22926_, _22854_, _22821_);
  and _27508_ (_22927_, _22926_, _22925_);
  not _27509_ (_22928_, _22927_);
  and _27510_ (_22930_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nor _27511_ (_22931_, _22930_, _22829_);
  and _27512_ (_22932_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _27513_ (_22933_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _27514_ (_22934_, _22933_, _22932_);
  and _27515_ (_22935_, _22934_, _22931_);
  and _27516_ (_22936_, _22935_, _22928_);
  not _27517_ (_22937_, _22936_);
  and _27518_ (_22938_, _22937_, _22871_);
  nor _27519_ (_22940_, _22816_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _27520_ (_22941_, _22940_, _22817_);
  and _27521_ (_22942_, _22941_, _22815_);
  and _27522_ (_22943_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _27523_ (_22945_, _22943_, _22942_);
  and _27524_ (_22946_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _27525_ (_22947_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _27526_ (_22948_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _27527_ (_22949_, _22948_, _22947_);
  nor _27528_ (_22950_, _22949_, _22946_);
  and _27529_ (_22951_, _22950_, _22945_);
  nor _27530_ (_22952_, _22951_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27531_ (_22953_, _22952_, _22938_);
  nor _27532_ (_22954_, _22953_, _22849_);
  nor _27533_ (_22956_, _22821_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _27534_ (_22957_, _22956_);
  nor _27535_ (_22958_, _22854_, _22822_);
  and _27536_ (_22960_, _22958_, _22957_);
  not _27537_ (_22961_, _22960_);
  and _27538_ (_22962_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  nor _27539_ (_22963_, _22962_, _22829_);
  and _27540_ (_22964_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and _27541_ (_22965_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _27542_ (_22966_, _22965_, _22964_);
  and _27543_ (_22967_, _22966_, _22963_);
  and _27544_ (_22968_, _22967_, _22961_);
  not _27545_ (_22969_, _22968_);
  and _27546_ (_22970_, _22969_, _22871_);
  nor _27547_ (_22971_, _22871_, _22867_);
  nor _27548_ (_22972_, _22971_, _22970_);
  and _27549_ (_22973_, _22972_, _22954_);
  and _27550_ (_22974_, _22973_, _22923_);
  nor _27551_ (_22975_, _22905_, _22871_);
  and _27552_ (_22976_, _22975_, _22847_);
  and _27553_ (_22977_, _22976_, _22936_);
  and _27554_ (_22978_, _22810_, _22869_);
  not _27555_ (_22979_, _22978_);
  or _27556_ (_22980_, _22979_, _22968_);
  nor _27557_ (_22981_, _22980_, _22844_);
  and _27558_ (_22982_, _22981_, _22977_);
  and _27559_ (_22983_, _22982_, _22974_);
  not _27560_ (_22984_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor _27561_ (_22985_, _22984_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  not _27562_ (_22986_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _27563_ (_22987_, _22986_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand _27564_ (_22988_, _22987_, _22985_);
  and _27565_ (_22989_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _22735_);
  and _27566_ (_22990_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _22735_);
  nor _27567_ (_22991_, _22990_, _22989_);
  not _27568_ (_22992_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _27569_ (_22993_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22735_);
  and _27570_ (_22994_, _22993_, _22992_);
  and _27571_ (_22995_, _22994_, _22991_);
  not _27572_ (_22996_, _22995_);
  not _27573_ (_22997_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _27574_ (_22998_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _27575_ (_22999_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _27576_ (_23000_, _22999_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _27577_ (_23001_, _23000_, _22998_);
  or _27578_ (_23002_, _23001_, _22997_);
  not _27579_ (_23003_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _27580_ (_23004_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _27581_ (_23005_, _23004_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _27582_ (_23006_, _23005_, _23003_);
  and _27583_ (_23007_, _23006_, _23002_);
  not _27584_ (_23008_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or _27585_ (_23009_, _23000_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _27586_ (_23010_, _23009_, _23008_);
  not _27587_ (_23011_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  or _27588_ (_23012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _27589_ (_23013_, _23012_, _22999_);
  or _27590_ (_23015_, _23013_, _23011_);
  and _27591_ (_23016_, _23015_, _23010_);
  and _27592_ (_23017_, _23016_, _23007_);
  or _27593_ (_23018_, _23012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or _27594_ (_23019_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not _27595_ (_23020_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27596_ (_23022_, _23020_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and _27597_ (_23023_, _23022_, _23019_);
  not _27598_ (_23024_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _27599_ (_23025_, _23024_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _27600_ (_23026_, _23025_, _23023_);
  nand _27601_ (_23027_, _23024_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _27602_ (_23028_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _27603_ (_23029_, _23028_, _23026_);
  or _27604_ (_23030_, _23029_, _23018_);
  and _27605_ (_23031_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _27606_ (_23032_, _23031_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _27607_ (_23033_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  not _27608_ (_23034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand _27609_ (_23035_, _23031_, _22998_);
  or _27610_ (_23036_, _23035_, _23034_);
  and _27611_ (_23037_, _23036_, _23033_);
  and _27612_ (_23038_, _23037_, _23030_);
  and _27613_ (_23039_, _23038_, _23017_);
  or _27614_ (_23040_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _27615_ (_23041_, _23040_, _23029_);
  and _27616_ (_23042_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _27617_ (_23043_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not _27618_ (_23044_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _27619_ (_23045_, _23044_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor _27620_ (_23047_, _23045_, _23034_);
  nor _27621_ (_23048_, _23047_, _23043_);
  and _27622_ (_23049_, _23048_, _23041_);
  not _27623_ (_23050_, _23049_);
  and _27624_ (_23051_, _23050_, _23039_);
  nor _27625_ (_23052_, _23049_, _23039_);
  and _27626_ (_23053_, _23049_, _23039_);
  nor _27627_ (_23054_, _23053_, _23052_);
  not _27628_ (_23055_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _27629_ (_23056_, _23001_, _23055_);
  not _27630_ (_23057_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _27631_ (_23058_, _23005_, _23057_);
  and _27632_ (_23059_, _23058_, _23056_);
  not _27633_ (_23060_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or _27634_ (_23061_, _23013_, _23060_);
  not _27635_ (_23062_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or _27636_ (_23063_, _23009_, _23062_);
  and _27637_ (_23064_, _23063_, _23061_);
  and _27638_ (_23065_, _23064_, _23059_);
  or _27639_ (_23066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27640_ (_23067_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23020_);
  and _27641_ (_23068_, _23067_, _23066_);
  or _27642_ (_23069_, _23068_, _23025_);
  or _27643_ (_23070_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _27644_ (_23071_, _23070_, _23069_);
  or _27645_ (_23072_, _23071_, _23018_);
  nand _27646_ (_23073_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  not _27647_ (_23074_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _27648_ (_23075_, _23035_, _23074_);
  and _27649_ (_23076_, _23075_, _23073_);
  and _27650_ (_23078_, _23076_, _23072_);
  and _27651_ (_23079_, _23078_, _23065_);
  or _27652_ (_23080_, _23071_, _23040_);
  nand _27653_ (_23081_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or _27654_ (_23082_, _23045_, _23074_);
  and _27655_ (_23083_, _23082_, _23081_);
  nand _27656_ (_23084_, _23083_, _23080_);
  nor _27657_ (_23085_, _23084_, _23079_);
  not _27658_ (_23086_, _23084_);
  nor _27659_ (_23087_, _23086_, _23079_);
  and _27660_ (_23088_, _23086_, _23079_);
  nor _27661_ (_23089_, _23088_, _23087_);
  not _27662_ (_23090_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or _27663_ (_23091_, _23001_, _23090_);
  not _27664_ (_23092_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _27665_ (_23093_, _23005_, _23092_);
  and _27666_ (_23094_, _23093_, _23091_);
  not _27667_ (_23095_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  or _27668_ (_23096_, _23013_, _23095_);
  not _27669_ (_23097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or _27670_ (_23098_, _23009_, _23097_);
  and _27671_ (_23099_, _23098_, _23096_);
  and _27672_ (_23100_, _23099_, _23094_);
  or _27673_ (_23101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27674_ (_23103_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23020_);
  and _27675_ (_23104_, _23103_, _23101_);
  or _27676_ (_23105_, _23104_, _23025_);
  or _27677_ (_23106_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _27678_ (_23107_, _23106_, _23105_);
  or _27679_ (_23108_, _23107_, _23018_);
  not _27680_ (_23109_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _27681_ (_23111_, _23035_, _23109_);
  nand _27682_ (_23112_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _27683_ (_23113_, _23112_, _23111_);
  and _27684_ (_23114_, _23113_, _23108_);
  nand _27685_ (_23115_, _23114_, _23100_);
  or _27686_ (_23116_, _23107_, _23040_);
  nand _27687_ (_23117_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or _27688_ (_23118_, _23045_, _23109_);
  and _27689_ (_23119_, _23118_, _23117_);
  and _27690_ (_23120_, _23119_, _23116_);
  and _27691_ (_23121_, _23120_, _23115_);
  nand _27692_ (_23122_, _23119_, _23116_);
  and _27693_ (_23123_, _23122_, _23115_);
  nor _27694_ (_23124_, _23122_, _23115_);
  nor _27695_ (_23125_, _23124_, _23123_);
  not _27696_ (_23126_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _27697_ (_23127_, _23001_, _23126_);
  not _27698_ (_23128_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _27699_ (_23129_, _23005_, _23128_);
  and _27700_ (_23130_, _23129_, _23127_);
  not _27701_ (_23131_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or _27702_ (_23132_, _23013_, _23131_);
  not _27703_ (_23133_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or _27704_ (_23134_, _23009_, _23133_);
  and _27705_ (_23136_, _23134_, _23132_);
  and _27706_ (_23137_, _23136_, _23130_);
  or _27707_ (_23138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27708_ (_23139_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23020_);
  and _27709_ (_23140_, _23139_, _23138_);
  or _27710_ (_23141_, _23140_, _23025_);
  or _27711_ (_23142_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _27712_ (_23143_, _23142_, _23141_);
  or _27713_ (_23144_, _23143_, _23018_);
  not _27714_ (_23145_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _27715_ (_23146_, _23035_, _23145_);
  nand _27716_ (_23147_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and _27717_ (_23148_, _23147_, _23146_);
  and _27718_ (_23149_, _23148_, _23144_);
  and _27719_ (_23150_, _23149_, _23137_);
  or _27720_ (_23151_, _23143_, _23040_);
  nand _27721_ (_23152_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or _27722_ (_23154_, _23045_, _23145_);
  and _27723_ (_23155_, _23154_, _23152_);
  nand _27724_ (_23156_, _23155_, _23151_);
  and _27725_ (_23157_, _23156_, _23150_);
  nor _27726_ (_23158_, _23157_, _23125_);
  nor _27727_ (_23159_, _23158_, _23121_);
  nor _27728_ (_23160_, _23159_, _23089_);
  nor _27729_ (_23161_, _23160_, _23085_);
  and _27730_ (_23162_, _23159_, _23089_);
  nor _27731_ (_23163_, _23162_, _23160_);
  not _27732_ (_23164_, _23163_);
  and _27733_ (_23166_, _23157_, _23125_);
  nor _27734_ (_23167_, _23166_, _23158_);
  not _27735_ (_23168_, _23167_);
  and _27736_ (_23169_, _23155_, _23151_);
  nor _27737_ (_23170_, _23169_, _23150_);
  and _27738_ (_23172_, _23169_, _23150_);
  nor _27739_ (_23173_, _23172_, _23170_);
  not _27740_ (_23174_, _23173_);
  not _27741_ (_23175_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _27742_ (_23176_, _23001_, _23175_);
  not _27743_ (_23177_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _27744_ (_23178_, _23005_, _23177_);
  and _27745_ (_23179_, _23178_, _23176_);
  not _27746_ (_23181_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or _27747_ (_23182_, _23013_, _23181_);
  not _27748_ (_23183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or _27749_ (_23184_, _23009_, _23183_);
  and _27750_ (_23185_, _23184_, _23182_);
  and _27751_ (_23186_, _23185_, _23179_);
  or _27752_ (_23187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27753_ (_23188_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23020_);
  and _27754_ (_23189_, _23188_, _23187_);
  or _27755_ (_23190_, _23189_, _23025_);
  or _27756_ (_23191_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _27757_ (_23192_, _23191_, _23190_);
  or _27758_ (_23193_, _23192_, _23018_);
  nand _27759_ (_23194_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not _27760_ (_23195_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _27761_ (_23196_, _23035_, _23195_);
  and _27762_ (_23197_, _23196_, _23194_);
  and _27763_ (_23198_, _23197_, _23193_);
  and _27764_ (_23199_, _23198_, _23186_);
  or _27765_ (_23201_, _23192_, _23040_);
  nand _27766_ (_23202_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or _27767_ (_23203_, _23045_, _23195_);
  and _27768_ (_23204_, _23203_, _23202_);
  and _27769_ (_23205_, _23204_, _23201_);
  and _27770_ (_23206_, _23205_, _23199_);
  nor _27771_ (_23207_, _23205_, _23199_);
  nor _27772_ (_23208_, _23207_, _23206_);
  nand _27773_ (_23209_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not _27774_ (_23210_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _27775_ (_23211_, _23035_, _23210_);
  and _27776_ (_23212_, _23211_, _23209_);
  not _27777_ (_23213_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _27778_ (_23214_, _23001_, _23213_);
  not _27779_ (_23215_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _27780_ (_23216_, _23005_, _23215_);
  and _27781_ (_23217_, _23216_, _23214_);
  and _27782_ (_23218_, _23217_, _23212_);
  or _27783_ (_23219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27784_ (_23220_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23020_);
  and _27785_ (_23221_, _23220_, _23219_);
  or _27786_ (_23222_, _23221_, _23025_);
  or _27787_ (_23223_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _27788_ (_23224_, _23223_, _23222_);
  or _27789_ (_23225_, _23224_, _23018_);
  not _27790_ (_23226_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _27791_ (_23227_, _23009_, _23226_);
  not _27792_ (_23228_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or _27793_ (_23229_, _23013_, _23228_);
  and _27794_ (_23230_, _23229_, _23227_);
  and _27795_ (_23231_, _23230_, _23225_);
  nand _27796_ (_23232_, _23231_, _23218_);
  or _27797_ (_23233_, _23224_, _23040_);
  nand _27798_ (_23234_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _27799_ (_23235_, _23045_, _23210_);
  and _27800_ (_23236_, _23235_, _23234_);
  nand _27801_ (_23237_, _23236_, _23233_);
  and _27802_ (_23238_, _23237_, _23232_);
  nor _27803_ (_23239_, _23237_, _23232_);
  nor _27804_ (_23240_, _23239_, _23238_);
  not _27805_ (_23241_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _27806_ (_23242_, _23001_, _23241_);
  not _27807_ (_23243_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _27808_ (_23244_, _23005_, _23243_);
  and _27809_ (_23245_, _23244_, _23242_);
  not _27810_ (_23246_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or _27811_ (_23247_, _23013_, _23246_);
  not _27812_ (_23248_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _27813_ (_23249_, _23009_, _23248_);
  and _27814_ (_23250_, _23249_, _23247_);
  and _27815_ (_23251_, _23250_, _23245_);
  or _27816_ (_23252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27817_ (_23253_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23020_);
  and _27818_ (_23254_, _23253_, _23252_);
  or _27819_ (_23255_, _23254_, _23025_);
  or _27820_ (_23256_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _27821_ (_23257_, _23256_, _23255_);
  or _27822_ (_23258_, _23257_, _23018_);
  nand _27823_ (_23259_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  not _27824_ (_23260_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _27825_ (_23261_, _23035_, _23260_);
  and _27826_ (_23262_, _23261_, _23259_);
  and _27827_ (_23263_, _23262_, _23258_);
  nand _27828_ (_23264_, _23263_, _23251_);
  or _27829_ (_23265_, _23257_, _23040_);
  nand _27830_ (_23266_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _27831_ (_23267_, _23045_, _23260_);
  and _27832_ (_23268_, _23267_, _23266_);
  nand _27833_ (_23269_, _23268_, _23265_);
  nor _27834_ (_23270_, _23269_, _23264_);
  and _27835_ (_23271_, _23269_, _23264_);
  nor _27836_ (_23272_, _23271_, _23270_);
  not _27837_ (_23273_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _27838_ (_23274_, _23001_, _23273_);
  not _27839_ (_23275_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _27840_ (_23276_, _23005_, _23275_);
  nor _27841_ (_23277_, _23276_, _23274_);
  not _27842_ (_23278_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor _27843_ (_23279_, _23013_, _23278_);
  not _27844_ (_23280_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _27845_ (_23281_, _23009_, _23280_);
  nor _27846_ (_23282_, _23281_, _23279_);
  and _27847_ (_23283_, _23282_, _23277_);
  or _27848_ (_23284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27849_ (_23285_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23020_);
  and _27850_ (_23286_, _23285_, _23284_);
  or _27851_ (_23287_, _23286_, _23025_);
  or _27852_ (_23288_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _27853_ (_23289_, _23288_, _23287_);
  or _27854_ (_23290_, _23289_, _23018_);
  not _27855_ (_23291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _27856_ (_23292_, _23035_, _23291_);
  and _27857_ (_23293_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor _27858_ (_23294_, _23293_, _23292_);
  and _27859_ (_23295_, _23294_, _23290_);
  and _27860_ (_23296_, _23295_, _23283_);
  or _27861_ (_23297_, _23289_, _23040_);
  nand _27862_ (_23298_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or _27863_ (_23299_, _23045_, _23291_);
  and _27864_ (_23300_, _23299_, _23298_);
  nand _27865_ (_23301_, _23300_, _23297_);
  and _27866_ (_23302_, _23301_, _23296_);
  nor _27867_ (_23304_, _23302_, _23272_);
  not _27868_ (_23305_, _23269_);
  and _27869_ (_23306_, _23305_, _23264_);
  nor _27870_ (_23308_, _23306_, _23304_);
  nor _27871_ (_23309_, _23308_, _23240_);
  and _27872_ (_23310_, _23236_, _23233_);
  and _27873_ (_23311_, _23310_, _23232_);
  nor _27874_ (_23312_, _23311_, _23309_);
  nor _27875_ (_23313_, _23312_, _23208_);
  and _27876_ (_23314_, _23312_, _23208_);
  nor _27877_ (_23316_, _23314_, _23313_);
  and _27878_ (_23317_, _23308_, _23240_);
  nor _27879_ (_23318_, _23317_, _23309_);
  not _27880_ (_23319_, _23318_);
  and _27881_ (_23320_, _23302_, _23272_);
  nor _27882_ (_23321_, _23320_, _23304_);
  not _27883_ (_23322_, _23321_);
  not _27884_ (_23323_, _23301_);
  nor _27885_ (_23324_, _23323_, _23296_);
  and _27886_ (_23325_, _23323_, _23296_);
  nor _27887_ (_23327_, _23325_, _23324_);
  and _27888_ (_23328_, _22984_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _27889_ (_23329_, _23068_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _27890_ (_23330_, _23221_, _22986_);
  nand _27891_ (_23331_, _23330_, _23329_);
  nand _27892_ (_23333_, _23331_, _23328_);
  and _27893_ (_23334_, _22985_, _22986_);
  nand _27894_ (_23335_, _23334_, _23254_);
  and _27895_ (_23336_, _22985_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _27896_ (_23337_, _23336_, _23104_);
  and _27897_ (_23338_, _23337_, _23335_);
  and _27898_ (_23340_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _27899_ (_23341_, _23340_, _22986_);
  nand _27900_ (_23342_, _23341_, _23189_);
  and _27901_ (_23343_, _23340_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _27902_ (_23344_, _23343_, _23023_);
  and _27903_ (_23345_, _23344_, _23342_);
  nor _27904_ (_23346_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _27905_ (_23347_, _23346_, _22986_);
  nand _27906_ (_23348_, _23347_, _23286_);
  and _27907_ (_23349_, _23346_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _27908_ (_23350_, _23349_, _23140_);
  and _27909_ (_23351_, _23350_, _23348_);
  and _27910_ (_23352_, _23351_, _23345_);
  and _27911_ (_23353_, _23352_, _23338_);
  nand _27912_ (_23354_, _23353_, _23333_);
  nand _27913_ (_23355_, _23354_, _23027_);
  and _27914_ (_23356_, _23025_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not _27915_ (_23357_, _23356_);
  and _27916_ (_23358_, _23357_, _23355_);
  and _27917_ (_23359_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _27918_ (_23360_, _23359_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor _27919_ (_23361_, _23360_, _23358_);
  not _27920_ (_23362_, _23360_);
  and _27921_ (_23363_, _23362_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _27922_ (_23364_, _23363_, _23361_);
  nor _27923_ (_23366_, _23364_, _23327_);
  and _27924_ (_23367_, _23366_, _23322_);
  and _27925_ (_23368_, _23367_, _23319_);
  not _27926_ (_23369_, _23368_);
  nor _27927_ (_23370_, _23369_, _23316_);
  nand _27928_ (_23371_, _23204_, _23201_);
  or _27929_ (_23372_, _23371_, _23199_);
  and _27930_ (_23373_, _23371_, _23199_);
  or _27931_ (_23374_, _23312_, _23373_);
  and _27932_ (_23375_, _23374_, _23372_);
  or _27933_ (_23376_, _23375_, _23370_);
  and _27934_ (_23377_, _23376_, _23174_);
  and _27935_ (_23378_, _23377_, _23168_);
  and _27936_ (_23379_, _23378_, _23164_);
  nor _27937_ (_23380_, _23379_, _23161_);
  nor _27938_ (_23381_, _23380_, _23054_);
  nor _27939_ (_23382_, _23381_, _23051_);
  nor _27940_ (_23383_, _23382_, _22996_);
  not _27941_ (_23385_, _23383_);
  not _27942_ (_23386_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _27943_ (_23387_, _22735_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _27944_ (_23388_, _23387_, _23386_);
  and _27945_ (_23390_, _23388_, _22991_);
  not _27946_ (_23391_, _23390_);
  not _27947_ (_23392_, _23052_);
  not _27948_ (_23393_, _23054_);
  not _27949_ (_23395_, _23240_);
  and _27950_ (_23396_, _23324_, _23272_);
  nor _27951_ (_23397_, _23396_, _23271_);
  nor _27952_ (_23398_, _23397_, _23395_);
  nor _27953_ (_23399_, _23398_, _23238_);
  nor _27954_ (_23400_, _23399_, _23208_);
  and _27955_ (_23401_, _23399_, _23208_);
  nor _27956_ (_23402_, _23401_, _23400_);
  not _27957_ (_23403_, _23327_);
  nor _27958_ (_23404_, _23364_, _23403_);
  and _27959_ (_23405_, _23404_, _23272_);
  and _27960_ (_23406_, _23397_, _23395_);
  nor _27961_ (_23407_, _23406_, _23398_);
  and _27962_ (_23408_, _23407_, _23405_);
  not _27963_ (_23409_, _23408_);
  nor _27964_ (_23410_, _23409_, _23402_);
  nor _27965_ (_23411_, _23399_, _23206_);
  or _27966_ (_23412_, _23411_, _23207_);
  or _27967_ (_23413_, _23412_, _23410_);
  and _27968_ (_23414_, _23413_, _23173_);
  and _27969_ (_23415_, _23170_, _23125_);
  nor _27970_ (_23416_, _23170_, _23125_);
  nor _27971_ (_23417_, _23416_, _23415_);
  and _27972_ (_23418_, _23417_, _23414_);
  not _27973_ (_23419_, _23089_);
  nor _27974_ (_23420_, _23415_, _23123_);
  nor _27975_ (_23421_, _23420_, _23419_);
  and _27976_ (_23422_, _23420_, _23419_);
  nor _27977_ (_23423_, _23422_, _23421_);
  and _27978_ (_23424_, _23423_, _23418_);
  not _27979_ (_23425_, _23424_);
  nor _27980_ (_23426_, _23421_, _23087_);
  and _27981_ (_23427_, _23426_, _23425_);
  or _27982_ (_23429_, _23427_, _23393_);
  and _27983_ (_23430_, _23429_, _23392_);
  nor _27984_ (_23432_, _23430_, _23391_);
  not _27985_ (_23433_, _23363_);
  not _27986_ (_23434_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _27987_ (_23436_, _22990_, _23434_);
  and _27988_ (_23437_, _23436_, _22994_);
  and _27989_ (_23438_, _23437_, _23433_);
  nor _27990_ (_23439_, _23387_, _22993_);
  and _27991_ (_23440_, _22989_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _27992_ (_23441_, _23440_, _23439_);
  and _27993_ (_23442_, _23441_, _23363_);
  nor _27994_ (_23443_, _23442_, _23438_);
  nor _27995_ (_23444_, _23443_, _23361_);
  not _27996_ (_23445_, _23444_);
  and _27997_ (_23446_, _23433_, _23358_);
  not _27998_ (_23447_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _27999_ (_23448_, _22989_, _23447_);
  and _28000_ (_23449_, _23448_, _23388_);
  and _28001_ (_23450_, _23439_, _23448_);
  not _28002_ (_23451_, _23450_);
  nor _28003_ (_23452_, _23451_, _23361_);
  nor _28004_ (_23453_, _23452_, _23449_);
  nor _28005_ (_23454_, _23453_, _23446_);
  not _28006_ (_23455_, _23454_);
  not _28007_ (_23456_, _23364_);
  not _28008_ (_23457_, _23115_);
  and _28009_ (_23458_, _23457_, _23079_);
  not _28010_ (_23459_, _23458_);
  not _28011_ (_23460_, _23150_);
  and _28012_ (_23461_, _23436_, _23388_);
  nor _28013_ (_23462_, _23264_, _23232_);
  nor _28014_ (_23463_, _23462_, _23199_);
  and _28015_ (_23464_, _23463_, _23461_);
  and _28016_ (_23465_, _23464_, _23460_);
  nor _28017_ (_23466_, _23465_, _23459_);
  nor _28018_ (_23467_, _23466_, _23039_);
  nor _28019_ (_23468_, _23467_, _23456_);
  not _28020_ (_23469_, _23468_);
  not _28021_ (_23470_, _23461_);
  not _28022_ (_23471_, _23466_);
  nor _28023_ (_23472_, _23364_, _23039_);
  and _28024_ (_23473_, _23472_, _23471_);
  nor _28025_ (_23474_, _23473_, _23470_);
  and _28026_ (_23475_, _23474_, _23469_);
  nor _28027_ (_23476_, _23362_, _23358_);
  and _28028_ (_23477_, _23448_, _22994_);
  not _28029_ (_23478_, _23358_);
  and _28030_ (_23479_, _22993_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _28031_ (_23480_, _23479_, _23436_);
  and _28032_ (_23481_, _23480_, _23478_);
  nor _28033_ (_23482_, _23481_, _23477_);
  nor _28034_ (_23483_, _23482_, _23476_);
  and _28035_ (_23484_, _23439_, _22991_);
  and _28036_ (_23485_, _23484_, _23456_);
  not _28037_ (_23486_, _23485_);
  not _28038_ (_23487_, _23039_);
  and _28039_ (_23488_, _23479_, _23448_);
  and _28040_ (_23489_, _23488_, _23487_);
  not _28041_ (_23490_, _23489_);
  not _28042_ (_23491_, _23296_);
  and _28043_ (_23492_, _23440_, _23388_);
  and _28044_ (_23493_, _23492_, _23491_);
  nor _28045_ (_23494_, _23493_, _23464_);
  and _28046_ (_23495_, _23494_, _23490_);
  nand _28047_ (_23496_, _23495_, _23486_);
  or _28048_ (_23497_, _23496_, _23483_);
  nor _28049_ (_23498_, _23497_, _23475_);
  and _28050_ (_23499_, _23498_, _23455_);
  and _28051_ (_23500_, _23499_, _23445_);
  not _28052_ (_23501_, _23500_);
  nor _28053_ (_23503_, _23501_, _23432_);
  and _28054_ (_23504_, _23503_, _23385_);
  nor _28055_ (_23505_, _23504_, _22988_);
  and _28056_ (_23506_, _23440_, _23479_);
  and _28057_ (_23507_, _23506_, _23269_);
  and _28058_ (_23508_, _23491_, _23264_);
  not _28059_ (_23509_, _23264_);
  and _28060_ (_23510_, _23296_, _23509_);
  nor _28061_ (_23511_, _23510_, _23508_);
  not _28062_ (_23512_, _23511_);
  nand _28063_ (_23513_, _23512_, _23364_);
  and _28064_ (_23514_, _23440_, _22994_);
  or _28065_ (_23515_, _23512_, _23364_);
  and _28066_ (_23516_, _23515_, _23514_);
  and _28067_ (_23517_, _23516_, _23513_);
  nor _28068_ (_23518_, _23517_, _23507_);
  and _28069_ (_23519_, _23450_, _23272_);
  not _28070_ (_23520_, _23449_);
  nor _28071_ (_23521_, _23520_, _23270_);
  or _28072_ (_23522_, _23521_, _23519_);
  not _28073_ (_23523_, _23522_);
  and _28074_ (_23524_, _23480_, _23271_);
  and _28075_ (_23525_, _23437_, _23509_);
  nor _28076_ (_23526_, _23525_, _23524_);
  and _28077_ (_23527_, _23526_, _23523_);
  and _28078_ (_23528_, _23439_, _23436_);
  not _28079_ (_23529_, _23528_);
  and _28080_ (_23530_, _23388_, _23434_);
  and _28081_ (_23531_, _23479_, _22991_);
  nor _28082_ (_23532_, _23531_, _23530_);
  and _28083_ (_23533_, _23532_, _23529_);
  and _28084_ (_23534_, _23440_, _23386_);
  and _28085_ (_23535_, _23448_, _22993_);
  or _28086_ (_23536_, _23535_, _23534_);
  nor _28087_ (_23537_, _23536_, _23484_);
  and _28088_ (_23538_, _23537_, _23533_);
  nor _28089_ (_23539_, _23538_, _23509_);
  not _28090_ (_23540_, _23539_);
  and _28091_ (_23541_, _23540_, _23527_);
  and _28092_ (_23542_, _23541_, _23518_);
  nor _28093_ (_23543_, _23542_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28094_ (_23544_, _23334_, _22869_);
  and _28095_ (_23545_, _23544_, _23254_);
  or _28096_ (_23546_, _23545_, _23543_);
  or _28097_ (_23547_, _23546_, _23505_);
  and _28098_ (_23548_, _23547_, _22847_);
  and _28099_ (_23549_, _23548_, _22983_);
  not _28100_ (_23550_, _22983_);
  and _28101_ (_23551_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or _28102_ (_03395_, _23551_, _23549_);
  nand _28103_ (_23552_, _23340_, _22987_);
  nor _28104_ (_23553_, _23552_, _23504_);
  and _28105_ (_23554_, _23450_, _23208_);
  nor _28106_ (_23555_, _23520_, _23206_);
  or _28107_ (_23556_, _23555_, _23554_);
  and _28108_ (_23557_, _23480_, _23207_);
  and _28109_ (_23558_, _23437_, _23199_);
  nor _28110_ (_23559_, _23558_, _23557_);
  not _28111_ (_23560_, _23559_);
  nor _28112_ (_23561_, _23560_, _23556_);
  nor _28113_ (_23562_, _23538_, _23199_);
  not _28114_ (_23563_, _23199_);
  nand _28115_ (_23564_, _23508_, _23232_);
  or _28116_ (_23565_, _23564_, _23456_);
  nand _28117_ (_23566_, _23462_, _23296_);
  or _28118_ (_23567_, _23566_, _23364_);
  nand _28119_ (_23568_, _23567_, _23565_);
  nand _28120_ (_23569_, _23568_, _23563_);
  or _28121_ (_23570_, _23568_, _23563_);
  and _28122_ (_23571_, _23570_, _23514_);
  nand _28123_ (_23572_, _23571_, _23569_);
  and _28124_ (_23573_, _23506_, _23371_);
  not _28125_ (_23574_, _23573_);
  nand _28126_ (_23575_, _23574_, _23572_);
  nor _28127_ (_23576_, _23575_, _23562_);
  nand _28128_ (_23577_, _23576_, _23561_);
  and _28129_ (_23578_, _23577_, _22869_);
  nor _28130_ (_23579_, _23341_, _22869_);
  and _28131_ (_23580_, _23579_, _23189_);
  or _28132_ (_23581_, _23580_, _23578_);
  or _28133_ (_23582_, _23581_, _23553_);
  and _28134_ (_23583_, _23582_, _22847_);
  and _28135_ (_23584_, _23583_, _22983_);
  and _28136_ (_23585_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or _28137_ (_04137_, _23585_, _23584_);
  and _28138_ (_23586_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _28139_ (_23587_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _28140_ (_23588_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _28141_ (_23589_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _28142_ (_23590_, _23589_, _23588_);
  nand _28143_ (_23591_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _28144_ (_23592_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _28145_ (_23593_, _23592_, _23588_);
  nand _28146_ (_23594_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and _28147_ (_23595_, _23594_, _23591_);
  nor _28148_ (_23596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _28149_ (_23597_, _23596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nand _28150_ (_23598_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not _28151_ (_23599_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _28152_ (_23600_, _23599_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _28153_ (_23601_, _23600_, _23588_);
  not _28154_ (_23602_, _23601_);
  nand _28155_ (_23603_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _28156_ (_23604_, _23603_, _23598_);
  nor _28157_ (_23605_, _23589_, _23588_);
  nand _28158_ (_23606_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _28159_ (_23607_, _23589_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _28160_ (_23608_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _28161_ (_23609_, _23608_, _23606_);
  and _28162_ (_23610_, _23609_, _23604_);
  and _28163_ (_23611_, _23610_, _23595_);
  or _28164_ (_23612_, _23611_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _28165_ (_23613_, _23612_, _23587_);
  nor _28166_ (_23614_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _23587_);
  or _28167_ (_23615_, _23614_, _23613_);
  and _28168_ (_23616_, _23615_, _22738_);
  not _28169_ (_23617_, _23616_);
  not _28170_ (_23618_, _22734_);
  nor _28171_ (_23619_, _22737_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _28172_ (_23620_, _23619_, _23618_);
  nand _28173_ (_23621_, _23620_, _23617_);
  not _28174_ (_23622_, _22738_);
  not _28175_ (_23623_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _28176_ (_23624_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and _28177_ (_23625_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _28178_ (_23626_, _23625_, _23624_);
  nand _28179_ (_23627_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand _28180_ (_23628_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _28181_ (_23629_, _23628_, _23627_);
  nand _28182_ (_23630_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand _28183_ (_23631_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _28184_ (_23632_, _23631_, _23630_);
  and _28185_ (_23633_, _23632_, _23629_);
  nand _28186_ (_23634_, _23633_, _23626_);
  nand _28187_ (_23635_, _23634_, _23623_);
  nand _28188_ (_23636_, _23635_, _23587_);
  nor _28189_ (_23637_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _23587_);
  not _28190_ (_23638_, _23637_);
  and _28191_ (_23639_, _23638_, _23636_);
  or _28192_ (_23640_, _23639_, _23622_);
  nor _28193_ (_23641_, _22737_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _28194_ (_23642_, _23641_, _23618_);
  and _28195_ (_23643_, _23642_, _23640_);
  and _28196_ (_23644_, _23643_, _23621_);
  nand _28197_ (_23645_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand _28198_ (_23646_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nand _28199_ (_23647_, _23646_, _23645_);
  and _28200_ (_23648_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _28201_ (_23649_, _23648_, _23647_);
  nand _28202_ (_23650_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _28203_ (_23651_, _23650_, _23623_);
  nand _28204_ (_23652_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _28205_ (_23653_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _28206_ (_23654_, _23653_, _23652_);
  and _28207_ (_23655_, _23654_, _23651_);
  nand _28208_ (_23656_, _23655_, _23649_);
  or _28209_ (_23657_, _23656_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _28210_ (_23658_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _23587_);
  not _28211_ (_23659_, _23658_);
  and _28212_ (_23660_, _23659_, _23657_);
  or _28213_ (_23661_, _23660_, _23622_);
  nor _28214_ (_23662_, _22737_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _28215_ (_23663_, _23662_, _23618_);
  and _28216_ (_23664_, _23663_, _23661_);
  nand _28217_ (_23665_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nand _28218_ (_23666_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _28219_ (_23667_, _23666_, _23665_);
  nand _28220_ (_23668_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _28221_ (_23669_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _28222_ (_23670_, _23669_, _23668_);
  nand _28223_ (_23671_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand _28224_ (_23672_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _28225_ (_23673_, _23672_, _23671_);
  and _28226_ (_23674_, _23673_, _23670_);
  and _28227_ (_23675_, _23674_, _23667_);
  or _28228_ (_23676_, _23675_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _28229_ (_23677_, _23676_, _23587_);
  nor _28230_ (_23679_, _23587_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  not _28231_ (_23680_, _23679_);
  and _28232_ (_23681_, _23680_, _23677_);
  or _28233_ (_23682_, _23681_, _23622_);
  nor _28234_ (_23683_, _22737_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _28235_ (_23684_, _23683_, _23618_);
  and _28236_ (_23685_, _23684_, _23682_);
  nor _28237_ (_23686_, _23685_, _23664_);
  and _28238_ (_23687_, _23686_, _23644_);
  and _28239_ (_23688_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _28240_ (_23689_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _28241_ (_23690_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _28242_ (_23691_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _28243_ (_23692_, _23691_, _23690_);
  and _28244_ (_23693_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and _28245_ (_23694_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _28246_ (_23695_, _23694_, _23693_);
  nand _28247_ (_23696_, _23695_, _23692_);
  or _28248_ (_23697_, _23696_, _23689_);
  or _28249_ (_23698_, _23697_, _23688_);
  or _28250_ (_23699_, _23698_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _28251_ (_23700_, _23699_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _28252_ (_23701_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _23587_);
  not _28253_ (_23702_, _23701_);
  and _28254_ (_23703_, _23702_, _23700_);
  or _28255_ (_23704_, _23703_, _23622_);
  nor _28256_ (_23705_, _22737_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _28257_ (_23706_, _23705_, _23618_);
  and _28258_ (_23707_, _23706_, _23704_);
  not _28259_ (_23708_, _23707_);
  nand _28260_ (_23709_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand _28261_ (_23710_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _28262_ (_23711_, _23710_, _23709_);
  nand _28263_ (_23712_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _28264_ (_23713_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _28265_ (_23714_, _23713_, _23712_);
  nand _28266_ (_23715_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _28267_ (_23716_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _28268_ (_23717_, _23716_, _23715_);
  and _28269_ (_23718_, _23717_, _23714_);
  nand _28270_ (_23719_, _23718_, _23711_);
  nand _28271_ (_23720_, _23719_, _23623_);
  nand _28272_ (_23721_, _23720_, _23587_);
  nor _28273_ (_23722_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _23587_);
  not _28274_ (_23723_, _23722_);
  and _28275_ (_23724_, _23723_, _23721_);
  or _28276_ (_23726_, _23724_, _23622_);
  nor _28277_ (_23727_, _22737_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _28278_ (_23728_, _23727_, _23618_);
  and _28279_ (_23729_, _23728_, _23726_);
  nand _28280_ (_23730_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand _28281_ (_23731_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _28282_ (_23732_, _23731_, _23730_);
  nand _28283_ (_23733_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nand _28284_ (_23734_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _28285_ (_23735_, _23734_, _23733_);
  and _28286_ (_23736_, _23735_, _23732_);
  nand _28287_ (_23737_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _28288_ (_23738_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _28289_ (_23739_, _23738_, _23737_);
  and _28290_ (_23740_, _23739_, _23736_);
  or _28291_ (_23741_, _23740_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _28292_ (_23742_, _23741_, _23587_);
  nor _28293_ (_23743_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _23587_);
  not _28294_ (_23744_, _23743_);
  and _28295_ (_23745_, _23744_, _23742_);
  or _28296_ (_23746_, _23745_, _23622_);
  nor _28297_ (_23747_, _22737_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _28298_ (_23748_, _23747_, _23618_);
  nand _28299_ (_23749_, _23748_, _23746_);
  nand _28300_ (_23750_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand _28301_ (_23751_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _28302_ (_23752_, _23751_, _23750_);
  nand _28303_ (_23753_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _28304_ (_23754_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _28305_ (_23755_, _23754_, _23753_);
  nand _28306_ (_23756_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _28307_ (_23757_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _28308_ (_23758_, _23757_, _23756_);
  and _28309_ (_23759_, _23758_, _23755_);
  nand _28310_ (_23760_, _23759_, _23752_);
  and _28311_ (_23761_, _23760_, _23623_);
  or _28312_ (_23762_, _23761_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _28313_ (_23763_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _23587_);
  not _28314_ (_23764_, _23763_);
  and _28315_ (_23765_, _23764_, _23762_);
  or _28316_ (_23766_, _23765_, _23622_);
  nor _28317_ (_23767_, _22737_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _28318_ (_23768_, _23767_, _23618_);
  nand _28319_ (_23769_, _23768_, _23766_);
  and _28320_ (_23770_, _23769_, _23749_);
  and _28321_ (_23771_, _23770_, _23729_);
  and _28322_ (_23772_, _23771_, _23708_);
  and _28323_ (_23773_, _23772_, _23687_);
  and _28324_ (_23774_, _23773_, _22735_);
  or _28325_ (_23775_, _23774_, _23586_);
  and _28326_ (_23776_, _23775_, _22731_);
  not _28327_ (_23777_, _23643_);
  and _28328_ (_23778_, _23777_, _23621_);
  and _28329_ (_23779_, _23778_, _23664_);
  and _28330_ (_23780_, _23779_, _23685_);
  and _28331_ (_23781_, _23768_, _23766_);
  and _28332_ (_23782_, _23781_, _23729_);
  and _28333_ (_23783_, _23782_, _23749_);
  and _28334_ (_23784_, _23783_, _23707_);
  and _28335_ (_23785_, _23784_, _23780_);
  and _28336_ (_23786_, _23748_, _23746_);
  and _28337_ (_23788_, _23782_, _23786_);
  and _28338_ (_23789_, _23788_, _23707_);
  and _28339_ (_23790_, _23789_, _23687_);
  not _28340_ (_23791_, _23685_);
  and _28341_ (_23792_, _23779_, _23791_);
  and _28342_ (_23793_, _23792_, _23784_);
  or _28343_ (_23794_, _23793_, _23790_);
  or _28344_ (_23795_, _23794_, _23785_);
  not _28345_ (_23796_, _23664_);
  and _28346_ (_23797_, _23796_, _23644_);
  not _28347_ (_23798_, _23729_);
  and _28348_ (_23799_, _23749_, _23798_);
  and _28349_ (_23800_, _23799_, _23769_);
  and _28350_ (_23801_, _23800_, _23708_);
  and _28351_ (_23802_, _23685_, _23796_);
  and _28352_ (_23803_, _23802_, _23644_);
  and _28353_ (_23804_, _23769_, _23786_);
  and _28354_ (_23805_, _23804_, _23729_);
  and _28355_ (_23806_, _23805_, _23707_);
  and _28356_ (_23807_, _23806_, _23803_);
  or _28357_ (_23808_, _23807_, _23801_);
  and _28358_ (_23809_, _23808_, _23797_);
  and _28359_ (_23810_, _23786_, _23798_);
  and _28360_ (_23811_, _23810_, _23769_);
  and _28361_ (_23812_, _23811_, _23707_);
  and _28362_ (_23813_, _23664_, _23643_);
  and _28363_ (_23814_, _23813_, _23621_);
  and _28364_ (_23815_, _23814_, _23812_);
  and _28365_ (_23816_, _23778_, _23686_);
  and _28366_ (_23817_, _23816_, _23784_);
  and _28367_ (_23818_, _23800_, _23707_);
  and _28368_ (_23819_, _23818_, _23797_);
  or _28369_ (_23820_, _23819_, _23817_);
  or _28370_ (_23821_, _23820_, _23815_);
  or _28371_ (_23822_, _23821_, _23809_);
  or _28372_ (_23823_, _23822_, _23795_);
  not _28373_ (_23824_, _23621_);
  and _28374_ (_23825_, _23707_, _23824_);
  and _28375_ (_23826_, _23825_, _23811_);
  or _28376_ (_23827_, _23806_, _23800_);
  and _28377_ (_23828_, _23827_, _23824_);
  nor _28378_ (_23829_, _23828_, _23826_);
  and _28379_ (_23830_, _23812_, _23779_);
  and _28380_ (_23831_, _23792_, _23772_);
  or _28381_ (_23832_, _23831_, _23830_);
  and _28382_ (_23833_, _23812_, _23797_);
  nor _28383_ (_23834_, _23833_, _23832_);
  nand _28384_ (_23835_, _23834_, _23829_);
  and _28385_ (_23836_, _23799_, _23780_);
  and _28386_ (_23837_, _23836_, _23769_);
  nor _28387_ (_23838_, _23707_, _23621_);
  and _28388_ (_23839_, _23838_, _23805_);
  and _28389_ (_23840_, _23814_, _23800_);
  and _28390_ (_23841_, _23814_, _23805_);
  or _28391_ (_23842_, _23841_, _23840_);
  or _28392_ (_23843_, _23842_, _23839_);
  and _28393_ (_23844_, _23805_, _23708_);
  and _28394_ (_23845_, _23844_, _23803_);
  and _28395_ (_23846_, _23806_, _23687_);
  or _28396_ (_23847_, _23846_, _23845_);
  or _28397_ (_23848_, _23847_, _23843_);
  or _28398_ (_23850_, _23848_, _23837_);
  or _28399_ (_23851_, _23850_, _23835_);
  or _28400_ (_23853_, _23851_, _23823_);
  nor _28401_ (_23854_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and _28402_ (_23855_, _23854_, _22736_);
  and _28403_ (_23856_, _23855_, _23853_);
  or _28404_ (_26851_[2], _23856_, _23776_);
  nand _28405_ (_23857_, _23328_, _22987_);
  nor _28406_ (_23858_, _23857_, _23504_);
  and _28407_ (_23859_, _23506_, _23237_);
  or _28408_ (_23860_, _23510_, _23364_);
  or _28409_ (_23861_, _23508_, _23456_);
  and _28410_ (_23862_, _23861_, _23860_);
  nand _28411_ (_23863_, _23862_, _23232_);
  or _28412_ (_23864_, _23862_, _23232_);
  and _28413_ (_23865_, _23864_, _23514_);
  and _28414_ (_23867_, _23865_, _23863_);
  nor _28415_ (_23868_, _23867_, _23859_);
  and _28416_ (_23869_, _23450_, _23240_);
  and _28417_ (_23870_, _23480_, _23238_);
  nor _28418_ (_23871_, _23520_, _23239_);
  not _28419_ (_23872_, _23232_);
  and _28420_ (_23873_, _23437_, _23872_);
  or _28421_ (_23874_, _23873_, _23871_);
  or _28422_ (_23875_, _23874_, _23870_);
  nor _28423_ (_23876_, _23875_, _23869_);
  nor _28424_ (_23877_, _23538_, _23872_);
  not _28425_ (_23878_, _23877_);
  and _28426_ (_23879_, _23878_, _23876_);
  nand _28427_ (_23880_, _23879_, _23868_);
  and _28428_ (_23881_, _23880_, _22869_);
  nand _28429_ (_23882_, _23328_, _22986_);
  and _28430_ (_23883_, _23221_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _28431_ (_23884_, _23883_, _23882_);
  or _28432_ (_23885_, _23884_, _23881_);
  or _28433_ (_23886_, _23885_, _23858_);
  and _28434_ (_23887_, _23886_, _22847_);
  and _28435_ (_23888_, _23887_, _22983_);
  and _28436_ (_23889_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or _28437_ (_06732_, _23889_, _23888_);
  and _28438_ (_23890_, \oc8051_top_1.oc8051_sfr1.wait_data , _22731_);
  and _28439_ (_23891_, _23890_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and _28440_ (_23892_, _23783_, _23708_);
  and _28441_ (_23893_, _23892_, _23792_);
  and _28442_ (_23894_, _23844_, _23780_);
  or _28443_ (_23895_, _23894_, _23893_);
  or _28444_ (_23896_, _23813_, _23824_);
  and _28445_ (_23897_, _23896_, _23784_);
  and _28446_ (_23898_, _23797_, _23784_);
  or _28447_ (_23899_, _23898_, _23897_);
  or _28448_ (_23900_, _23899_, _23895_);
  or _28449_ (_23901_, _23846_, _23785_);
  nor _28450_ (_23902_, _23831_, _23817_);
  and _28451_ (_23903_, _23799_, _23781_);
  and _28452_ (_23904_, _23903_, _23780_);
  nand _28453_ (_23905_, _23904_, _23707_);
  nand _28454_ (_23906_, _23905_, _23902_);
  or _28455_ (_23907_, _23906_, _23901_);
  or _28456_ (_23908_, _23907_, _23900_);
  and _28457_ (_23909_, _23814_, _23707_);
  and _28458_ (_23910_, _23909_, _23771_);
  and _28459_ (_23911_, _23771_, _23707_);
  and _28460_ (_23912_, _23911_, _23797_);
  or _28461_ (_23913_, _23912_, _23910_);
  and _28462_ (_23914_, _23903_, _23814_);
  and _28463_ (_23915_, _23825_, _23770_);
  and _28464_ (_23916_, _23915_, _23729_);
  or _28465_ (_23917_, _23916_, _23914_);
  and _28466_ (_23918_, _23903_, _23824_);
  and _28467_ (_23919_, _23903_, _23797_);
  or _28468_ (_23920_, _23919_, _23918_);
  or _28469_ (_23921_, _23920_, _23917_);
  or _28470_ (_23922_, _23921_, _23913_);
  and _28471_ (_23923_, _23806_, _23779_);
  and _28472_ (_23924_, _23923_, _23685_);
  and _28473_ (_23925_, _23818_, _23780_);
  and _28474_ (_23926_, _23810_, _23781_);
  and _28475_ (_23927_, _23926_, _23707_);
  and _28476_ (_23928_, _23927_, _23792_);
  and _28477_ (_23929_, _23816_, _23783_);
  and _28478_ (_23930_, _23929_, _23708_);
  nor _28479_ (_23931_, _23930_, _23928_);
  not _28480_ (_23932_, _23931_);
  or _28481_ (_23933_, _23932_, _23925_);
  or _28482_ (_23934_, _23933_, _23924_);
  or _28483_ (_23935_, _23934_, _23922_);
  or _28484_ (_23936_, _23935_, _23908_);
  and _28485_ (_23937_, _23936_, _23855_);
  or _28486_ (_26852_[0], _23937_, _23891_);
  and _28487_ (_23938_, _22922_, _22888_);
  nor _28488_ (_23939_, _22972_, _22849_);
  and _28489_ (_23940_, _23939_, _22953_);
  and _28490_ (_23941_, _23940_, _23938_);
  and _28491_ (_23943_, _22976_, _22937_);
  and _28492_ (_23944_, _22968_, _22844_);
  and _28493_ (_23945_, _23944_, _23943_);
  and _28494_ (_23946_, _23945_, _23941_);
  and _28495_ (_23947_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand _28496_ (_23948_, _23947_, _23340_);
  nor _28497_ (_23950_, _23948_, _23504_);
  nor _28498_ (_23951_, _23538_, _23039_);
  not _28499_ (_23952_, _23951_);
  not _28500_ (_23953_, _23514_);
  nor _28501_ (_23954_, _23566_, _23563_);
  and _28502_ (_23955_, _23954_, _23150_);
  and _28503_ (_23957_, _23955_, _23458_);
  nor _28504_ (_23958_, _23957_, _23364_);
  not _28505_ (_23959_, _23079_);
  nor _28506_ (_23960_, _23564_, _23199_);
  and _28507_ (_23962_, _23960_, _23460_);
  and _28508_ (_23963_, _23962_, _23115_);
  and _28509_ (_23964_, _23963_, _23959_);
  nor _28510_ (_23965_, _23964_, _23456_);
  or _28511_ (_23966_, _23965_, _23958_);
  nor _28512_ (_23967_, _23966_, _23487_);
  and _28513_ (_23968_, _23966_, _23487_);
  nor _28514_ (_23969_, _23968_, _23967_);
  nor _28515_ (_23970_, _23969_, _23953_);
  nor _28516_ (_23971_, _23364_, _23050_);
  not _28517_ (_23973_, _23971_);
  not _28518_ (_23974_, _23506_);
  and _28519_ (_23975_, _23364_, _23039_);
  nor _28520_ (_23976_, _23975_, _23974_);
  and _28521_ (_23977_, _23976_, _23973_);
  and _28522_ (_23978_, _23450_, _23054_);
  and _28523_ (_23979_, _23480_, _23052_);
  nor _28524_ (_23980_, _23520_, _23053_);
  and _28525_ (_23981_, _23437_, _23039_);
  or _28526_ (_23982_, _23981_, _23980_);
  or _28527_ (_23983_, _23982_, _23979_);
  nor _28528_ (_23984_, _23983_, _23978_);
  not _28529_ (_23985_, _23984_);
  nor _28530_ (_23986_, _23985_, _23977_);
  not _28531_ (_23987_, _23986_);
  nor _28532_ (_23988_, _23987_, _23970_);
  and _28533_ (_23989_, _23988_, _23952_);
  nor _28534_ (_23990_, _23989_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28535_ (_23991_, _23343_, _22869_);
  and _28536_ (_23992_, _23991_, _23023_);
  or _28537_ (_23994_, _23992_, _23990_);
  or _28538_ (_23995_, _23994_, _23950_);
  and _28539_ (_23996_, _23995_, _22847_);
  and _28540_ (_23997_, _23996_, _23946_);
  not _28541_ (_23998_, _23946_);
  and _28542_ (_23999_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or _28543_ (_09147_, _23999_, _23997_);
  nor _28544_ (_24000_, _22937_, _22871_);
  not _28545_ (_24001_, _24000_);
  and _28546_ (_24002_, _24001_, _22847_);
  nor _28547_ (_24003_, _24002_, _22976_);
  and _28548_ (_24004_, _22969_, _22844_);
  and _28549_ (_24005_, _24004_, _22847_);
  and _28550_ (_24006_, _24005_, _24003_);
  and _28551_ (_24008_, _24006_, _23941_);
  and _28552_ (_24009_, _24008_, _23996_);
  not _28553_ (_24011_, _24008_);
  and _28554_ (_24013_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or _28555_ (_13109_, _24013_, _24009_);
  and _28556_ (_24014_, _22921_, _22890_);
  and _28557_ (_24015_, _23939_, _22954_);
  and _28558_ (_24016_, _24015_, _24014_);
  and _28559_ (_24017_, _24016_, _23945_);
  nand _28560_ (_24018_, _23947_, _22985_);
  nor _28561_ (_24019_, _24018_, _23504_);
  and _28562_ (_24020_, _23364_, _23457_);
  not _28563_ (_24021_, _24020_);
  nor _28564_ (_24022_, _23364_, _23122_);
  nor _28565_ (_24023_, _24022_, _23974_);
  and _28566_ (_24024_, _24023_, _24021_);
  nor _28567_ (_24025_, _23962_, _23456_);
  nor _28568_ (_24026_, _23955_, _23364_);
  nor _28569_ (_24027_, _24026_, _24025_);
  nor _28570_ (_24028_, _24027_, _23115_);
  and _28571_ (_24029_, _24027_, _23115_);
  or _28572_ (_24030_, _24029_, _23953_);
  nor _28573_ (_24031_, _24030_, _24028_);
  nor _28574_ (_24032_, _24031_, _24024_);
  and _28575_ (_24033_, _23450_, _23125_);
  and _28576_ (_24034_, _23480_, _23123_);
  nor _28577_ (_24035_, _23520_, _23124_);
  and _28578_ (_24036_, _23437_, _23457_);
  or _28579_ (_24037_, _24036_, _24035_);
  or _28580_ (_24038_, _24037_, _24034_);
  nor _28581_ (_24039_, _24038_, _24033_);
  nor _28582_ (_24040_, _23538_, _23457_);
  not _28583_ (_24041_, _24040_);
  and _28584_ (_24042_, _24041_, _24039_);
  and _28585_ (_24043_, _24042_, _24032_);
  nor _28586_ (_24044_, _24043_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28587_ (_24045_, _23336_, _22869_);
  and _28588_ (_24047_, _24045_, _23104_);
  or _28589_ (_24048_, _24047_, _24044_);
  or _28590_ (_24050_, _24048_, _24019_);
  and _28591_ (_24051_, _24050_, _22847_);
  and _28592_ (_24052_, _24051_, _24017_);
  not _28593_ (_24053_, _24017_);
  and _28594_ (_24054_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or _28595_ (_18267_, _24054_, _24052_);
  and _28596_ (_24055_, _22922_, _22890_);
  and _28597_ (_24056_, _24055_, _22973_);
  and _28598_ (_24057_, _24056_, _22982_);
  nand _28599_ (_24058_, _23947_, _23346_);
  nor _28600_ (_24059_, _24058_, _23504_);
  nand _28601_ (_24060_, _23960_, _23364_);
  nand _28602_ (_24061_, _23954_, _23456_);
  and _28603_ (_24062_, _24061_, _24060_);
  or _28604_ (_24063_, _24062_, _23150_);
  nand _28605_ (_24064_, _24062_, _23150_);
  and _28606_ (_24065_, _24064_, _24063_);
  nand _28607_ (_24066_, _24065_, _23514_);
  and _28608_ (_24067_, _23364_, _23150_);
  nor _28609_ (_24068_, _23364_, _23156_);
  or _28610_ (_24069_, _24068_, _23974_);
  nor _28611_ (_24070_, _24069_, _24067_);
  not _28612_ (_24071_, _24070_);
  and _28613_ (_24072_, _24071_, _24066_);
  and _28614_ (_24073_, _23480_, _23170_);
  and _28615_ (_24074_, _23437_, _23150_);
  nor _28616_ (_24075_, _24074_, _24073_);
  nor _28617_ (_24076_, _23538_, _23150_);
  and _28618_ (_24077_, _23450_, _23173_);
  nor _28619_ (_24078_, _23520_, _23172_);
  or _28620_ (_24079_, _24078_, _24077_);
  nor _28621_ (_24080_, _24079_, _24076_);
  and _28622_ (_24081_, _24080_, _24075_);
  and _28623_ (_24082_, _24081_, _24072_);
  nor _28624_ (_24083_, _24082_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28625_ (_24085_, _23349_, _22869_);
  and _28626_ (_24086_, _24085_, _23140_);
  or _28627_ (_24087_, _24086_, _24083_);
  or _28628_ (_24088_, _24087_, _24059_);
  and _28629_ (_24089_, _24088_, _22847_);
  and _28630_ (_24091_, _24089_, _24057_);
  not _28631_ (_24092_, _24057_);
  and _28632_ (_24093_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or _28633_ (_27284_, _24093_, _24091_);
  nor _28634_ (_24094_, _23939_, _22954_);
  and _28635_ (_24095_, _24094_, _24055_);
  not _28636_ (_24096_, _22975_);
  and _28637_ (_24097_, _24002_, _24096_);
  and _28638_ (_24098_, _24097_, _22981_);
  and _28639_ (_24099_, _24098_, _24095_);
  nand _28640_ (_24100_, _23947_, _23328_);
  nor _28641_ (_24101_, _24100_, _23504_);
  nor _28642_ (_24102_, _23364_, _23086_);
  and _28643_ (_24104_, _23364_, _23959_);
  nor _28644_ (_24105_, _24104_, _24102_);
  nor _28645_ (_24106_, _24105_, _23974_);
  or _28646_ (_24107_, _23963_, _23959_);
  and _28647_ (_24108_, _24107_, _23965_);
  and _28648_ (_24109_, _23955_, _23457_);
  nor _28649_ (_24110_, _24109_, _23079_);
  or _28650_ (_24111_, _24110_, _23957_);
  and _28651_ (_24112_, _24111_, _23456_);
  or _28652_ (_24113_, _24112_, _24108_);
  and _28653_ (_24114_, _24113_, _23514_);
  nor _28654_ (_24115_, _24114_, _24106_);
  and _28655_ (_24116_, _23450_, _23089_);
  and _28656_ (_24117_, _23480_, _23087_);
  nor _28657_ (_24118_, _23520_, _23088_);
  and _28658_ (_24119_, _23437_, _23079_);
  or _28659_ (_24120_, _24119_, _24118_);
  or _28660_ (_24121_, _24120_, _24117_);
  nor _28661_ (_24122_, _24121_, _24116_);
  nor _28662_ (_24123_, _23538_, _23079_);
  not _28663_ (_24124_, _24123_);
  and _28664_ (_24125_, _24124_, _24122_);
  and _28665_ (_24126_, _24125_, _24115_);
  nor _28666_ (_24127_, _24126_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand _28667_ (_24129_, _23328_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _28668_ (_24130_, _23068_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _28669_ (_24131_, _24130_, _24129_);
  or _28670_ (_24132_, _24131_, _24127_);
  or _28671_ (_24133_, _24132_, _24101_);
  and _28672_ (_24134_, _24133_, _22847_);
  and _28673_ (_24136_, _24134_, _24099_);
  not _28674_ (_24137_, _24099_);
  and _28675_ (_24139_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _28676_ (_27310_, _24139_, _24136_);
  and _28677_ (_24140_, _24094_, _22923_);
  and _28678_ (_24141_, _23943_, _22981_);
  and _28679_ (_24142_, _24141_, _24140_);
  and _28680_ (_24143_, _24142_, _23548_);
  not _28681_ (_24144_, _24142_);
  and _28682_ (_24145_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or _28683_ (_22611_, _24145_, _24143_);
  and _28684_ (_24146_, _24094_, _24014_);
  and _28685_ (_24147_, _24146_, _24141_);
  and _28686_ (_24148_, _24147_, _23548_);
  not _28687_ (_24149_, _24147_);
  and _28688_ (_24150_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _28689_ (_22616_, _24150_, _24148_);
  and _28690_ (_24151_, _24142_, _24134_);
  and _28691_ (_24152_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or _28692_ (_22620_, _24152_, _24151_);
  and _28693_ (_24153_, _24147_, _23887_);
  and _28694_ (_24154_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _28695_ (_22688_, _24154_, _24153_);
  and _28696_ (_24155_, _24095_, _22982_);
  and _28697_ (_24156_, _24155_, _24051_);
  not _28698_ (_24157_, _24155_);
  and _28699_ (_24158_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or _28700_ (_22689_, _24158_, _24156_);
  and _28701_ (_24159_, _24055_, _24015_);
  and _28702_ (_24160_, _24159_, _24098_);
  and _28703_ (_24161_, _24160_, _23887_);
  not _28704_ (_24162_, _24160_);
  and _28705_ (_24163_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or _28706_ (_23787_, _24163_, _24161_);
  and _28707_ (_24164_, _24147_, _23996_);
  and _28708_ (_24165_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _28709_ (_23949_, _24165_, _24164_);
  and _28710_ (_24166_, _24147_, _24089_);
  and _28711_ (_24167_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _28712_ (_23972_, _24167_, _24166_);
  and _28713_ (_24169_, _23946_, _23548_);
  and _28714_ (_24170_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or _28715_ (_23993_, _24170_, _24169_);
  and _28716_ (_24171_, _24147_, _24051_);
  and _28717_ (_24172_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _28718_ (_26923_, _24172_, _24171_);
  and _28719_ (_24173_, _22936_, _22905_);
  and _28720_ (_24174_, _24173_, _23944_);
  not _28721_ (_24175_, _22886_);
  and _28722_ (_24176_, _22951_, _22919_);
  and _28723_ (_24177_, _24176_, _24175_);
  nor _28724_ (_24178_, _22814_, _22811_);
  and _28725_ (_24179_, _24178_, _22869_);
  not _28726_ (_24180_, _24179_);
  nor _28727_ (_24181_, _24180_, _22867_);
  and _28728_ (_24182_, _24181_, _24177_);
  and _28729_ (_24184_, _24182_, _24174_);
  or _28730_ (_24185_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _28731_ (_24186_, _24185_, _22731_);
  and _28732_ (_24187_, _24177_, _22868_);
  and _28733_ (_24188_, _24174_, _24179_);
  and _28734_ (_24189_, _24188_, _24187_);
  nand _28735_ (_24190_, _24189_, _24126_);
  and _28736_ (_24427_, _24190_, _24186_);
  nand _28737_ (_24192_, _23346_, _22987_);
  nor _28738_ (_24193_, _24192_, _23504_);
  nor _28739_ (_24194_, _23451_, _23324_);
  nor _28740_ (_24196_, _24194_, _23449_);
  or _28741_ (_24197_, _24196_, _23325_);
  and _28742_ (_24198_, _23480_, _23324_);
  and _28743_ (_24200_, _23437_, _23296_);
  nor _28744_ (_24201_, _24200_, _24198_);
  and _28745_ (_24203_, _23506_, _23301_);
  and _28746_ (_24204_, _23514_, _23296_);
  nor _28747_ (_24206_, _24204_, _24203_);
  or _28748_ (_24207_, _23538_, _23296_);
  and _28749_ (_24208_, _24207_, _24206_);
  and _28750_ (_24209_, _24208_, _24201_);
  and _28751_ (_24210_, _24209_, _24197_);
  nor _28752_ (_24212_, _24210_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand _28753_ (_24214_, _23286_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28754_ (_24216_, _24214_, _23347_);
  or _28755_ (_24217_, _24216_, _24212_);
  or _28756_ (_24218_, _24217_, _24193_);
  and _28757_ (_24219_, _24218_, _22847_);
  and _28758_ (_24220_, _24219_, _23946_);
  and _28759_ (_24221_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or _28760_ (_27056_, _24221_, _24220_);
  and _28761_ (_24223_, _23938_, _22973_);
  and _28762_ (_24224_, _24223_, _22982_);
  and _28763_ (_24225_, _24224_, _23996_);
  not _28764_ (_24226_, _24224_);
  and _28765_ (_24228_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _28766_ (_24683_, _24228_, _24225_);
  and _28767_ (_24229_, _24224_, _24134_);
  and _28768_ (_24230_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _28769_ (_24796_, _24230_, _24229_);
  and _28770_ (_24231_, _24224_, _24051_);
  and _28771_ (_24232_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _28772_ (_24901_, _24232_, _24231_);
  and _28773_ (_24233_, _24134_, _24008_);
  and _28774_ (_24234_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _28775_ (_25095_, _24234_, _24233_);
  and _28776_ (_24236_, _24015_, _22923_);
  and _28777_ (_24237_, _24236_, _23945_);
  and _28778_ (_24238_, _24237_, _24089_);
  not _28779_ (_24239_, _24237_);
  and _28780_ (_24240_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _28781_ (_25114_, _24240_, _24238_);
  and _28782_ (_24243_, _23890_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _28783_ (_24244_, _23892_, _23687_);
  or _28784_ (_24245_, _24244_, _23833_);
  and _28785_ (_24246_, _23780_, _23771_);
  and _28786_ (_24247_, _23903_, _23707_);
  and _28787_ (_24248_, _24247_, _23797_);
  or _28788_ (_24249_, _24248_, _24246_);
  or _28789_ (_24250_, _24249_, _24245_);
  and _28790_ (_24251_, _23927_, _23780_);
  and _28791_ (_24253_, _23892_, _23780_);
  nor _28792_ (_24254_, _24253_, _24251_);
  not _28793_ (_24255_, _24254_);
  and _28794_ (_24257_, _23811_, _23708_);
  and _28795_ (_24258_, _24257_, _23687_);
  and _28796_ (_24259_, _24257_, _23779_);
  nor _28797_ (_24260_, _24259_, _23928_);
  not _28798_ (_24261_, _24260_);
  or _28799_ (_24262_, _24261_, _24258_);
  or _28800_ (_24263_, _24262_, _24255_);
  or _28801_ (_24264_, _24263_, _24250_);
  nor _28802_ (_24265_, _23831_, _23830_);
  nand _28803_ (_24266_, _23905_, _24265_);
  or _28804_ (_24267_, _23918_, _23826_);
  and _28805_ (_24268_, _23909_, _23811_);
  or _28806_ (_24269_, _23914_, _24268_);
  or _28807_ (_24270_, _24269_, _24267_);
  or _28808_ (_24271_, _24270_, _24266_);
  and _28809_ (_24272_, _23903_, _23708_);
  and _28810_ (_24273_, _24272_, _23797_);
  and _28811_ (_24274_, _24257_, _23803_);
  and _28812_ (_24275_, _23844_, _23797_);
  or _28813_ (_24276_, _24275_, _24274_);
  or _28814_ (_24277_, _24276_, _24273_);
  or _28815_ (_24278_, _22736_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _28816_ (_24279_, _24278_);
  and _28817_ (_24281_, _23838_, _23804_);
  or _28818_ (_24283_, _24281_, _24279_);
  or _28819_ (_24284_, _24283_, _23841_);
  or _28820_ (_24286_, _24284_, _23846_);
  and _28821_ (_24287_, _24257_, _23814_);
  or _28822_ (_24289_, _24287_, _23925_);
  or _28823_ (_24290_, _24289_, _24286_);
  or _28824_ (_24291_, _24290_, _24277_);
  or _28825_ (_24292_, _24291_, _24271_);
  or _28826_ (_24293_, _24292_, _24264_);
  or _28827_ (_24294_, _24244_, _24278_);
  and _28828_ (_24295_, _24294_, _23854_);
  and _28829_ (_24296_, _24295_, _24293_);
  or _28830_ (_26851_[0], _24296_, _24243_);
  and _28831_ (_24297_, _24015_, _23938_);
  nor _28832_ (_24298_, _22969_, _22844_);
  nor _28833_ (_24299_, _24298_, _22871_);
  not _28834_ (_24300_, _24299_);
  and _28835_ (_24301_, _24300_, _23943_);
  and _28836_ (_24302_, _24301_, _24297_);
  and _28837_ (_24303_, _24302_, _23548_);
  not _28838_ (_24304_, _24302_);
  and _28839_ (_24305_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or _28840_ (_25352_, _24305_, _24303_);
  and _28841_ (_24306_, _24057_, _23887_);
  and _28842_ (_24307_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or _28843_ (_25419_, _24307_, _24306_);
  and _28844_ (_24308_, _24057_, _23548_);
  and _28845_ (_24309_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or _28846_ (_25474_, _24309_, _24308_);
  and _28847_ (_24310_, _23946_, _23583_);
  and _28848_ (_24311_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or _28849_ (_25595_, _24311_, _24310_);
  and _28850_ (_24312_, _24219_, _24057_);
  and _28851_ (_24313_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or _28852_ (_25624_, _24313_, _24312_);
  and _28853_ (_24314_, _24237_, _24134_);
  and _28854_ (_24315_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _28855_ (_27064_, _24315_, _24314_);
  and _28856_ (_24317_, _23946_, _23887_);
  and _28857_ (_24318_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or _28858_ (_25749_, _24318_, _24317_);
  and _28859_ (_24319_, _24014_, _22973_);
  and _28860_ (_24320_, _24319_, _22982_);
  and _28861_ (_24321_, _24320_, _24134_);
  not _28862_ (_24322_, _24320_);
  and _28863_ (_24323_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _28864_ (_25824_, _24323_, _24321_);
  and _28865_ (_24324_, _24224_, _24219_);
  and _28866_ (_24325_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _28867_ (_25843_, _24325_, _24324_);
  and _28868_ (_24327_, _24320_, _23996_);
  and _28869_ (_24328_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _28870_ (_25943_, _24328_, _24327_);
  and _28871_ (_24330_, _24223_, _23945_);
  and _28872_ (_24331_, _24330_, _23548_);
  not _28873_ (_24332_, _24330_);
  and _28874_ (_24333_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _28875_ (_26134_, _24333_, _24331_);
  or _28876_ (_24334_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _28877_ (_24336_, _24334_, _22731_);
  nand _28878_ (_24337_, _24189_, _24082_);
  and _28879_ (_26179_, _24337_, _24336_);
  and _28880_ (_24339_, _24330_, _24219_);
  and _28881_ (_24340_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _28882_ (_26270_, _24340_, _24339_);
  and _28883_ (_24341_, _24224_, _23583_);
  and _28884_ (_24342_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _28885_ (_27282_, _24342_, _24341_);
  and _28886_ (_24343_, _24224_, _23887_);
  and _28887_ (_24345_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _28888_ (_27281_, _24345_, _24343_);
  and _28889_ (_24347_, _24224_, _23548_);
  and _28890_ (_24348_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _28891_ (_27280_, _24348_, _24347_);
  and _28892_ (_24349_, _24055_, _23940_);
  and _28893_ (_24350_, _24349_, _23945_);
  and _28894_ (_24351_, _24350_, _24051_);
  not _28895_ (_24352_, _24350_);
  and _28896_ (_24353_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _28897_ (_27061_, _24353_, _24351_);
  and _28898_ (_24354_, _24330_, _24089_);
  and _28899_ (_24355_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _28900_ (_27049_, _24355_, _24354_);
  and _28901_ (_24357_, _24320_, _24089_);
  and _28902_ (_24358_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _28903_ (_27278_, _24358_, _24357_);
  and _28904_ (_24360_, _24330_, _23583_);
  and _28905_ (_24361_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _28906_ (_27048_, _24361_, _24360_);
  and _28907_ (_24362_, _24330_, _23887_);
  and _28908_ (_24364_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _28909_ (_27047_, _24364_, _24362_);
  and _28910_ (_24365_, _24300_, _24097_);
  and _28911_ (_24367_, _24365_, _24349_);
  and _28912_ (_24368_, _24367_, _23996_);
  not _28913_ (_24369_, _24367_);
  and _28914_ (_24371_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or _28915_ (_27202_, _24371_, _24368_);
  and _28916_ (_24372_, _24094_, _23938_);
  and _28917_ (_24373_, _24372_, _22982_);
  and _28918_ (_24374_, _24373_, _23887_);
  not _28919_ (_24375_, _24373_);
  and _28920_ (_24376_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _28921_ (_27270_, _24376_, _24374_);
  and _28922_ (_24377_, _24373_, _23548_);
  and _28923_ (_24378_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _28924_ (_27269_, _24378_, _24377_);
  and _28925_ (_24379_, _24373_, _24219_);
  and _28926_ (_24380_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _28927_ (_27268_, _24380_, _24379_);
  and _28928_ (_24381_, _24319_, _23945_);
  and _28929_ (_24382_, _24381_, _23887_);
  not _28930_ (_24383_, _24381_);
  and _28931_ (_24384_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _28932_ (_27043_, _24384_, _24382_);
  and _28933_ (_24385_, _24381_, _23583_);
  and _28934_ (_24386_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _28935_ (_27044_, _24386_, _24385_);
  and _28936_ (_24387_, _24373_, _24051_);
  and _28937_ (_24388_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _28938_ (_27273_, _24388_, _24387_);
  and _28939_ (_24389_, _24373_, _24089_);
  and _28940_ (_24391_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _28941_ (_27272_, _24391_, _24389_);
  and _28942_ (_24392_, _24373_, _23583_);
  and _28943_ (_24393_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _28944_ (_27271_, _24393_, _24392_);
  and _28945_ (_24394_, _24146_, _22982_);
  and _28946_ (_24395_, _24394_, _24089_);
  not _28947_ (_24396_, _24394_);
  and _28948_ (_24397_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _28949_ (_27264_, _24397_, _24395_);
  and _28950_ (_24398_, _24381_, _24134_);
  and _28951_ (_24399_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _28952_ (_27046_, _24399_, _24398_);
  and _28953_ (_24400_, _24394_, _23583_);
  and _28954_ (_24401_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _28955_ (_27263_, _24401_, _24400_);
  and _28956_ (_24402_, _24381_, _24051_);
  and _28957_ (_24403_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _28958_ (_27045_, _24403_, _24402_);
  and _28959_ (_24404_, _24394_, _23996_);
  and _28960_ (_24405_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _28961_ (_27267_, _24405_, _24404_);
  and _28962_ (_24406_, _24394_, _24134_);
  and _28963_ (_24407_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _28964_ (_27266_, _24407_, _24406_);
  and _28965_ (_24408_, _24097_, _24004_);
  and _28966_ (_24409_, _24408_, _24319_);
  and _28967_ (_24410_, _24409_, _24219_);
  not _28968_ (_24411_, _24409_);
  and _28969_ (_24412_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or _28970_ (_27118_, _24412_, _24410_);
  and _28971_ (_24413_, _24394_, _24051_);
  and _28972_ (_24414_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _28973_ (_27265_, _24414_, _24413_);
  and _28974_ (_24415_, _23945_, _22974_);
  and _28975_ (_24416_, _24415_, _24134_);
  not _28976_ (_24417_, _24415_);
  and _28977_ (_24418_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or _28978_ (_27041_, _24418_, _24416_);
  and _28979_ (_24420_, _24415_, _24051_);
  and _28980_ (_24421_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or _28981_ (_27040_, _24421_, _24420_);
  or _28982_ (_24422_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _28983_ (_24424_, _24422_, _22731_);
  nand _28984_ (_24425_, _24189_, _23989_);
  and _28985_ (_02924_, _24425_, _24424_);
  and _28986_ (_24426_, _24155_, _23548_);
  and _28987_ (_24428_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or _28988_ (_27275_, _24428_, _24426_);
  and _28989_ (_24430_, _24219_, _24155_);
  and _28990_ (_24431_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or _28991_ (_27274_, _24431_, _24430_);
  and _28992_ (_24433_, _24350_, _23583_);
  and _28993_ (_24434_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _28994_ (_27059_, _24434_, _24433_);
  and _28995_ (_03359_, t1_i, _22731_);
  and _28996_ (_24436_, _24381_, _24219_);
  and _28997_ (_24437_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _28998_ (_27042_, _24437_, _24436_);
  and _28999_ (_24438_, _24155_, _23583_);
  and _29000_ (_24439_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or _29001_ (_27277_, _24439_, _24438_);
  and _29002_ (_24440_, _24155_, _23887_);
  and _29003_ (_24441_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or _29004_ (_27276_, _24441_, _24440_);
  and _29005_ (_24442_, _24146_, _24006_);
  and _29006_ (_24443_, _24442_, _23887_);
  not _29007_ (_24444_, _24442_);
  and _29008_ (_24446_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or _29009_ (_27074_, _24446_, _24443_);
  and _29010_ (_24447_, _24302_, _23996_);
  and _29011_ (_24448_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or _29012_ (_04393_, _24448_, _24447_);
  and _29013_ (_24449_, _24415_, _24219_);
  and _29014_ (_24450_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or _29015_ (_27039_, _24450_, _24449_);
  and _29016_ (_24451_, _24301_, _24146_);
  and _29017_ (_24452_, _24451_, _24134_);
  not _29018_ (_24453_, _24451_);
  and _29019_ (_24454_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _29020_ (_04780_, _24454_, _24452_);
  nor _29021_ (_24455_, _22737_, _23183_);
  and _29022_ (_24457_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _29023_ (_24458_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _29024_ (_24459_, _24458_, _24457_);
  and _29025_ (_24460_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _29026_ (_24461_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _29027_ (_24462_, _24461_, _24460_);
  and _29028_ (_24464_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _29029_ (_24465_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _29030_ (_24467_, _24465_, _24464_);
  and _29031_ (_24468_, _24467_, _24462_);
  and _29032_ (_24469_, _24468_, _24459_);
  and _29033_ (_24470_, _22737_, _23623_);
  not _29034_ (_24471_, _24470_);
  nor _29035_ (_24472_, _24471_, _24469_);
  nor _29036_ (_24473_, _24472_, _24455_);
  nor _29037_ (_26867_[3], _24473_, rst);
  and _29038_ (_24474_, _23940_, _22923_);
  and _29039_ (_24476_, _24300_, _22977_);
  and _29040_ (_24478_, _24476_, _24474_);
  and _29041_ (_24479_, _24478_, _23548_);
  not _29042_ (_24480_, _24478_);
  and _29043_ (_24481_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _29044_ (_27171_, _24481_, _24479_);
  and _29045_ (_24482_, _24478_, _24219_);
  and _29046_ (_24484_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _29047_ (_04945_, _24484_, _24482_);
  and _29048_ (_24485_, _24095_, _23945_);
  and _29049_ (_24486_, _24485_, _23996_);
  not _29050_ (_24487_, _24485_);
  and _29051_ (_24489_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or _29052_ (_05303_, _24489_, _24486_);
  and _29053_ (_24490_, _24365_, _24095_);
  and _29054_ (_24491_, _24490_, _24134_);
  not _29055_ (_24492_, _24490_);
  and _29056_ (_24493_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _29057_ (_05608_, _24493_, _24491_);
  and _29058_ (_24494_, _24409_, _23887_);
  and _29059_ (_24495_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or _29060_ (_05764_, _24495_, _24494_);
  and _29061_ (_24496_, _24003_, _22981_);
  and _29062_ (_24497_, _24496_, _24474_);
  and _29063_ (_24499_, _24497_, _23548_);
  not _29064_ (_24500_, _24497_);
  and _29065_ (_24502_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or _29066_ (_05861_, _24502_, _24499_);
  and _29067_ (_24503_, _24365_, _22974_);
  and _29068_ (_24504_, _24503_, _23548_);
  not _29069_ (_24505_, _24503_);
  and _29070_ (_24507_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _29071_ (_05882_, _24507_, _24504_);
  and _29072_ (_24508_, _24503_, _23887_);
  and _29073_ (_24509_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _29074_ (_05940_, _24509_, _24508_);
  and _29075_ (_24510_, _24365_, _24140_);
  and _29076_ (_24511_, _24510_, _24089_);
  not _29077_ (_24512_, _24510_);
  and _29078_ (_24513_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _29079_ (_06025_, _24513_, _24511_);
  and _29080_ (_24514_, _24415_, _23887_);
  and _29081_ (_24515_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or _29082_ (_06056_, _24515_, _24514_);
  and _29083_ (_24516_, _24510_, _24051_);
  and _29084_ (_24517_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _29085_ (_06076_, _24517_, _24516_);
  and _29086_ (_24518_, _24301_, _24056_);
  and _29087_ (_24519_, _24518_, _23548_);
  not _29088_ (_24520_, _24518_);
  and _29089_ (_24521_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or _29090_ (_27219_, _24521_, _24519_);
  and _29091_ (_24522_, _24510_, _23996_);
  and _29092_ (_24523_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _29093_ (_06235_, _24523_, _24522_);
  and _29094_ (_24525_, _24365_, _24146_);
  and _29095_ (_24526_, _24525_, _24219_);
  not _29096_ (_24527_, _24525_);
  and _29097_ (_24528_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or _29098_ (_06304_, _24528_, _24526_);
  and _29099_ (_24529_, _24525_, _23583_);
  and _29100_ (_24530_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or _29101_ (_06382_, _24530_, _24529_);
  not _29102_ (_24531_, _23504_);
  nor _29103_ (_24532_, _22919_, _22886_);
  and _29104_ (_24533_, _24532_, _22951_);
  and _29105_ (_24534_, _24533_, _24531_);
  nand _29106_ (_24535_, _22951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor _29107_ (_24536_, _24535_, _24532_);
  or _29108_ (_24537_, _24536_, _24534_);
  and _29109_ (_24538_, _22968_, _22937_);
  and _29110_ (_24539_, _24178_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not _29111_ (_24540_, _24539_);
  nor _29112_ (_24541_, _24540_, _22867_);
  and _29113_ (_24542_, _24541_, _22906_);
  and _29114_ (_24543_, _24542_, _22844_);
  and _29115_ (_24544_, _24543_, _24538_);
  and _29116_ (_24545_, _24544_, _24537_);
  nand _29117_ (_24546_, _24544_, _22951_);
  and _29118_ (_24547_, _24546_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor _29119_ (_24548_, _22936_, _22905_);
  and _29120_ (_24549_, _24548_, _23944_);
  not _29121_ (_24550_, _22951_);
  and _29122_ (_24551_, _24550_, _22867_);
  and _29123_ (_24552_, _24532_, _24179_);
  and _29124_ (_24553_, _24552_, _24551_);
  and _29125_ (_24554_, _24553_, _24549_);
  or _29126_ (_24555_, _24554_, _24547_);
  or _29127_ (_24556_, _24555_, _24545_);
  not _29128_ (_24557_, _24554_);
  or _29129_ (_24558_, _24557_, _23577_);
  and _29130_ (_24559_, _24558_, _22731_);
  and _29131_ (_06442_, _24559_, _24556_);
  not _29132_ (_24560_, _22919_);
  and _29133_ (_24561_, _24560_, _22886_);
  and _29134_ (_24562_, _24561_, _22951_);
  and _29135_ (_24563_, _24544_, _24562_);
  or _29136_ (_24564_, _24563_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _29137_ (_24565_, _24564_, _24557_);
  nand _29138_ (_24566_, _24563_, _23504_);
  and _29139_ (_24567_, _24566_, _24565_);
  and _29140_ (_24568_, _24554_, _23880_);
  or _29141_ (_24569_, _24568_, _24567_);
  and _29142_ (_06510_, _24569_, _22731_);
  and _29143_ (_24570_, _24544_, _24177_);
  and _29144_ (_24571_, _24570_, _23504_);
  nor _29145_ (_24572_, _24570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _29146_ (_24573_, _24572_, _24571_);
  nand _29147_ (_24574_, _24573_, _24557_);
  nand _29148_ (_24575_, _24554_, _23542_);
  and _29149_ (_24576_, _24575_, _22731_);
  and _29150_ (_06536_, _24576_, _24574_);
  and _29151_ (_24577_, _24176_, _22886_);
  and _29152_ (_24578_, _24544_, _24577_);
  and _29153_ (_24579_, _24578_, _23504_);
  nor _29154_ (_24580_, _24578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _29155_ (_24581_, _24580_, _24579_);
  nand _29156_ (_24582_, _24581_, _24557_);
  nand _29157_ (_24583_, _24554_, _24210_);
  and _29158_ (_24584_, _24583_, _22731_);
  and _29159_ (_06560_, _24584_, _24582_);
  and _29160_ (_24585_, _24415_, _23583_);
  and _29161_ (_24586_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or _29162_ (_06601_, _24586_, _24585_);
  and _29163_ (_24587_, _24525_, _24089_);
  and _29164_ (_24588_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or _29165_ (_06622_, _24588_, _24587_);
  and _29166_ (_24589_, _24525_, _24134_);
  and _29167_ (_24590_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or _29168_ (_27194_, _24590_, _24589_);
  and _29169_ (_24591_, _24525_, _23996_);
  and _29170_ (_24592_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or _29171_ (_06722_, _24592_, _24591_);
  nor _29172_ (_24593_, _22951_, _22919_);
  and _29173_ (_24594_, _24593_, _22886_);
  and _29174_ (_24595_, _24594_, _24544_);
  and _29175_ (_24596_, _24595_, _23504_);
  nor _29176_ (_24597_, _24595_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _29177_ (_24598_, _24597_, _24596_);
  nand _29178_ (_24599_, _24598_, _24557_);
  nand _29179_ (_24600_, _24554_, _24126_);
  and _29180_ (_24601_, _24600_, _22731_);
  and _29181_ (_06752_, _24601_, _24599_);
  and _29182_ (_24602_, _24372_, _24365_);
  and _29183_ (_24603_, _24602_, _23548_);
  not _29184_ (_24604_, _24602_);
  and _29185_ (_24605_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or _29186_ (_06772_, _24605_, _24603_);
  and _29187_ (_24606_, _22919_, _24175_);
  and _29188_ (_24607_, _24606_, _24550_);
  and _29189_ (_24608_, _24607_, _24544_);
  nand _29190_ (_24609_, _24608_, _23504_);
  or _29191_ (_24610_, _24608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _29192_ (_24611_, _24610_, _24557_);
  and _29193_ (_24612_, _24611_, _24609_);
  nor _29194_ (_24613_, _24557_, _24043_);
  or _29195_ (_24614_, _24613_, _24612_);
  and _29196_ (_06793_, _24614_, _22731_);
  and _29197_ (_24615_, _24602_, _23583_);
  and _29198_ (_24616_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or _29199_ (_06814_, _24616_, _24615_);
  and _29200_ (_24617_, _24602_, _24051_);
  and _29201_ (_24618_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or _29202_ (_06894_, _24618_, _24617_);
  and _29203_ (_24619_, _24541_, _22905_);
  and _29204_ (_24620_, _24619_, _22844_);
  and _29205_ (_24621_, _24620_, _24538_);
  and _29206_ (_24622_, _24621_, _24177_);
  nand _29207_ (_24623_, _24622_, _23504_);
  or _29208_ (_24624_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _29209_ (_24625_, _22937_, _22905_);
  and _29210_ (_24626_, _24625_, _23944_);
  and _29211_ (_24627_, _24577_, _22868_);
  and _29212_ (_24628_, _24627_, _24179_);
  and _29213_ (_24629_, _24628_, _24626_);
  not _29214_ (_24630_, _24629_);
  and _29215_ (_24631_, _24630_, _24624_);
  and _29216_ (_24632_, _24631_, _24623_);
  nor _29217_ (_24633_, _24630_, _23542_);
  or _29218_ (_24634_, _24633_, _24632_);
  and _29219_ (_06967_, _24634_, _22731_);
  and _29220_ (_24635_, _22919_, _22886_);
  and _29221_ (_24636_, _24635_, _24550_);
  and _29222_ (_24637_, _24636_, _24531_);
  nor _29223_ (_24638_, _24635_, _24550_);
  and _29224_ (_24639_, _24638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _29225_ (_24640_, _24639_, _24637_);
  and _29226_ (_24641_, _24640_, _24621_);
  not _29227_ (_24642_, _24621_);
  nor _29228_ (_24643_, _24638_, _24636_);
  or _29229_ (_24644_, _24643_, _24642_);
  and _29230_ (_24645_, _24644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _29231_ (_24646_, _24645_, _24629_);
  or _29232_ (_24647_, _24646_, _24641_);
  nand _29233_ (_24648_, _24629_, _24082_);
  and _29234_ (_24649_, _24648_, _22731_);
  and _29235_ (_07024_, _24649_, _24647_);
  and _29236_ (_24650_, _24602_, _24134_);
  and _29237_ (_24651_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or _29238_ (_07047_, _24651_, _24650_);
  and _29239_ (_24652_, _24621_, _24533_);
  nand _29240_ (_24653_, _24652_, _23504_);
  or _29241_ (_24654_, _24652_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _29242_ (_24655_, _24654_, _24630_);
  and _29243_ (_24656_, _24655_, _24653_);
  and _29244_ (_24657_, _24629_, _23577_);
  or _29245_ (_24658_, _24657_, _24656_);
  and _29246_ (_07072_, _24658_, _22731_);
  and _29247_ (_24659_, _24621_, _24562_);
  nand _29248_ (_24660_, _24659_, _23504_);
  or _29249_ (_24661_, _24659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _29250_ (_24662_, _24661_, _24630_);
  and _29251_ (_24663_, _24662_, _24660_);
  and _29252_ (_24664_, _24629_, _23880_);
  or _29253_ (_24665_, _24664_, _24663_);
  and _29254_ (_07135_, _24665_, _22731_);
  and _29255_ (_24666_, _24621_, _24577_);
  nand _29256_ (_24667_, _24666_, _23504_);
  or _29257_ (_24668_, _24666_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _29258_ (_24669_, _24668_, _24630_);
  and _29259_ (_24670_, _24669_, _24667_);
  not _29260_ (_24671_, _24210_);
  and _29261_ (_24672_, _24629_, _24671_);
  or _29262_ (_24673_, _24672_, _24670_);
  and _29263_ (_07156_, _24673_, _22731_);
  and _29264_ (_24674_, _24490_, _24219_);
  and _29265_ (_24675_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _29266_ (_07199_, _24675_, _24674_);
  and _29267_ (_24676_, _24490_, _23887_);
  and _29268_ (_24677_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _29269_ (_07223_, _24677_, _24676_);
  and _29270_ (_24678_, _24490_, _24089_);
  and _29271_ (_24679_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _29272_ (_07276_, _24679_, _24678_);
  and _29273_ (_24680_, _24490_, _24051_);
  and _29274_ (_24681_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _29275_ (_07366_, _24681_, _24680_);
  and _29276_ (_24682_, _24503_, _24051_);
  and _29277_ (_24684_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _29278_ (_07386_, _24684_, _24682_);
  and _29279_ (_24685_, _24621_, _24594_);
  nand _29280_ (_24686_, _24685_, _23504_);
  or _29281_ (_24687_, _24685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _29282_ (_24688_, _24687_, _24630_);
  and _29283_ (_24689_, _24688_, _24686_);
  nor _29284_ (_24690_, _24630_, _24126_);
  or _29285_ (_24691_, _24690_, _24689_);
  and _29286_ (_07479_, _24691_, _22731_);
  and _29287_ (_24692_, _24503_, _24134_);
  and _29288_ (_24693_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _29289_ (_07614_, _24693_, _24692_);
  and _29290_ (_24694_, _24365_, _24319_);
  and _29291_ (_24695_, _24694_, _24219_);
  not _29292_ (_24696_, _24694_);
  and _29293_ (_24697_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or _29294_ (_07645_, _24697_, _24695_);
  and _29295_ (_24698_, _22968_, _22936_);
  and _29296_ (_24699_, _24698_, _24620_);
  and _29297_ (_24700_, _24699_, _24636_);
  nand _29298_ (_24701_, _24700_, _23504_);
  or _29299_ (_24702_, _24700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _29300_ (_24703_, _24628_, _24174_);
  not _29301_ (_24704_, _24703_);
  and _29302_ (_24705_, _24704_, _24702_);
  and _29303_ (_24706_, _24705_, _24701_);
  nor _29304_ (_24707_, _24704_, _24082_);
  or _29305_ (_24708_, _24707_, _24706_);
  and _29306_ (_07703_, _24708_, _22731_);
  and _29307_ (_24709_, _24699_, _24562_);
  nand _29308_ (_24710_, _24709_, _23504_);
  or _29309_ (_24711_, _24709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _29310_ (_24712_, _24711_, _24704_);
  and _29311_ (_24713_, _24712_, _24710_);
  and _29312_ (_24714_, _24703_, _23880_);
  or _29313_ (_24715_, _24714_, _24713_);
  and _29314_ (_07723_, _24715_, _22731_);
  and _29315_ (_24716_, _24699_, _24577_);
  or _29316_ (_24717_, _24716_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _29317_ (_24718_, _24717_, _24704_);
  nand _29318_ (_24719_, _24716_, _23504_);
  and _29319_ (_24720_, _24719_, _24718_);
  and _29320_ (_24721_, _24703_, _24671_);
  or _29321_ (_24722_, _24721_, _24720_);
  and _29322_ (_07742_, _24722_, _22731_);
  and _29323_ (_24723_, _24694_, _23548_);
  and _29324_ (_24724_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or _29325_ (_07762_, _24724_, _24723_);
  and _29326_ (_24725_, _24694_, _24089_);
  and _29327_ (_24726_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or _29328_ (_07812_, _24726_, _24725_);
  and _29329_ (_24727_, _24485_, _24219_);
  and _29330_ (_24728_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or _29331_ (_07894_, _24728_, _24727_);
  and _29332_ (_24729_, _24694_, _24051_);
  and _29333_ (_24730_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or _29334_ (_07923_, _24730_, _24729_);
  and _29335_ (_24731_, _24694_, _23996_);
  and _29336_ (_24732_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or _29337_ (_07944_, _24732_, _24731_);
  and _29338_ (_24733_, _24302_, _24134_);
  and _29339_ (_24734_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or _29340_ (_08017_, _24734_, _24733_);
  and _29341_ (_24735_, _24365_, _24223_);
  and _29342_ (_24736_, _24735_, _24219_);
  not _29343_ (_24737_, _24735_);
  and _29344_ (_24738_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or _29345_ (_08087_, _24738_, _24736_);
  and _29346_ (_24739_, _24485_, _23887_);
  and _29347_ (_24740_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or _29348_ (_08103_, _24740_, _24739_);
  and _29349_ (_24741_, _24735_, _23583_);
  and _29350_ (_24742_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or _29351_ (_08123_, _24742_, _24741_);
  and _29352_ (_24743_, _24735_, _24051_);
  and _29353_ (_24744_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or _29354_ (_08142_, _24744_, _24743_);
  and _29355_ (_24745_, _24735_, _23996_);
  and _29356_ (_24746_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or _29357_ (_08169_, _24746_, _24745_);
  and _29358_ (_24747_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _29359_ (_24748_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _29360_ (_24749_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _29361_ (_24750_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _29362_ (_24751_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _24750_);
  and _29363_ (_24752_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29364_ (_24753_, _24752_, _24751_);
  and _29365_ (_24754_, _24753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _29366_ (_24755_, _24754_, _24749_);
  and _29367_ (_24756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _29368_ (_24757_, _24756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _29369_ (_24758_, _24757_);
  and _29370_ (_24759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _29371_ (_24760_, _24759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29372_ (_24761_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _29373_ (_24762_, _24761_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _29374_ (_24763_, _24762_, _24760_);
  and _29375_ (_24764_, _24763_, _24758_);
  nor _29376_ (_24765_, _24764_, _24755_);
  not _29377_ (_24766_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _29378_ (_24767_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _29379_ (_24768_, _24767_, _24766_);
  nand _29380_ (_24769_, _24768_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _29381_ (_24770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _29382_ (_24771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _29383_ (_24772_, _24771_, _24770_);
  and _29384_ (_24773_, _24772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _29385_ (_24774_, _24773_);
  and _29386_ (_24775_, _24774_, _24769_);
  and _29387_ (_24776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _29388_ (_24777_, _24776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _29389_ (_24778_, _24777_);
  and _29390_ (_24779_, _24778_, _24775_);
  nor _29391_ (_24780_, _24779_, _24755_);
  nor _29392_ (_24781_, _24780_, _24765_);
  and _29393_ (_24782_, _24749_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not _29394_ (_24783_, _24782_);
  not _29395_ (_24784_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _29396_ (_24785_, _24768_, _24784_);
  not _29397_ (_24786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _29398_ (_24787_, _24772_, _24786_);
  nor _29399_ (_24788_, _24787_, _24785_);
  not _29400_ (_24789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _29401_ (_24790_, _24776_, _24789_);
  not _29402_ (_24791_, _24790_);
  and _29403_ (_24792_, _24791_, _24788_);
  nor _29404_ (_24793_, _24792_, _24783_);
  not _29405_ (_24794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _29406_ (_24795_, _24756_, _24794_);
  not _29407_ (_24797_, _24795_);
  not _29408_ (_24798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29409_ (_24799_, _24759_, _24798_);
  not _29410_ (_24800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _29411_ (_24801_, _24761_, _24800_);
  nor _29412_ (_24802_, _24801_, _24799_);
  and _29413_ (_24803_, _24802_, _24797_);
  nor _29414_ (_24804_, _24803_, _24783_);
  nor _29415_ (_24805_, _24804_, _24793_);
  not _29416_ (_24806_, _24805_);
  and _29417_ (_24807_, _24806_, _24781_);
  nand _29418_ (_24808_, _24807_, _24748_);
  not _29419_ (_24809_, _24781_);
  and _29420_ (_24810_, _24809_, _24748_);
  or _29421_ (_24811_, _24810_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _29422_ (_24812_, _24811_, _22731_);
  and _29423_ (_08233_, _24812_, _24808_);
  and _29424_ (_24813_, _24365_, _24056_);
  and _29425_ (_24814_, _24813_, _24219_);
  not _29426_ (_24815_, _24813_);
  and _29427_ (_24816_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _29428_ (_08294_, _24816_, _24814_);
  and _29429_ (_24817_, _24485_, _23548_);
  and _29430_ (_24818_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or _29431_ (_08331_, _24818_, _24817_);
  and _29432_ (_24819_, _24813_, _23887_);
  and _29433_ (_24820_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _29434_ (_08378_, _24820_, _24819_);
  and _29435_ (_24821_, _24813_, _24089_);
  and _29436_ (_24822_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _29437_ (_08397_, _24822_, _24821_);
  and _29438_ (_26840_[6], _23745_, _22731_);
  and _29439_ (_24823_, _24813_, _24134_);
  and _29440_ (_24824_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _29441_ (_08490_, _24824_, _24823_);
  and _29442_ (_24825_, _24813_, _23996_);
  and _29443_ (_24826_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _29444_ (_27196_, _24826_, _24825_);
  nor _29445_ (_24827_, _24747_, _24750_);
  nand _29446_ (_24828_, _24827_, _24807_);
  and _29447_ (_24829_, _24827_, _24809_);
  or _29448_ (_24830_, _24829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _29449_ (_24831_, _24830_, _22731_);
  and _29450_ (_08572_, _24831_, _24828_);
  and _29451_ (_24832_, _24474_, _24365_);
  and _29452_ (_24833_, _24832_, _23887_);
  not _29453_ (_24834_, _24832_);
  and _29454_ (_24835_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or _29455_ (_08606_, _24835_, _24833_);
  and _29456_ (_24836_, _24832_, _24089_);
  and _29457_ (_24837_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or _29458_ (_27198_, _24837_, _24836_);
  and _29459_ (_24838_, _24832_, _24134_);
  and _29460_ (_24839_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or _29461_ (_08724_, _24839_, _24838_);
  and _29462_ (_24840_, _24805_, _24781_);
  nor _29463_ (_24841_, _24840_, _24747_);
  not _29464_ (_24842_, _24841_);
  and _29465_ (_24843_, _24842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _29466_ (_24844_, _24747_);
  nor _29467_ (_24845_, _24769_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29468_ (_24846_, _24845_, _24777_);
  not _29469_ (_24847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _29470_ (_24848_, _24773_, _24750_);
  or _29471_ (_24849_, _24848_, _24847_);
  nand _29472_ (_24850_, _24849_, _24846_);
  and _29473_ (_24851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29474_ (_24852_, _24851_, _24778_);
  and _29475_ (_24853_, _24852_, _24850_);
  or _29476_ (_24854_, _24853_, _24762_);
  not _29477_ (_24855_, _24760_);
  not _29478_ (_24856_, _24762_);
  or _29479_ (_24857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _24750_);
  or _29480_ (_24858_, _24857_, _24856_);
  and _29481_ (_24859_, _24858_, _24855_);
  and _29482_ (_24860_, _24859_, _24854_);
  and _29483_ (_24861_, _24851_, _24760_);
  or _29484_ (_24862_, _24861_, _24757_);
  or _29485_ (_24863_, _24862_, _24860_);
  nor _29486_ (_24864_, _24857_, _24758_);
  nor _29487_ (_24865_, _24864_, _24781_);
  and _29488_ (_24866_, _24865_, _24863_);
  or _29489_ (_24867_, _24857_, _24797_);
  and _29490_ (_24868_, _24785_, _24750_);
  nor _29491_ (_24869_, _24868_, _24790_);
  and _29492_ (_24870_, _24787_, _24750_);
  or _29493_ (_24871_, _24870_, _24847_);
  nand _29494_ (_24872_, _24871_, _24869_);
  or _29495_ (_24873_, _24851_, _24791_);
  and _29496_ (_24874_, _24873_, _24872_);
  or _29497_ (_24875_, _24874_, _24801_);
  not _29498_ (_24876_, _24799_);
  not _29499_ (_24877_, _24801_);
  or _29500_ (_24878_, _24857_, _24877_);
  and _29501_ (_24879_, _24878_, _24876_);
  and _29502_ (_24880_, _24879_, _24875_);
  and _29503_ (_24881_, _24851_, _24799_);
  or _29504_ (_24882_, _24881_, _24795_);
  or _29505_ (_24883_, _24882_, _24880_);
  and _29506_ (_24884_, _24883_, _24807_);
  and _29507_ (_24885_, _24884_, _24867_);
  or _29508_ (_24886_, _24885_, _24866_);
  and _29509_ (_24887_, _24886_, _24844_);
  or _29510_ (_24888_, _24887_, _24843_);
  and _29511_ (_08746_, _24888_, _22731_);
  and _29512_ (_24889_, _24006_, _22974_);
  and _29513_ (_24890_, _24889_, _24219_);
  not _29514_ (_24891_, _24889_);
  and _29515_ (_24892_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or _29516_ (_08767_, _24892_, _24890_);
  nand _29517_ (_24893_, _24840_, _24748_);
  and _29518_ (_24894_, _24781_, _24844_);
  or _29519_ (_24895_, _24894_, _24750_);
  and _29520_ (_24896_, _24895_, _22731_);
  and _29521_ (_08845_, _24896_, _24893_);
  and _29522_ (_24897_, _24832_, _23996_);
  and _29523_ (_24898_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or _29524_ (_08971_, _24898_, _24897_);
  and _29525_ (_24899_, _24014_, _23940_);
  and _29526_ (_24900_, _24899_, _24365_);
  and _29527_ (_24902_, _24900_, _23548_);
  not _29528_ (_24903_, _24900_);
  and _29529_ (_24904_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _29530_ (_09008_, _24904_, _24902_);
  and _29531_ (_24905_, _24900_, _23583_);
  and _29532_ (_24906_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _29533_ (_09032_, _24906_, _24905_);
  and _29534_ (_24907_, _24900_, _24051_);
  and _29535_ (_24908_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _29536_ (_09093_, _24908_, _24907_);
  not _29537_ (_24909_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor _29538_ (_24910_, _24841_, _24909_);
  or _29539_ (_24911_, _24778_, _24762_);
  and _29540_ (_24912_, _24911_, _24855_);
  and _29541_ (_24913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _24750_);
  or _29542_ (_24914_, _24913_, _24912_);
  and _29543_ (_24915_, _24773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29544_ (_24916_, _24915_, _24909_);
  nor _29545_ (_24917_, _24769_, _24750_);
  nor _29546_ (_24918_, _24917_, _24777_);
  nand _29547_ (_24919_, _24918_, _24763_);
  or _29548_ (_24920_, _24919_, _24916_);
  and _29549_ (_24921_, _24920_, _24914_);
  or _29550_ (_24922_, _24921_, _24757_);
  or _29551_ (_24923_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29552_ (_24924_, _24856_, _24760_);
  and _29553_ (_24925_, _24924_, _24758_);
  nor _29554_ (_24926_, _24925_, _24923_);
  nor _29555_ (_24927_, _24926_, _24781_);
  and _29556_ (_24928_, _24927_, _24922_);
  and _29557_ (_24929_, _24785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29558_ (_24930_, _24929_, _24790_);
  and _29559_ (_24931_, _24787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29560_ (_24932_, _24931_, _24909_);
  nand _29561_ (_24933_, _24932_, _24930_);
  or _29562_ (_24934_, _24913_, _24791_);
  and _29563_ (_24935_, _24934_, _24933_);
  or _29564_ (_24936_, _24935_, _24801_);
  or _29565_ (_24937_, _24923_, _24877_);
  and _29566_ (_24938_, _24937_, _24876_);
  and _29567_ (_24939_, _24938_, _24936_);
  and _29568_ (_24940_, _24913_, _24799_);
  or _29569_ (_24941_, _24940_, _24795_);
  or _29570_ (_24942_, _24941_, _24939_);
  and _29571_ (_24943_, _24807_, _24797_);
  and _29572_ (_24944_, _24923_, _24807_);
  or _29573_ (_24945_, _24944_, _24943_);
  and _29574_ (_24946_, _24945_, _24942_);
  or _29575_ (_24947_, _24946_, _24928_);
  and _29576_ (_24948_, _24947_, _24844_);
  or _29577_ (_24949_, _24948_, _24910_);
  and _29578_ (_09118_, _24949_, _22731_);
  and _29579_ (_24950_, _24900_, _24134_);
  and _29580_ (_24951_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _29581_ (_27200_, _24951_, _24950_);
  and _29582_ (_24952_, _24365_, _23941_);
  and _29583_ (_24953_, _24952_, _23548_);
  not _29584_ (_24954_, _24952_);
  and _29585_ (_24955_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _29586_ (_27201_, _24955_, _24953_);
  and _29587_ (_24956_, _24952_, _23887_);
  and _29588_ (_24957_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _29589_ (_09448_, _24957_, _24956_);
  and _29590_ (_24959_, _24952_, _24089_);
  and _29591_ (_24960_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _29592_ (_09479_, _24960_, _24959_);
  and _29593_ (_24961_, _24952_, _24134_);
  and _29594_ (_24962_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _29595_ (_09499_, _24962_, _24961_);
  and _29596_ (_24963_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _29597_ (_24964_, _24963_, _24841_);
  and _29598_ (_09539_, _24964_, _22731_);
  or _29599_ (_24965_, _24801_, _24790_);
  nor _29600_ (_24966_, _24799_, _24795_);
  nand _29601_ (_24967_, _24966_, _24782_);
  or _29602_ (_24968_, _24967_, _24965_);
  nor _29603_ (_24969_, _24968_, _24788_);
  and _29604_ (_24970_, _24969_, _24781_);
  and _29605_ (_24971_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor _29606_ (_24972_, _24777_, _24755_);
  not _29607_ (_24973_, _24764_);
  nor _29608_ (_24974_, _24775_, _24973_);
  and _29609_ (_24975_, _24974_, _24972_);
  and _29610_ (_24976_, _24975_, _24844_);
  or _29611_ (_24977_, _24976_, _24971_);
  or _29612_ (_24978_, _24977_, _24970_);
  and _29613_ (_09560_, _24978_, _22731_);
  and _29614_ (_24979_, _24788_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _29615_ (_24980_, _24979_, _24965_);
  and _29616_ (_24981_, _24980_, _24966_);
  and _29617_ (_24982_, _24981_, _24807_);
  nor _29618_ (_24983_, _24760_, _24757_);
  or _29619_ (_24984_, _24777_, _24762_);
  and _29620_ (_24985_, _24775_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _29621_ (_24986_, _24985_, _24984_);
  nand _29622_ (_24987_, _24986_, _24983_);
  nor _29623_ (_24988_, _24987_, _24781_);
  or _29624_ (_24989_, _24988_, _24747_);
  or _29625_ (_24990_, _24989_, _24982_);
  or _29626_ (_24991_, _24844_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _29627_ (_24992_, _24991_, _22731_);
  and _29628_ (_09580_, _24992_, _24990_);
  and _29629_ (_24993_, _24367_, _24219_);
  and _29630_ (_24994_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or _29631_ (_09600_, _24994_, _24993_);
  nor _29632_ (_24995_, _24787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _29633_ (_24996_, _24995_, _24785_);
  or _29634_ (_24997_, _24996_, _24790_);
  and _29635_ (_24998_, _24997_, _24877_);
  or _29636_ (_24999_, _24998_, _24799_);
  and _29637_ (_25000_, _24999_, _24943_);
  or _29638_ (_25001_, _24773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _29639_ (_25002_, _25001_, _24769_);
  or _29640_ (_25003_, _25002_, _24777_);
  and _29641_ (_25004_, _25003_, _24856_);
  or _29642_ (_25005_, _25004_, _24760_);
  nor _29643_ (_25006_, _24781_, _24757_);
  and _29644_ (_25007_, _25006_, _25005_);
  or _29645_ (_25008_, _25007_, _24747_);
  or _29646_ (_25009_, _25008_, _25000_);
  not _29647_ (_25010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nand _29648_ (_25011_, _24747_, _25010_);
  and _29649_ (_25012_, _25011_, _22731_);
  and _29650_ (_09621_, _25012_, _25009_);
  and _29651_ (_25013_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _22731_);
  and _29652_ (_09650_, _25013_, _24747_);
  and _29653_ (_25014_, _24367_, _23548_);
  and _29654_ (_25015_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or _29655_ (_09745_, _25015_, _25014_);
  and _29656_ (_25016_, _22906_, _22867_);
  and _29657_ (_25017_, _25016_, _22844_);
  and _29658_ (_25018_, _25017_, _24538_);
  and _29659_ (_25019_, _25018_, _24533_);
  nand _29660_ (_25020_, _25019_, _23504_);
  or _29661_ (_25021_, _25019_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _29662_ (_25022_, _25021_, _24539_);
  and _29663_ (_25023_, _25022_, _25020_);
  and _29664_ (_25024_, _24577_, _22867_);
  and _29665_ (_25025_, _25024_, _24548_);
  and _29666_ (_25026_, _25025_, _23944_);
  not _29667_ (_25027_, _25026_);
  or _29668_ (_25028_, _25027_, _23577_);
  or _29669_ (_25029_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _29670_ (_25030_, _25029_, _24179_);
  and _29671_ (_25032_, _25030_, _25028_);
  not _29672_ (_25033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor _29673_ (_25034_, _24178_, _25033_);
  or _29674_ (_25035_, _25034_, rst);
  or _29675_ (_25036_, _25035_, _25032_);
  or _29676_ (_09786_, _25036_, _25023_);
  and _29677_ (_25038_, _24367_, _23583_);
  and _29678_ (_25039_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or _29679_ (_09809_, _25039_, _25038_);
  and _29680_ (_25040_, _25018_, _24562_);
  nand _29681_ (_25041_, _25040_, _23504_);
  or _29682_ (_25042_, _25040_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _29683_ (_25043_, _25042_, _24539_);
  and _29684_ (_25044_, _25043_, _25041_);
  or _29685_ (_25045_, _25027_, _23880_);
  or _29686_ (_25046_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _29687_ (_25047_, _25046_, _24179_);
  and _29688_ (_25048_, _25047_, _25045_);
  not _29689_ (_25049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor _29690_ (_25050_, _24178_, _25049_);
  or _29691_ (_25051_, _25050_, rst);
  or _29692_ (_25052_, _25051_, _25048_);
  or _29693_ (_09868_, _25052_, _25044_);
  and _29694_ (_25053_, _25018_, _24177_);
  nand _29695_ (_25054_, _25053_, _23504_);
  or _29696_ (_25055_, _25053_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _29697_ (_25056_, _25055_, _24539_);
  and _29698_ (_25057_, _25056_, _25054_);
  nand _29699_ (_25058_, _25026_, _23542_);
  or _29700_ (_25059_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _29701_ (_25060_, _25059_, _24179_);
  and _29702_ (_25061_, _25060_, _25058_);
  not _29703_ (_25062_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor _29704_ (_25063_, _24178_, _25062_);
  or _29705_ (_25064_, _25063_, rst);
  or _29706_ (_25065_, _25064_, _25061_);
  or _29707_ (_09894_, _25065_, _25057_);
  and _29708_ (_25066_, _25018_, _24577_);
  nand _29709_ (_25067_, _25066_, _23504_);
  or _29710_ (_25068_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _29711_ (_25069_, _25068_, _24539_);
  and _29712_ (_25070_, _25069_, _25067_);
  nand _29713_ (_25071_, _25026_, _24210_);
  and _29714_ (_25072_, _25071_, _24179_);
  and _29715_ (_25073_, _25072_, _25068_);
  not _29716_ (_25074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _29717_ (_25075_, _24178_, _25074_);
  or _29718_ (_25077_, _25075_, rst);
  or _29719_ (_25078_, _25077_, _25073_);
  or _29720_ (_09922_, _25078_, _25070_);
  and _29721_ (_25080_, _24367_, _24051_);
  and _29722_ (_25081_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or _29723_ (_09986_, _25081_, _25080_);
  and _29724_ (_25083_, _24485_, _24051_);
  and _29725_ (_25084_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or _29726_ (_10012_, _25084_, _25083_);
  and _29727_ (_25085_, _24485_, _24089_);
  and _29728_ (_25086_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or _29729_ (_10107_, _25086_, _25085_);
  and _29730_ (_25088_, _25018_, _24594_);
  nand _29731_ (_25089_, _25088_, _23504_);
  or _29732_ (_25090_, _25088_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _29733_ (_25091_, _25090_, _24539_);
  and _29734_ (_25092_, _25091_, _25089_);
  nand _29735_ (_25093_, _25026_, _24126_);
  or _29736_ (_25094_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _29737_ (_25096_, _25094_, _24179_);
  and _29738_ (_25097_, _25096_, _25093_);
  not _29739_ (_25098_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _29740_ (_25099_, _24178_, _25098_);
  or _29741_ (_25100_, _25099_, rst);
  or _29742_ (_25101_, _25100_, _25097_);
  or _29743_ (_10136_, _25101_, _25092_);
  and _29744_ (_25102_, _24478_, _23583_);
  and _29745_ (_25103_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _29746_ (_10250_, _25103_, _25102_);
  and _29747_ (_25104_, _25018_, _24607_);
  nand _29748_ (_25105_, _25104_, _23504_);
  or _29749_ (_25106_, _25104_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _29750_ (_25107_, _25106_, _24539_);
  and _29751_ (_25108_, _25107_, _25105_);
  nand _29752_ (_25109_, _25026_, _24043_);
  or _29753_ (_25110_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _29754_ (_25111_, _25110_, _24179_);
  and _29755_ (_25112_, _25111_, _25109_);
  not _29756_ (_25113_, _24178_);
  and _29757_ (_25115_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _29758_ (_25116_, _25115_, rst);
  or _29759_ (_25117_, _25116_, _25112_);
  or _29760_ (_10293_, _25117_, _25108_);
  and _29761_ (_25118_, _24485_, _23583_);
  and _29762_ (_25119_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or _29763_ (_10347_, _25119_, _25118_);
  and _29764_ (_25120_, _24478_, _23887_);
  and _29765_ (_25121_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _29766_ (_10382_, _25121_, _25120_);
  and _29767_ (_25122_, _22905_, _22867_);
  and _29768_ (_25123_, _25122_, _22844_);
  and _29769_ (_25124_, _25123_, _24538_);
  and _29770_ (_25125_, _25124_, _24177_);
  nand _29771_ (_25126_, _25125_, _23504_);
  or _29772_ (_25127_, _25125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _29773_ (_25128_, _25127_, _24539_);
  and _29774_ (_25129_, _25128_, _25126_);
  and _29775_ (_25130_, _25024_, _24626_);
  nand _29776_ (_25131_, _25130_, _23542_);
  or _29777_ (_25132_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _29778_ (_25133_, _25132_, _24179_);
  and _29779_ (_25134_, _25133_, _25131_);
  not _29780_ (_25135_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor _29781_ (_25136_, _24178_, _25135_);
  or _29782_ (_25137_, _25136_, rst);
  or _29783_ (_25138_, _25137_, _25134_);
  or _29784_ (_10460_, _25138_, _25129_);
  and _29785_ (_25139_, _25124_, _24607_);
  nand _29786_ (_25140_, _25139_, _23504_);
  or _29787_ (_25141_, _25139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _29788_ (_25142_, _25141_, _24539_);
  and _29789_ (_25143_, _25142_, _25140_);
  nand _29790_ (_25144_, _25130_, _24043_);
  or _29791_ (_25145_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _29792_ (_25146_, _25145_, _24179_);
  and _29793_ (_25147_, _25146_, _25144_);
  and _29794_ (_25148_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _29795_ (_25149_, _25148_, rst);
  or _29796_ (_25150_, _25149_, _25147_);
  or _29797_ (_10482_, _25150_, _25143_);
  and _29798_ (_25151_, _25124_, _24636_);
  nand _29799_ (_25152_, _25151_, _23504_);
  or _29800_ (_25153_, _25151_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _29801_ (_25154_, _25153_, _24539_);
  and _29802_ (_25155_, _25154_, _25152_);
  nand _29803_ (_25156_, _25130_, _24082_);
  or _29804_ (_25157_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _29805_ (_25158_, _25157_, _24179_);
  and _29806_ (_25159_, _25158_, _25156_);
  not _29807_ (_25160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _29808_ (_25161_, _24178_, _25160_);
  or _29809_ (_25162_, _25161_, rst);
  or _29810_ (_25163_, _25162_, _25159_);
  or _29811_ (_10516_, _25163_, _25155_);
  and _29812_ (_25164_, _25124_, _24533_);
  nand _29813_ (_25165_, _25164_, _23504_);
  or _29814_ (_25166_, _25164_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _29815_ (_25167_, _25166_, _24539_);
  and _29816_ (_25168_, _25167_, _25165_);
  not _29817_ (_25169_, _25130_);
  or _29818_ (_25171_, _25169_, _23577_);
  or _29819_ (_25172_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _29820_ (_25173_, _25172_, _24179_);
  and _29821_ (_25174_, _25173_, _25171_);
  not _29822_ (_25175_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor _29823_ (_25176_, _24178_, _25175_);
  or _29824_ (_25177_, _25176_, rst);
  or _29825_ (_25178_, _25177_, _25174_);
  or _29826_ (_10541_, _25178_, _25168_);
  and _29827_ (_25179_, _25124_, _24562_);
  nand _29828_ (_25180_, _25179_, _23504_);
  or _29829_ (_25181_, _25179_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _29830_ (_25182_, _25181_, _24539_);
  and _29831_ (_25183_, _25182_, _25180_);
  or _29832_ (_25184_, _25169_, _23880_);
  or _29833_ (_25185_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _29834_ (_25186_, _25185_, _24179_);
  and _29835_ (_25187_, _25186_, _25184_);
  not _29836_ (_25188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor _29837_ (_25189_, _24178_, _25188_);
  or _29838_ (_25190_, _25189_, rst);
  or _29839_ (_25191_, _25190_, _25187_);
  or _29840_ (_10565_, _25191_, _25183_);
  and _29841_ (_25192_, _25124_, _24577_);
  nand _29842_ (_25193_, _25192_, _23504_);
  or _29843_ (_25194_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _29844_ (_25195_, _25194_, _24539_);
  and _29845_ (_25196_, _25195_, _25193_);
  nand _29846_ (_25197_, _25130_, _24210_);
  and _29847_ (_25198_, _25197_, _24179_);
  and _29848_ (_25199_, _25198_, _25194_);
  not _29849_ (_25200_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _29850_ (_25201_, _24178_, _25200_);
  or _29851_ (_25202_, _25201_, rst);
  or _29852_ (_25203_, _25202_, _25199_);
  or _29853_ (_10592_, _25203_, _25196_);
  and _29854_ (_25204_, _24237_, _23996_);
  and _29855_ (_25205_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _29856_ (_27065_, _25205_, _25204_);
  and _29857_ (_25206_, _24372_, _23945_);
  and _29858_ (_25207_, _25206_, _24089_);
  not _29859_ (_25208_, _25206_);
  and _29860_ (_25209_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _29861_ (_10727_, _25209_, _25207_);
  and _29862_ (_25210_, _24476_, _24056_);
  and _29863_ (_25211_, _25210_, _23583_);
  not _29864_ (_25212_, _25210_);
  and _29865_ (_25213_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or _29866_ (_10764_, _25213_, _25211_);
  and _29867_ (_25214_, _25210_, _23887_);
  and _29868_ (_25215_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or _29869_ (_10780_, _25215_, _25214_);
  and _29870_ (_25216_, _25210_, _23548_);
  and _29871_ (_25217_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or _29872_ (_10796_, _25217_, _25216_);
  and _29873_ (_25218_, _25206_, _24051_);
  and _29874_ (_25219_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _29875_ (_10814_, _25219_, _25218_);
  and _29876_ (_25220_, _25017_, _24698_);
  and _29877_ (_25221_, _25220_, _24533_);
  nand _29878_ (_25222_, _25221_, _23504_);
  or _29879_ (_25223_, _25221_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _29880_ (_25224_, _25223_, _24539_);
  and _29881_ (_25225_, _25224_, _25222_);
  and _29882_ (_25226_, _22936_, _22906_);
  and _29883_ (_25227_, _25226_, _23944_);
  and _29884_ (_25228_, _25227_, _25024_);
  not _29885_ (_25229_, _25228_);
  or _29886_ (_25230_, _25229_, _23577_);
  or _29887_ (_25231_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _29888_ (_25232_, _25231_, _24179_);
  and _29889_ (_25233_, _25232_, _25230_);
  not _29890_ (_25234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor _29891_ (_25235_, _24178_, _25234_);
  or _29892_ (_25236_, _25235_, rst);
  or _29893_ (_25238_, _25236_, _25233_);
  or _29894_ (_10934_, _25238_, _25225_);
  and _29895_ (_25240_, _25220_, _24562_);
  nand _29896_ (_25241_, _25240_, _23504_);
  or _29897_ (_25242_, _25240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _29898_ (_25243_, _25242_, _24539_);
  and _29899_ (_25244_, _25243_, _25241_);
  or _29900_ (_25246_, _25229_, _23880_);
  or _29901_ (_25247_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _29902_ (_25248_, _25247_, _24179_);
  and _29903_ (_25249_, _25248_, _25246_);
  not _29904_ (_25250_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor _29905_ (_25251_, _24178_, _25250_);
  or _29906_ (_25252_, _25251_, rst);
  or _29907_ (_25253_, _25252_, _25249_);
  or _29908_ (_10960_, _25253_, _25244_);
  and _29909_ (_25254_, _25220_, _24177_);
  nand _29910_ (_25255_, _25254_, _23504_);
  or _29911_ (_25256_, _25254_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _29912_ (_25257_, _25256_, _24539_);
  and _29913_ (_25258_, _25257_, _25255_);
  nand _29914_ (_25259_, _25228_, _23542_);
  or _29915_ (_25260_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _29916_ (_25261_, _25260_, _24179_);
  and _29917_ (_25262_, _25261_, _25259_);
  not _29918_ (_25263_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor _29919_ (_25264_, _24178_, _25263_);
  or _29920_ (_25266_, _25264_, rst);
  or _29921_ (_25267_, _25266_, _25262_);
  or _29922_ (_10987_, _25267_, _25258_);
  and _29923_ (_25268_, _25220_, _24577_);
  nand _29924_ (_25269_, _25268_, _23504_);
  or _29925_ (_25270_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _29926_ (_25271_, _25270_, _24539_);
  and _29927_ (_25272_, _25271_, _25269_);
  nand _29928_ (_25274_, _25228_, _24210_);
  and _29929_ (_25275_, _25274_, _24179_);
  and _29930_ (_25276_, _25275_, _25270_);
  not _29931_ (_25277_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _29932_ (_25278_, _24178_, _25277_);
  or _29933_ (_25279_, _25278_, rst);
  or _29934_ (_25280_, _25279_, _25276_);
  or _29935_ (_11035_, _25280_, _25272_);
  and _29936_ (_25281_, _25210_, _24134_);
  and _29937_ (_25283_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or _29938_ (_27155_, _25283_, _25281_);
  and _29939_ (_25284_, _25210_, _24051_);
  and _29940_ (_25285_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or _29941_ (_11161_, _25285_, _25284_);
  and _29942_ (_25286_, _25220_, _24594_);
  nand _29943_ (_25287_, _25286_, _23504_);
  or _29944_ (_25288_, _25286_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _29945_ (_25289_, _25288_, _24539_);
  and _29946_ (_25290_, _25289_, _25287_);
  nand _29947_ (_25291_, _25228_, _24126_);
  or _29948_ (_25292_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _29949_ (_25293_, _25292_, _24179_);
  and _29950_ (_25294_, _25293_, _25291_);
  not _29951_ (_25295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _29952_ (_25296_, _24178_, _25295_);
  or _29953_ (_25297_, _25296_, rst);
  or _29954_ (_25298_, _25297_, _25294_);
  or _29955_ (_11255_, _25298_, _25290_);
  and _29956_ (_25299_, _25220_, _24607_);
  nand _29957_ (_25300_, _25299_, _23504_);
  or _29958_ (_25301_, _25299_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _29959_ (_25302_, _25301_, _24539_);
  and _29960_ (_25303_, _25302_, _25300_);
  nand _29961_ (_25305_, _25228_, _24043_);
  or _29962_ (_25306_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _29963_ (_25307_, _25306_, _24179_);
  and _29964_ (_25308_, _25307_, _25305_);
  and _29965_ (_25309_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _29966_ (_25310_, _25309_, rst);
  or _29967_ (_25311_, _25310_, _25308_);
  or _29968_ (_11356_, _25311_, _25303_);
  and _29969_ (_25312_, _25206_, _24134_);
  and _29970_ (_25313_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _29971_ (_11416_, _25313_, _25312_);
  and _29972_ (_25314_, _24476_, _24223_);
  and _29973_ (_25315_, _25314_, _24051_);
  not _29974_ (_25316_, _25314_);
  and _29975_ (_25318_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _29976_ (_11589_, _25318_, _25315_);
  and _29977_ (_25319_, _25123_, _24698_);
  and _29978_ (_25320_, _25319_, _24562_);
  nand _29979_ (_25321_, _25320_, _23504_);
  or _29980_ (_25322_, _25320_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _29981_ (_25323_, _25322_, _24539_);
  and _29982_ (_25325_, _25323_, _25321_);
  and _29983_ (_25327_, _25319_, _24577_);
  not _29984_ (_25328_, _25327_);
  or _29985_ (_25329_, _25328_, _23880_);
  or _29986_ (_25330_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _29987_ (_25331_, _25330_, _24179_);
  and _29988_ (_25332_, _25331_, _25329_);
  not _29989_ (_25333_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor _29990_ (_25334_, _24178_, _25333_);
  or _29991_ (_25335_, _25334_, rst);
  or _29992_ (_25336_, _25335_, _25332_);
  or _29993_ (_11618_, _25336_, _25325_);
  and _29994_ (_25338_, _25319_, _24177_);
  nand _29995_ (_25339_, _25338_, _23504_);
  or _29996_ (_25340_, _25338_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _29997_ (_25341_, _25340_, _24539_);
  and _29998_ (_25342_, _25341_, _25339_);
  nand _29999_ (_25343_, _25327_, _23542_);
  or _30000_ (_25344_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _30001_ (_25345_, _25344_, _24179_);
  and _30002_ (_25346_, _25345_, _25343_);
  not _30003_ (_25347_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor _30004_ (_25349_, _24178_, _25347_);
  or _30005_ (_25350_, _25349_, rst);
  or _30006_ (_25351_, _25350_, _25346_);
  or _30007_ (_11644_, _25351_, _25342_);
  nand _30008_ (_25353_, _25327_, _23504_);
  or _30009_ (_25354_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _30010_ (_25355_, _25354_, _24539_);
  and _30011_ (_25356_, _25355_, _25353_);
  nand _30012_ (_25357_, _25327_, _24210_);
  and _30013_ (_25358_, _25357_, _24179_);
  and _30014_ (_25359_, _25358_, _25354_);
  not _30015_ (_25360_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _30016_ (_25361_, _24178_, _25360_);
  or _30017_ (_25362_, _25361_, rst);
  or _30018_ (_25363_, _25362_, _25359_);
  or _30019_ (_11669_, _25363_, _25356_);
  and _30020_ (_25364_, _25314_, _24089_);
  and _30021_ (_25365_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _30022_ (_27122_, _25365_, _25364_);
  and _30023_ (_25366_, _25319_, _24607_);
  nand _30024_ (_25367_, _25366_, _23504_);
  or _30025_ (_25368_, _25366_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _30026_ (_25369_, _25368_, _24539_);
  and _30027_ (_25370_, _25369_, _25367_);
  nand _30028_ (_25371_, _25327_, _24043_);
  or _30029_ (_25372_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _30030_ (_25374_, _25372_, _24179_);
  and _30031_ (_25375_, _25374_, _25371_);
  and _30032_ (_25376_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _30033_ (_25377_, _25376_, rst);
  or _30034_ (_25378_, _25377_, _25375_);
  or _30035_ (_11891_, _25378_, _25370_);
  and _30036_ (_25380_, _25206_, _24219_);
  and _30037_ (_25381_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _30038_ (_27036_, _25381_, _25380_);
  and _30039_ (_25382_, _25319_, _24594_);
  nand _30040_ (_25383_, _25382_, _23504_);
  or _30041_ (_25384_, _25382_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _30042_ (_25385_, _25384_, _24539_);
  and _30043_ (_25386_, _25385_, _25383_);
  nand _30044_ (_25387_, _25327_, _24126_);
  or _30045_ (_25388_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _30046_ (_25390_, _25388_, _24179_);
  and _30047_ (_25391_, _25390_, _25387_);
  not _30048_ (_25392_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _30049_ (_25393_, _24178_, _25392_);
  or _30050_ (_25394_, _25393_, rst);
  or _30051_ (_25395_, _25394_, _25391_);
  or _30052_ (_11973_, _25395_, _25386_);
  not _30053_ (_25396_, _25319_);
  or _30054_ (_25397_, _25396_, _24643_);
  and _30055_ (_25398_, _25397_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _30056_ (_25400_, _24638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _30057_ (_25401_, _25400_, _24637_);
  and _30058_ (_25402_, _25401_, _25319_);
  or _30059_ (_25403_, _25402_, _25398_);
  and _30060_ (_25404_, _25403_, _24539_);
  nand _30061_ (_25405_, _25327_, _24082_);
  or _30062_ (_25406_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _30063_ (_25407_, _25406_, _24179_);
  and _30064_ (_25408_, _25407_, _25405_);
  not _30065_ (_25409_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor _30066_ (_25410_, _24178_, _25409_);
  or _30067_ (_25411_, _25410_, rst);
  or _30068_ (_25412_, _25411_, _25408_);
  or _30069_ (_11994_, _25412_, _25404_);
  and _30070_ (_25413_, _24004_, _23943_);
  and _30071_ (_25414_, _25413_, _24146_);
  and _30072_ (_25415_, _25414_, _23548_);
  not _30073_ (_25416_, _25414_);
  and _30074_ (_25417_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or _30075_ (_12065_, _25417_, _25415_);
  and _30076_ (_25418_, _25314_, _23996_);
  and _30077_ (_25420_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _30078_ (_12243_, _25420_, _25418_);
  and _30079_ (_25421_, _25314_, _24134_);
  and _30080_ (_25422_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _30081_ (_12266_, _25422_, _25421_);
  and _30082_ (_25423_, _25206_, _23887_);
  and _30083_ (_25424_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _30084_ (_12515_, _25424_, _25423_);
  and _30085_ (_25425_, _25206_, _23548_);
  and _30086_ (_25426_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _30087_ (_12616_, _25426_, _25425_);
  and _30088_ (_25428_, _25314_, _24219_);
  and _30089_ (_25429_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _30090_ (_12637_, _25429_, _25428_);
  and _30091_ (_25430_, _24302_, _24051_);
  and _30092_ (_25431_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or _30093_ (_27231_, _25431_, _25430_);
  and _30094_ (_25432_, _24476_, _24319_);
  and _30095_ (_25433_, _25432_, _23996_);
  not _30096_ (_25434_, _25432_);
  and _30097_ (_25435_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _30098_ (_27100_, _25435_, _25433_);
  and _30099_ (_25436_, _25432_, _24134_);
  and _30100_ (_25438_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _30101_ (_12748_, _25438_, _25436_);
  and _30102_ (_25440_, _24302_, _24089_);
  and _30103_ (_25441_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or _30104_ (_14268_, _25441_, _25440_);
  and _30105_ (_25442_, _24146_, _23945_);
  and _30106_ (_25443_, _25442_, _24089_);
  not _30107_ (_25444_, _25442_);
  and _30108_ (_25445_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _30109_ (_15162_, _25445_, _25443_);
  and _30110_ (_25446_, _25314_, _23887_);
  and _30111_ (_25447_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _30112_ (_15213_, _25447_, _25446_);
  and _30113_ (_25448_, _25442_, _23583_);
  and _30114_ (_25449_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _30115_ (_15234_, _25449_, _25448_);
  and _30116_ (_25450_, _25314_, _23548_);
  and _30117_ (_25451_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _30118_ (_15619_, _25451_, _25450_);
  nor _30119_ (_25453_, _22737_, _23011_);
  not _30120_ (_25454_, _22737_);
  and _30121_ (_25455_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _30122_ (_25456_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  not _30123_ (_25457_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _30124_ (_25458_, _23601_, _25457_);
  nor _30125_ (_25459_, _25458_, _25456_);
  and _30126_ (_25460_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _30127_ (_25461_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _30128_ (_25462_, _25461_, _25460_);
  and _30129_ (_25463_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _30130_ (_25465_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _30131_ (_25466_, _25465_, _25463_);
  and _30132_ (_25467_, _25466_, _25462_);
  and _30133_ (_25469_, _25467_, _25459_);
  nor _30134_ (_25470_, _25469_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _30135_ (_25472_, _25470_, _25455_);
  nor _30136_ (_25473_, _25472_, _25454_);
  nor _30137_ (_25475_, _25473_, _25453_);
  nor _30138_ (_26877_[7], _25475_, rst);
  nor _30139_ (_26840_[3], _23615_, rst);
  or _30140_ (_25477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _30141_ (_25478_, _22968_, _22937_);
  and _30142_ (_25479_, _25478_, _24620_);
  or _30143_ (_25480_, _25479_, _25477_);
  and _30144_ (_25481_, _24532_, _24550_);
  and _30145_ (_25482_, _25481_, _24531_);
  not _30146_ (_25483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _30147_ (_25484_, _25481_, _25483_);
  nand _30148_ (_25485_, _25484_, _25479_);
  or _30149_ (_25486_, _25485_, _25482_);
  and _30150_ (_25487_, _25486_, _25480_);
  and _30151_ (_25488_, _24173_, _24004_);
  and _30152_ (_25489_, _25488_, _24628_);
  or _30153_ (_25490_, _25489_, _25487_);
  nand _30154_ (_25491_, _25489_, _23989_);
  and _30155_ (_25492_, _25491_, _22731_);
  and _30156_ (_17618_, _25492_, _25490_);
  and _30157_ (_25493_, _25442_, _24134_);
  and _30158_ (_25494_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _30159_ (_27034_, _25494_, _25493_);
  and _30160_ (_25495_, _25432_, _24219_);
  and _30161_ (_25496_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _30162_ (_27099_, _25496_, _25495_);
  and _30163_ (_25497_, _24636_, _24181_);
  and _30164_ (_25499_, _25497_, _25488_);
  and _30165_ (_25500_, _24607_, _24181_);
  and _30166_ (_25501_, _25500_, _25488_);
  nor _30167_ (_25502_, _25501_, _25499_);
  or _30168_ (_25503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _30169_ (_25504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _30170_ (_25505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _25504_);
  and _30171_ (_25506_, _25505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _30172_ (_25507_, _25506_, _25503_);
  and _30173_ (_25508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _30174_ (_25509_, _25508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _30175_ (_25510_, _25509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _30176_ (_25511_, _25510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _30177_ (_25512_, _25511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _30178_ (_25513_, _25512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _30179_ (_25514_, _25513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _30180_ (_25515_, _25514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _30181_ (_25516_, _25515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _30182_ (_25517_, _25516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _30183_ (_25518_, _25517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _30184_ (_25519_, _25518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _30185_ (_25520_, _25519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _30186_ (_25521_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _30187_ (_25522_, _25521_, _25520_);
  and _30188_ (_25523_, _25522_, _25507_);
  nor _30189_ (_25524_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not _30190_ (_25526_, _25524_);
  not _30191_ (_25527_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _30192_ (_25528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _30193_ (_25529_, _25528_, _25524_);
  and _30194_ (_25531_, _25529_, _25527_);
  nor _30195_ (_25532_, _25531_, _25526_);
  nand _30196_ (_25533_, _25532_, _25523_);
  nand _30197_ (_25534_, _25533_, _25502_);
  or _30198_ (_25535_, _25502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _30199_ (_25536_, _25535_, _22731_);
  and _30200_ (_17752_, _25536_, _25534_);
  and _30201_ (_25538_, _25524_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not _30202_ (_25539_, _25538_);
  or _30203_ (_25540_, _25529_, _25523_);
  and _30204_ (_25541_, _25540_, _25539_);
  and _30205_ (_25542_, _25541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _30206_ (_25543_, _25520_, _25507_);
  and _30207_ (_25544_, _25543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _30208_ (_25545_, _25544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor _30209_ (_25546_, _25531_, _25523_);
  or _30210_ (_25547_, _25546_, _25499_);
  and _30211_ (_25548_, _25547_, _25545_);
  or _30212_ (_25549_, _25548_, _25542_);
  not _30213_ (_25550_, _25499_);
  nor _30214_ (_25551_, _25550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor _30215_ (_25552_, _25551_, _25501_);
  and _30216_ (_25553_, _25552_, _25549_);
  not _30217_ (_25554_, _23989_);
  and _30218_ (_25556_, _24607_, _22868_);
  and _30219_ (_25557_, _25556_, _24179_);
  and _30220_ (_25558_, _25557_, _25488_);
  and _30221_ (_25560_, _25558_, _25554_);
  or _30222_ (_25561_, _25560_, _25553_);
  and _30223_ (_17768_, _25561_, _22731_);
  nor _30224_ (_25563_, _22737_, _23133_);
  and _30225_ (_25564_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _30226_ (_25565_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _30227_ (_25566_, _25565_, _25564_);
  and _30228_ (_25567_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _30229_ (_25568_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _30230_ (_25569_, _25568_, _25567_);
  and _30231_ (_25571_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _30232_ (_25572_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _30233_ (_25573_, _25572_, _25571_);
  and _30234_ (_25574_, _25573_, _25569_);
  and _30235_ (_25575_, _25574_, _25566_);
  nor _30236_ (_25576_, _25575_, _24471_);
  nor _30237_ (_25577_, _25576_, _25563_);
  nor _30238_ (_26867_[4], _25577_, rst);
  nor _30239_ (_25578_, _25550_, _23989_);
  not _30240_ (_25579_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _30241_ (_25580_, _25538_, _25579_);
  and _30242_ (_25581_, _25580_, _25523_);
  and _30243_ (_25582_, _25513_, _25507_);
  or _30244_ (_25583_, _25582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _30245_ (_25584_, _25582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _30246_ (_25585_, _25584_, _25583_);
  or _30247_ (_25586_, _25585_, _25531_);
  or _30248_ (_25587_, _25586_, _25581_);
  nand _30249_ (_25588_, _25531_, _25579_);
  and _30250_ (_25589_, _25588_, _25502_);
  and _30251_ (_25590_, _25589_, _25587_);
  and _30252_ (_25591_, _25558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _30253_ (_25592_, _25591_, _25590_);
  or _30254_ (_25593_, _25592_, _25578_);
  and _30255_ (_17818_, _25593_, _22731_);
  and _30256_ (_25594_, _25526_, _25507_);
  and _30257_ (_25596_, _25594_, _25502_);
  or _30258_ (_25597_, _25596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _30259_ (_25598_, _25522_);
  nand _30260_ (_25599_, _25596_, _25598_);
  and _30261_ (_25600_, _25599_, _22731_);
  and _30262_ (_17853_, _25600_, _25597_);
  and _30263_ (_25601_, _24533_, _22868_);
  and _30264_ (_25602_, _25601_, _24179_);
  and _30265_ (_25603_, _25602_, _25488_);
  nand _30266_ (_25604_, _25603_, _23989_);
  and _30267_ (_25605_, _25538_, _25528_);
  not _30268_ (_25606_, _25605_);
  and _30269_ (_25607_, _24562_, _24181_);
  and _30270_ (_25608_, _25607_, _25488_);
  nor _30271_ (_25609_, _25608_, _25606_);
  not _30272_ (_25610_, _25609_);
  and _30273_ (_25611_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _30274_ (_25612_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _30275_ (_25613_, _25612_, _25611_);
  or _30276_ (_25614_, _25603_, _25613_);
  and _30277_ (_25615_, _25614_, _22731_);
  and _30278_ (_17922_, _25615_, _25604_);
  nand _30279_ (_25616_, _25608_, _23989_);
  not _30280_ (_25617_, _25603_);
  nor _30281_ (_25618_, _25605_, _25579_);
  and _30282_ (_25619_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _30283_ (_25620_, _25619_, _25618_);
  or _30284_ (_25621_, _25620_, _25608_);
  and _30285_ (_25622_, _25621_, _25617_);
  and _30286_ (_25623_, _25622_, _25616_);
  and _30287_ (_25625_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _30288_ (_25626_, _25625_, _25623_);
  and _30289_ (_17942_, _25626_, _22731_);
  and _30290_ (_17956_, t2ex_i, _22731_);
  and _30291_ (_25627_, _24476_, _22974_);
  and _30292_ (_25628_, _25627_, _23996_);
  not _30293_ (_25629_, _25627_);
  and _30294_ (_25630_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or _30295_ (_17998_, _25630_, _25628_);
  and _30296_ (_25631_, _24350_, _24089_);
  and _30297_ (_25632_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _30298_ (_27060_, _25632_, _25631_);
  nand _30299_ (_25633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _22731_);
  nor _30300_ (_18105_, _25633_, t2ex_i);
  nor _30301_ (_25634_, t2_i, rst);
  and _30302_ (_18119_, _25634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and _30303_ (_18134_, t2_i, _22731_);
  and _30304_ (_25635_, _24350_, _23996_);
  and _30305_ (_25636_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _30306_ (_18155_, _25636_, _25635_);
  and _30307_ (_25637_, _24301_, _24223_);
  and _30308_ (_25639_, _25637_, _24219_);
  not _30309_ (_25640_, _25637_);
  and _30310_ (_25642_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _30311_ (_18176_, _25642_, _25639_);
  and _30312_ (_25643_, _25432_, _23887_);
  and _30313_ (_25644_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _30314_ (_18441_, _25644_, _25643_);
  and _30315_ (_25645_, _25432_, _23583_);
  and _30316_ (_25647_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _30317_ (_18950_, _25647_, _25645_);
  and _30318_ (_25648_, _24140_, _23945_);
  and _30319_ (_25649_, _25648_, _23996_);
  not _30320_ (_25650_, _25648_);
  and _30321_ (_25651_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or _30322_ (_19201_, _25651_, _25649_);
  and _30323_ (_25652_, _25627_, _24219_);
  and _30324_ (_25654_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or _30325_ (_19605_, _25654_, _25652_);
  and _30326_ (_25656_, _25627_, _23887_);
  and _30327_ (_25657_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or _30328_ (_19639_, _25657_, _25656_);
  and _30329_ (_25658_, _24496_, _24056_);
  and _30330_ (_25659_, _25658_, _24134_);
  not _30331_ (_25660_, _25658_);
  and _30332_ (_25661_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _30333_ (_19907_, _25661_, _25659_);
  and _30334_ (_25662_, _25627_, _23548_);
  and _30335_ (_25663_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or _30336_ (_27090_, _25663_, _25662_);
  and _30337_ (_25664_, _25442_, _24219_);
  and _30338_ (_25665_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _30339_ (_27033_, _25665_, _25664_);
  and _30340_ (_25666_, _25627_, _24051_);
  and _30341_ (_25668_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or _30342_ (_21388_, _25668_, _25666_);
  and _30343_ (_25669_, _25627_, _24089_);
  and _30344_ (_25670_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or _30345_ (_21519_, _25670_, _25669_);
  and _30346_ (_25672_, _24365_, _24016_);
  and _30347_ (_25673_, _25672_, _24051_);
  not _30348_ (_25674_, _25672_);
  and _30349_ (_25675_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _30350_ (_21620_, _25675_, _25673_);
  and _30351_ (_25677_, _25627_, _23583_);
  and _30352_ (_25679_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or _30353_ (_21642_, _25679_, _25677_);
  and _30354_ (_26865_[0], _23685_, _22731_);
  and _30355_ (_26865_[1], _23664_, _22731_);
  and _30356_ (_26865_[2], _23643_, _22731_);
  and _30357_ (_25681_, _25024_, _24179_);
  and _30358_ (_25682_, _25226_, _24004_);
  and _30359_ (_25683_, _25682_, _25681_);
  not _30360_ (_25684_, _25683_);
  and _30361_ (_25685_, _25684_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _30362_ (_25686_, _25683_, _23577_);
  or _30363_ (_25687_, _25686_, _25685_);
  and _30364_ (_26865_[3], _25687_, _22731_);
  and _30365_ (_25689_, _25648_, _24089_);
  and _30366_ (_25691_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or _30367_ (_27031_, _25691_, _25689_);
  nor _30368_ (_25692_, _23592_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _30369_ (_25693_, _25692_, _25454_);
  nor _30370_ (_25694_, _25693_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _30371_ (_25695_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  not _30372_ (_25696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand _30373_ (_25697_, _25694_, _25696_);
  and _30374_ (_25698_, _25697_, _22731_);
  and _30375_ (_26883_[0], _25698_, _25695_);
  or _30376_ (_25699_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  not _30377_ (_25700_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand _30378_ (_25701_, _25694_, _25700_);
  and _30379_ (_25703_, _25701_, _22731_);
  and _30380_ (_26883_[1], _25703_, _25699_);
  or _30381_ (_25704_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  not _30382_ (_25705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand _30383_ (_25707_, _25694_, _25705_);
  and _30384_ (_25709_, _25707_, _22731_);
  and _30385_ (_26883_[2], _25709_, _25704_);
  or _30386_ (_25710_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not _30387_ (_25711_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand _30388_ (_25712_, _25694_, _25711_);
  and _30389_ (_25713_, _25712_, _22731_);
  and _30390_ (_26883_[3], _25713_, _25710_);
  or _30391_ (_25714_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not _30392_ (_25715_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand _30393_ (_25716_, _25694_, _25715_);
  and _30394_ (_25718_, _25716_, _22731_);
  and _30395_ (_26883_[4], _25718_, _25714_);
  or _30396_ (_25719_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not _30397_ (_25720_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand _30398_ (_25721_, _25694_, _25720_);
  and _30399_ (_25722_, _25721_, _22731_);
  and _30400_ (_26883_[5], _25722_, _25719_);
  or _30401_ (_25723_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  not _30402_ (_25724_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand _30403_ (_25726_, _25694_, _25724_);
  and _30404_ (_25727_, _25726_, _22731_);
  and _30405_ (_26883_[6], _25727_, _25723_);
  or _30406_ (_25728_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  not _30407_ (_25729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand _30408_ (_25730_, _25694_, _25729_);
  and _30409_ (_25732_, _25730_, _22731_);
  and _30410_ (_26883_[7], _25732_, _25728_);
  or _30411_ (_25734_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not _30412_ (_25735_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _30413_ (_25736_, _25694_, _25735_);
  and _30414_ (_25737_, _25736_, _22731_);
  and _30415_ (_26883_[8], _25737_, _25734_);
  or _30416_ (_25738_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  not _30417_ (_25739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _30418_ (_25740_, _25694_, _25739_);
  and _30419_ (_25741_, _25740_, _22731_);
  and _30420_ (_26883_[9], _25741_, _25738_);
  or _30421_ (_25743_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  not _30422_ (_25744_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand _30423_ (_25745_, _25694_, _25744_);
  and _30424_ (_25746_, _25745_, _22731_);
  and _30425_ (_26883_[10], _25746_, _25743_);
  or _30426_ (_25748_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  not _30427_ (_25750_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _30428_ (_25751_, _25694_, _25750_);
  and _30429_ (_25752_, _25751_, _22731_);
  and _30430_ (_26883_[11], _25752_, _25748_);
  or _30431_ (_25753_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  not _30432_ (_25754_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand _30433_ (_25755_, _25694_, _25754_);
  and _30434_ (_25756_, _25755_, _22731_);
  and _30435_ (_26883_[12], _25756_, _25753_);
  or _30436_ (_25757_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not _30437_ (_25758_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _30438_ (_25759_, _25694_, _25758_);
  and _30439_ (_25760_, _25759_, _22731_);
  and _30440_ (_26883_[13], _25760_, _25757_);
  or _30441_ (_25761_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  not _30442_ (_25763_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _30443_ (_25764_, _25694_, _25763_);
  and _30444_ (_25765_, _25764_, _22731_);
  and _30445_ (_26883_[14], _25765_, _25761_);
  or _30446_ (_25766_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  not _30447_ (_25767_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _30448_ (_25768_, _25694_, _25767_);
  and _30449_ (_25769_, _25768_, _22731_);
  and _30450_ (_26883_[15], _25769_, _25766_);
  or _30451_ (_25770_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  not _30452_ (_25771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _30453_ (_25772_, _25694_, _25771_);
  and _30454_ (_25773_, _25772_, _22731_);
  and _30455_ (_26883_[16], _25773_, _25770_);
  or _30456_ (_25775_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not _30457_ (_25776_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _30458_ (_25777_, _25694_, _25776_);
  and _30459_ (_25778_, _25777_, _22731_);
  and _30460_ (_26883_[17], _25778_, _25775_);
  or _30461_ (_25779_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not _30462_ (_25780_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _30463_ (_25781_, _25694_, _25780_);
  and _30464_ (_25782_, _25781_, _22731_);
  and _30465_ (_26883_[18], _25782_, _25779_);
  or _30466_ (_25783_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not _30467_ (_25784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _30468_ (_25785_, _25694_, _25784_);
  and _30469_ (_25786_, _25785_, _22731_);
  and _30470_ (_26883_[19], _25786_, _25783_);
  or _30471_ (_25787_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  not _30472_ (_25788_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand _30473_ (_25789_, _25694_, _25788_);
  and _30474_ (_25790_, _25789_, _22731_);
  and _30475_ (_26883_[20], _25790_, _25787_);
  or _30476_ (_25791_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  not _30477_ (_25792_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _30478_ (_25793_, _25694_, _25792_);
  and _30479_ (_25794_, _25793_, _22731_);
  and _30480_ (_26883_[21], _25794_, _25791_);
  or _30481_ (_25795_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not _30482_ (_25796_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _30483_ (_25797_, _25694_, _25796_);
  and _30484_ (_25798_, _25797_, _22731_);
  and _30485_ (_26883_[22], _25798_, _25795_);
  or _30486_ (_25799_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not _30487_ (_25800_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _30488_ (_25801_, _25694_, _25800_);
  and _30489_ (_25802_, _25801_, _22731_);
  and _30490_ (_26883_[23], _25802_, _25799_);
  or _30491_ (_25803_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  not _30492_ (_25804_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand _30493_ (_25805_, _25694_, _25804_);
  and _30494_ (_25806_, _25805_, _22731_);
  and _30495_ (_26883_[24], _25806_, _25803_);
  or _30496_ (_25807_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  not _30497_ (_25808_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _30498_ (_25809_, _25694_, _25808_);
  and _30499_ (_25810_, _25809_, _22731_);
  and _30500_ (_26883_[25], _25810_, _25807_);
  or _30501_ (_25811_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not _30502_ (_25812_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _30503_ (_25813_, _25694_, _25812_);
  and _30504_ (_25814_, _25813_, _22731_);
  and _30505_ (_26883_[26], _25814_, _25811_);
  or _30506_ (_25815_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not _30507_ (_25816_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _30508_ (_25817_, _25694_, _25816_);
  and _30509_ (_25818_, _25817_, _22731_);
  and _30510_ (_26883_[27], _25818_, _25815_);
  or _30511_ (_25819_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  not _30512_ (_25820_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand _30513_ (_25821_, _25694_, _25820_);
  and _30514_ (_25822_, _25821_, _22731_);
  and _30515_ (_26883_[28], _25822_, _25819_);
  or _30516_ (_25823_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not _30517_ (_25825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _30518_ (_25826_, _25694_, _25825_);
  and _30519_ (_25827_, _25826_, _22731_);
  and _30520_ (_26883_[29], _25827_, _25823_);
  or _30521_ (_25828_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not _30522_ (_25829_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand _30523_ (_25830_, _25694_, _25829_);
  and _30524_ (_25831_, _25830_, _22731_);
  and _30525_ (_26883_[30], _25831_, _25828_);
  and _30526_ (_25832_, _25684_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _30527_ (_25833_, _25684_, _24082_);
  nor _30528_ (_25834_, _25833_, _25832_);
  nor _30529_ (_25835_, _25834_, _22906_);
  and _30530_ (_25836_, _25834_, _22906_);
  nor _30531_ (_25837_, _25836_, _25835_);
  or _30532_ (_25838_, _25687_, _22867_);
  nor _30533_ (_25839_, _25686_, _25685_);
  or _30534_ (_25840_, _25839_, _22868_);
  and _30535_ (_25841_, _23685_, _22886_);
  nor _30536_ (_25842_, _23685_, _22886_);
  nor _30537_ (_25844_, _25842_, _25841_);
  and _30538_ (_25845_, _24176_, _22978_);
  and _30539_ (_25846_, _25845_, _24298_);
  and _30540_ (_25848_, _25846_, _25844_);
  and _30541_ (_25849_, _25848_, _22936_);
  and _30542_ (_25850_, _25849_, _25840_);
  and _30543_ (_25851_, _25850_, _25838_);
  and _30544_ (_25852_, _25851_, _25837_);
  and _30545_ (_25854_, _25852_, _24210_);
  not _30546_ (_25855_, _25834_);
  and _30547_ (_25856_, _25687_, _23685_);
  and _30548_ (_25858_, _25856_, _25855_);
  nand _30549_ (_25859_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _30550_ (_25860_, _25839_, _23791_);
  and _30551_ (_25861_, _25860_, _25834_);
  nand _30552_ (_25862_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _30553_ (_25863_, _25862_, _25859_);
  and _30554_ (_25864_, _25687_, _23791_);
  and _30555_ (_25865_, _25864_, _25855_);
  nand _30556_ (_25866_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _30557_ (_25867_, _25856_, _25834_);
  nand _30558_ (_25868_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _30559_ (_25869_, _25868_, _25866_);
  and _30560_ (_25870_, _25869_, _25863_);
  not _30561_ (_25872_, _25852_);
  and _30562_ (_25873_, _25839_, _23685_);
  and _30563_ (_25874_, _25873_, _25855_);
  nand _30564_ (_25876_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _30565_ (_25877_, _25873_, _25834_);
  nand _30566_ (_25878_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _30567_ (_25879_, _25878_, _25876_);
  and _30568_ (_25880_, _25860_, _25855_);
  nand _30569_ (_25881_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _30570_ (_25882_, _25864_, _25834_);
  nand _30571_ (_25884_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _30572_ (_25885_, _25884_, _25881_);
  and _30573_ (_25886_, _25885_, _25879_);
  and _30574_ (_25888_, _25886_, _25872_);
  and _30575_ (_25890_, _25888_, _25870_);
  nor _30576_ (_25891_, _25890_, _25854_);
  and _30577_ (_26866_[0], _25891_, _22731_);
  and _30578_ (_25892_, _25852_, _23542_);
  and _30579_ (_25893_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _30580_ (_25894_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _30581_ (_25895_, _25894_, _25893_);
  and _30582_ (_25896_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _30583_ (_25897_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _30584_ (_25898_, _25897_, _25896_);
  and _30585_ (_25899_, _25898_, _25895_);
  and _30586_ (_25900_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _30587_ (_25901_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _30588_ (_25902_, _25901_, _25900_);
  and _30589_ (_25903_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _30590_ (_25905_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _30591_ (_25907_, _25905_, _25903_);
  and _30592_ (_25908_, _25907_, _25902_);
  and _30593_ (_25909_, _25908_, _25872_);
  and _30594_ (_25910_, _25909_, _25899_);
  nor _30595_ (_25911_, _25910_, _25892_);
  and _30596_ (_26866_[1], _25911_, _22731_);
  nor _30597_ (_25912_, _25872_, _23880_);
  and _30598_ (_25913_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _30599_ (_25914_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _30600_ (_25915_, _25914_, _25913_);
  and _30601_ (_25916_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _30602_ (_25917_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _30603_ (_25918_, _25917_, _25916_);
  and _30604_ (_25919_, _25918_, _25915_);
  and _30605_ (_25920_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and _30606_ (_25921_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _30607_ (_25922_, _25921_, _25920_);
  and _30608_ (_25923_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _30609_ (_25924_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _30610_ (_25925_, _25924_, _25923_);
  and _30611_ (_25926_, _25925_, _25922_);
  and _30612_ (_25928_, _25926_, _25872_);
  and _30613_ (_25929_, _25928_, _25919_);
  nor _30614_ (_25930_, _25929_, _25912_);
  and _30615_ (_26866_[2], _25930_, _22731_);
  and _30616_ (_25931_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _30617_ (_25932_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _30618_ (_25933_, _25932_, _25931_);
  and _30619_ (_25934_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _30620_ (_25935_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _30621_ (_25936_, _25935_, _25934_);
  and _30622_ (_25937_, _25936_, _25933_);
  nand _30623_ (_25938_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nand _30624_ (_25940_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _30625_ (_25941_, _25940_, _25938_);
  nand _30626_ (_25942_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nand _30627_ (_25944_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _30628_ (_25945_, _25944_, _25942_);
  and _30629_ (_25947_, _25945_, _25941_);
  and _30630_ (_25948_, _25947_, _25872_);
  and _30631_ (_25950_, _25948_, _25937_);
  not _30632_ (_25951_, _23577_);
  and _30633_ (_25952_, _25852_, _25951_);
  nor _30634_ (_25954_, _25952_, _25950_);
  and _30635_ (_26866_[3], _25954_, _22731_);
  and _30636_ (_25955_, _25852_, _24082_);
  and _30637_ (_25956_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _30638_ (_25958_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _30639_ (_25959_, _25958_, _25956_);
  and _30640_ (_25961_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _30641_ (_25962_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _30642_ (_25963_, _25962_, _25961_);
  and _30643_ (_25964_, _25963_, _25959_);
  and _30644_ (_25965_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _30645_ (_25967_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor _30646_ (_25968_, _25967_, _25965_);
  and _30647_ (_25969_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _30648_ (_25970_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _30649_ (_25971_, _25970_, _25969_);
  and _30650_ (_25973_, _25971_, _25968_);
  and _30651_ (_25974_, _25973_, _25872_);
  and _30652_ (_25975_, _25974_, _25964_);
  nor _30653_ (_25976_, _25975_, _25955_);
  and _30654_ (_26866_[4], _25976_, _22731_);
  and _30655_ (_25977_, _25852_, _24043_);
  and _30656_ (_25978_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _30657_ (_25979_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _30658_ (_25980_, _25979_, _25978_);
  and _30659_ (_25981_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _30660_ (_25982_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _30661_ (_25983_, _25982_, _25981_);
  and _30662_ (_25984_, _25983_, _25980_);
  and _30663_ (_25985_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _30664_ (_25986_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _30665_ (_25987_, _25986_, _25985_);
  and _30666_ (_25988_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _30667_ (_25989_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _30668_ (_25990_, _25989_, _25988_);
  and _30669_ (_25991_, _25990_, _25987_);
  and _30670_ (_25992_, _25991_, _25872_);
  and _30671_ (_25994_, _25992_, _25984_);
  nor _30672_ (_25995_, _25994_, _25977_);
  and _30673_ (_26866_[5], _25995_, _22731_);
  and _30674_ (_25997_, _25852_, _24126_);
  and _30675_ (_25998_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _30676_ (_25999_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor _30677_ (_26000_, _25999_, _25998_);
  and _30678_ (_26001_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _30679_ (_26002_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor _30680_ (_26003_, _26002_, _26001_);
  and _30681_ (_26005_, _26003_, _26000_);
  and _30682_ (_26006_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _30683_ (_26007_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _30684_ (_26008_, _26007_, _26006_);
  and _30685_ (_26010_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _30686_ (_26011_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _30687_ (_26013_, _26011_, _26010_);
  and _30688_ (_26014_, _26013_, _26008_);
  and _30689_ (_26016_, _26014_, _25872_);
  and _30690_ (_26017_, _26016_, _26005_);
  nor _30691_ (_26018_, _26017_, _25997_);
  and _30692_ (_26866_[6], _26018_, _22731_);
  and _30693_ (_26020_, _24476_, _24095_);
  and _30694_ (_26021_, _26020_, _23583_);
  not _30695_ (_26022_, _26020_);
  and _30696_ (_26023_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or _30697_ (_22612_, _26023_, _26021_);
  and _30698_ (_26024_, _26020_, _23887_);
  and _30699_ (_26025_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or _30700_ (_22613_, _26025_, _26024_);
  and _30701_ (_26027_, _25648_, _23583_);
  and _30702_ (_26028_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or _30703_ (_27030_, _26028_, _26027_);
  and _30704_ (_26031_, _24051_, _22983_);
  and _30705_ (_26032_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or _30706_ (_22614_, _26032_, _26031_);
  and _30707_ (_26034_, _26020_, _23548_);
  and _30708_ (_26035_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or _30709_ (_22615_, _26035_, _26034_);
  nor _30710_ (_26036_, _22737_, _23097_);
  and _30711_ (_26037_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _30712_ (_26038_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _30713_ (_26039_, _26038_, _26037_);
  and _30714_ (_26040_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _30715_ (_26041_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _30716_ (_26042_, _26041_, _26040_);
  and _30717_ (_26043_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _30718_ (_26044_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _30719_ (_26045_, _26044_, _26043_);
  and _30720_ (_26047_, _26045_, _26042_);
  and _30721_ (_26048_, _26047_, _26039_);
  nor _30722_ (_26049_, _26048_, _24471_);
  nor _30723_ (_26050_, _26049_, _26036_);
  nor _30724_ (_26867_[5], _26050_, rst);
  nor _30725_ (_26051_, _22737_, _23248_);
  and _30726_ (_26053_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _30727_ (_26054_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _30728_ (_26055_, _26054_, _26053_);
  and _30729_ (_26057_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _30730_ (_26058_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _30731_ (_26059_, _26058_, _26057_);
  and _30732_ (_26060_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _30733_ (_26061_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _30734_ (_26063_, _26061_, _26060_);
  and _30735_ (_26064_, _26063_, _26059_);
  and _30736_ (_26066_, _26064_, _26055_);
  nor _30737_ (_26067_, _26066_, _24471_);
  nor _30738_ (_26068_, _26067_, _26051_);
  nor _30739_ (_26867_[1], _26068_, rst);
  and _30740_ (_26840_[4], _23703_, _22731_);
  nor _30741_ (_26070_, _22737_, _23095_);
  and _30742_ (_26071_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _30743_ (_26072_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _30744_ (_26073_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _30745_ (_26074_, _26073_, _26072_);
  and _30746_ (_26076_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _30747_ (_26077_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _30748_ (_26079_, _26077_, _26076_);
  and _30749_ (_26080_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _30750_ (_26081_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _30751_ (_26082_, _26081_, _26080_);
  and _30752_ (_26083_, _26082_, _26079_);
  and _30753_ (_26084_, _26083_, _26074_);
  nor _30754_ (_26085_, _26084_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _30755_ (_26087_, _26085_, _26071_);
  nor _30756_ (_26088_, _26087_, _25454_);
  nor _30757_ (_26089_, _26088_, _26070_);
  nor _30758_ (_26877_[5], _26089_, rst);
  nor _30759_ (_26090_, _22737_, _23060_);
  and _30760_ (_26091_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _30761_ (_26092_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _30762_ (_26093_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _30763_ (_26094_, _26093_, _26092_);
  and _30764_ (_26095_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _30765_ (_26097_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _30766_ (_26098_, _26097_, _26095_);
  and _30767_ (_26099_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _30768_ (_26100_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _30769_ (_26101_, _26100_, _26099_);
  and _30770_ (_26102_, _26101_, _26098_);
  and _30771_ (_26103_, _26102_, _26094_);
  nor _30772_ (_26104_, _26103_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _30773_ (_26106_, _26104_, _26091_);
  nor _30774_ (_26107_, _26106_, _25454_);
  nor _30775_ (_26108_, _26107_, _26090_);
  nor _30776_ (_26877_[6], _26108_, rst);
  and _30777_ (_26110_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _30778_ (_26111_, _22740_, _22806_);
  or _30779_ (_26112_, _26111_, _26110_);
  and _30780_ (_26862_[14], _26112_, _22731_);
  and _30781_ (_26113_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _30782_ (_26114_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _30783_ (_26115_, _22740_, _26114_);
  or _30784_ (_26116_, _26115_, _26113_);
  and _30785_ (_26862_[13], _26116_, _22731_);
  and _30786_ (_26118_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _30787_ (_26119_, _22740_, _22797_);
  or _30788_ (_26120_, _26119_, _26118_);
  and _30789_ (_26862_[12], _26120_, _22731_);
  and _30790_ (_26121_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _30791_ (_26122_, _22740_, _22793_);
  or _30792_ (_26123_, _26122_, _26121_);
  and _30793_ (_26862_[11], _26123_, _22731_);
  and _30794_ (_26124_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _30795_ (_26125_, _22740_, _22789_);
  or _30796_ (_26126_, _26125_, _26124_);
  and _30797_ (_26862_[10], _26126_, _22731_);
  and _30798_ (_26127_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not _30799_ (_26128_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _30800_ (_26129_, _22740_, _26128_);
  or _30801_ (_26130_, _26129_, _26127_);
  and _30802_ (_26862_[9], _26130_, _22731_);
  and _30803_ (_26131_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _30804_ (_26132_, _22740_, _22780_);
  or _30805_ (_26133_, _26132_, _26131_);
  and _30806_ (_26862_[8], _26133_, _22731_);
  and _30807_ (_26135_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _30808_ (_26136_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _30809_ (_26137_, _22740_, _26136_);
  or _30810_ (_26138_, _26137_, _26135_);
  and _30811_ (_26862_[7], _26138_, _22731_);
  and _30812_ (_26139_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _30813_ (_26140_, _22740_, _22772_);
  or _30814_ (_26141_, _26140_, _26139_);
  and _30815_ (_26862_[6], _26141_, _22731_);
  and _30816_ (_26142_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _30817_ (_26143_, _22740_, _22767_);
  or _30818_ (_26144_, _26143_, _26142_);
  and _30819_ (_26862_[5], _26144_, _22731_);
  and _30820_ (_26145_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _30821_ (_26146_, _22740_, _22762_);
  or _30822_ (_26147_, _26146_, _26145_);
  and _30823_ (_26862_[4], _26147_, _22731_);
  and _30824_ (_26148_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _30825_ (_26149_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _30826_ (_26150_, _22740_, _26149_);
  or _30827_ (_26151_, _26150_, _26148_);
  and _30828_ (_26862_[3], _26151_, _22731_);
  and _30829_ (_26152_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _30830_ (_26153_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _30831_ (_26154_, _22740_, _26153_);
  or _30832_ (_26155_, _26154_, _26152_);
  and _30833_ (_26862_[2], _26155_, _22731_);
  nor _30834_ (_26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _30835_ (_26157_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and _30836_ (_26158_, _26156_, _23296_);
  nor _30837_ (_26159_, _26158_, _26157_);
  not _30838_ (_26160_, _26159_);
  and _30839_ (_26161_, _23301_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _30840_ (_26162_, _26161_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _30841_ (_26163_, _23086_, _23049_);
  nor _30842_ (_26164_, _26163_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _30843_ (_26165_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _30844_ (_26166_, _23237_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _30845_ (_26167_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30846_ (_26168_, _23156_, _26167_);
  nand _30847_ (_26169_, _26168_, _26166_);
  or _30848_ (_26170_, _23156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30849_ (_26171_, _23084_, _26167_);
  nand _30850_ (_26172_, _26171_, _26170_);
  and _30851_ (_26173_, _26172_, _26169_);
  or _30852_ (_26174_, _23371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30853_ (_26175_, _23122_, _26167_);
  nand _30854_ (_26176_, _26175_, _26174_);
  or _30855_ (_26177_, _23122_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _30856_ (_26178_, _23049_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _30857_ (_26180_, _26178_, _26177_);
  and _30858_ (_26181_, _26180_, _26176_);
  nand _30859_ (_26182_, _26181_, _26173_);
  and _30860_ (_26183_, _26182_, _26165_);
  nor _30861_ (_26184_, _26183_, _26164_);
  or _30862_ (_26185_, _23269_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30863_ (_26186_, _23371_, _26167_);
  nand _30864_ (_26187_, _26186_, _26185_);
  and _30865_ (_26188_, _26187_, _26165_);
  and _30866_ (_26189_, _26180_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _30867_ (_26190_, _26189_, _26188_);
  not _30868_ (_26191_, _26190_);
  nand _30869_ (_26192_, _26156_, _23039_);
  nor _30870_ (_26193_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _30871_ (_26194_, _26193_);
  and _30872_ (_26195_, _26194_, _26192_);
  not _30873_ (_26196_, _26195_);
  or _30874_ (_26197_, _23301_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30875_ (_26198_, _23237_, _26167_);
  and _30876_ (_26199_, _26198_, _26197_);
  or _30877_ (_26200_, _26199_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _30878_ (_26201_, _26172_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _30879_ (_26202_, _26201_, _26200_);
  or _30880_ (_26203_, _26202_, _26196_);
  and _30881_ (_26204_, _23269_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30882_ (_26205_, _26204_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _30883_ (_26206_, _26176_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _30884_ (_26207_, _26206_, _26205_);
  nand _30885_ (_26208_, _26156_, _23079_);
  nor _30886_ (_26209_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _30887_ (_26210_, _26209_);
  and _30888_ (_26211_, _26210_, _26208_);
  not _30889_ (_26212_, _26211_);
  or _30890_ (_26213_, _26212_, _26207_);
  nand _30891_ (_26214_, _26201_, _26200_);
  or _30892_ (_26215_, _26214_, _26195_);
  and _30893_ (_26216_, _26215_, _26203_);
  not _30894_ (_26217_, _26216_);
  or _30895_ (_26218_, _26217_, _26213_);
  and _30896_ (_26219_, _26218_, _26203_);
  nand _30897_ (_26220_, _26206_, _26205_);
  or _30898_ (_26221_, _26211_, _26220_);
  and _30899_ (_26222_, _26221_, _26213_);
  and _30900_ (_26223_, _26222_, _26216_);
  not _30901_ (_26224_, _26156_);
  or _30902_ (_26225_, _26224_, _23115_);
  nor _30903_ (_26226_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _30904_ (_26227_, _26226_);
  and _30905_ (_26228_, _26227_, _26225_);
  or _30906_ (_26229_, _26161_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _30907_ (_26230_, _26169_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _30908_ (_26231_, _26230_, _26229_);
  nand _30909_ (_26232_, _26231_, _26228_);
  or _30910_ (_26233_, _26231_, _26228_);
  nand _30911_ (_26234_, _26233_, _26232_);
  nor _30912_ (_26235_, _26187_, _26165_);
  nand _30913_ (_26236_, _26156_, _23150_);
  nor _30914_ (_26237_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _30915_ (_26238_, _26237_);
  and _30916_ (_26239_, _26238_, _26236_);
  not _30917_ (_26240_, _26239_);
  or _30918_ (_26241_, _26240_, _26235_);
  or _30919_ (_26242_, _26241_, _26234_);
  nand _30920_ (_26243_, _26242_, _26232_);
  nand _30921_ (_26244_, _26243_, _26223_);
  and _30922_ (_26245_, _26244_, _26219_);
  and _30923_ (_26246_, _26199_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _30924_ (_26247_, _26246_);
  nor _30925_ (_26248_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _30926_ (_26249_, _26248_);
  nand _30927_ (_26250_, _26156_, _23199_);
  and _30928_ (_26251_, _26250_, _26249_);
  nand _30929_ (_26252_, _26251_, _26247_);
  or _30930_ (_26253_, _26251_, _26247_);
  nand _30931_ (_26254_, _26253_, _26252_);
  nand _30932_ (_26255_, _26204_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _30933_ (_26256_, _26224_, _23232_);
  nor _30934_ (_26257_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _30935_ (_26258_, _26257_);
  and _30936_ (_26259_, _26258_, _26256_);
  nand _30937_ (_26260_, _26259_, _26255_);
  or _30938_ (_26261_, _26224_, _23264_);
  nor _30939_ (_26262_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _30940_ (_26263_, _26262_);
  nand _30941_ (_26264_, _26263_, _26261_);
  and _30942_ (_26265_, _26264_, _26162_);
  or _30943_ (_26266_, _26259_, _26255_);
  nand _30944_ (_26267_, _26266_, _26260_);
  or _30945_ (_26268_, _26267_, _26265_);
  and _30946_ (_26269_, _26268_, _26260_);
  or _30947_ (_26271_, _26269_, _26254_);
  nand _30948_ (_26272_, _26271_, _26252_);
  and _30949_ (_26273_, _26233_, _26232_);
  not _30950_ (_26274_, _26235_);
  or _30951_ (_26275_, _26239_, _26274_);
  and _30952_ (_26276_, _26275_, _26241_);
  and _30953_ (_26277_, _26276_, _26273_);
  and _30954_ (_26278_, _26277_, _26223_);
  nand _30955_ (_26279_, _26278_, _26272_);
  nand _30956_ (_26280_, _26279_, _26245_);
  and _30957_ (_26281_, _26191_, _26184_);
  nand _30958_ (_26282_, _26281_, _26280_);
  and _30959_ (_26283_, _26282_, _26195_);
  not _30960_ (_26284_, _26283_);
  and _30961_ (_26285_, _26281_, _26280_);
  and _30962_ (_26286_, _26276_, _26272_);
  not _30963_ (_26287_, _26286_);
  and _30964_ (_26288_, _26287_, _26241_);
  or _30965_ (_26289_, _26288_, _26234_);
  and _30966_ (_26290_, _26289_, _26232_);
  not _30967_ (_26291_, _26290_);
  nand _30968_ (_26292_, _26291_, _26222_);
  and _30969_ (_26293_, _26292_, _26213_);
  nand _30970_ (_26294_, _26293_, _26216_);
  or _30971_ (_26295_, _26293_, _26216_);
  nand _30972_ (_26296_, _26295_, _26294_);
  nand _30973_ (_26297_, _26296_, _26285_);
  nand _30974_ (_26298_, _26297_, _26284_);
  or _30975_ (_26299_, _26298_, _26191_);
  nand _30976_ (_26300_, _26298_, _26191_);
  or _30977_ (_26301_, _26291_, _26222_);
  nand _30978_ (_26302_, _26301_, _26292_);
  nand _30979_ (_26303_, _26302_, _26285_);
  and _30980_ (_26304_, _26282_, _26212_);
  not _30981_ (_26305_, _26304_);
  and _30982_ (_26306_, _26305_, _26303_);
  and _30983_ (_26307_, _26306_, _26214_);
  not _30984_ (_26308_, _26307_);
  nand _30985_ (_26309_, _26308_, _26300_);
  nand _30986_ (_26310_, _26309_, _26299_);
  and _30987_ (_26311_, _26300_, _26299_);
  nor _30988_ (_26312_, _26306_, _26214_);
  nor _30989_ (_26313_, _26312_, _26307_);
  and _30990_ (_26314_, _26313_, _26311_);
  nand _30991_ (_26315_, _26288_, _26234_);
  nand _30992_ (_26316_, _26315_, _26289_);
  nand _30993_ (_26317_, _26316_, _26285_);
  nor _30994_ (_26318_, _26285_, _26228_);
  not _30995_ (_26319_, _26318_);
  and _30996_ (_26320_, _26319_, _26317_);
  and _30997_ (_26321_, _26320_, _26220_);
  nor _30998_ (_26322_, _26276_, _26272_);
  nor _30999_ (_26323_, _26322_, _26286_);
  nor _31000_ (_26324_, _26323_, _26282_);
  and _31001_ (_26325_, _26282_, _26240_);
  nor _31002_ (_26326_, _26325_, _26324_);
  and _31003_ (_26327_, _26326_, _26231_);
  not _31004_ (_26328_, _26327_);
  nor _31005_ (_26329_, _26320_, _26220_);
  or _31006_ (_26330_, _26321_, _26329_);
  nor _31007_ (_26331_, _26330_, _26328_);
  or _31008_ (_26332_, _26331_, _26321_);
  and _31009_ (_26333_, _26269_, _26254_);
  not _31010_ (_26334_, _26333_);
  and _31011_ (_26335_, _26334_, _26271_);
  or _31012_ (_26336_, _26335_, _26282_);
  or _31013_ (_26337_, _26285_, _26251_);
  and _31014_ (_26338_, _26337_, _26336_);
  nor _31015_ (_26339_, _26338_, _26274_);
  not _31016_ (_26340_, _26339_);
  not _31017_ (_26341_, _26162_);
  or _31018_ (_26342_, _26282_, _26341_);
  nand _31019_ (_26343_, _26342_, _26264_);
  or _31020_ (_26344_, _26342_, _26264_);
  and _31021_ (_26345_, _26344_, _26343_);
  nand _31022_ (_26346_, _26345_, _26255_);
  or _31023_ (_26347_, _26345_, _26255_);
  and _31024_ (_26348_, _26347_, _26346_);
  nor _31025_ (_26349_, _26341_, _26159_);
  not _31026_ (_26350_, _26349_);
  nand _31027_ (_26351_, _26350_, _26348_);
  and _31028_ (_26352_, _26351_, _26346_);
  and _31029_ (_26353_, _26267_, _26265_);
  not _31030_ (_26354_, _26353_);
  and _31031_ (_26355_, _26354_, _26268_);
  or _31032_ (_26356_, _26355_, _26282_);
  or _31033_ (_26357_, _26285_, _26259_);
  and _31034_ (_26358_, _26357_, _26356_);
  nand _31035_ (_26359_, _26358_, _26247_);
  or _31036_ (_26360_, _26358_, _26247_);
  and _31037_ (_26361_, _26360_, _26359_);
  not _31038_ (_26362_, _26361_);
  or _31039_ (_26363_, _26362_, _26352_);
  and _31040_ (_26364_, _26338_, _26274_);
  not _31041_ (_26365_, _26364_);
  and _31042_ (_26366_, _26365_, _26359_);
  nand _31043_ (_26367_, _26366_, _26363_);
  and _31044_ (_26368_, _26367_, _26340_);
  nor _31045_ (_26369_, _26326_, _26231_);
  nor _31046_ (_26370_, _26369_, _26327_);
  not _31047_ (_26371_, _26330_);
  and _31048_ (_26372_, _26371_, _26370_);
  and _31049_ (_26373_, _26372_, _26368_);
  or _31050_ (_26374_, _26373_, _26332_);
  nand _31051_ (_26375_, _26374_, _26314_);
  nand _31052_ (_26376_, _26375_, _26310_);
  and _31053_ (_26377_, _26376_, _26184_);
  and _31054_ (_26378_, _26377_, _26162_);
  nor _31055_ (_26379_, _26378_, _26160_);
  and _31056_ (_26380_, _26378_, _26160_);
  or _31057_ (_26381_, _26380_, _26379_);
  nand _31058_ (_26382_, _26381_, _23528_);
  and _31059_ (_26383_, _23364_, _23403_);
  nor _31060_ (_26384_, _26383_, _23404_);
  nand _31061_ (_26385_, _23390_, _26384_);
  and _31062_ (_26386_, _23477_, _23487_);
  nor _31063_ (_26387_, _23484_, _23461_);
  nor _31064_ (_26388_, _26387_, _23296_);
  nor _31065_ (_26389_, _26388_, _26386_);
  and _31066_ (_26390_, _26389_, _24197_);
  and _31067_ (_26391_, _26390_, _24201_);
  and _31068_ (_26392_, _26391_, _26385_);
  nor _31069_ (_26393_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _31070_ (_26394_, _26393_);
  and _31071_ (_26395_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand _31072_ (_26396_, _26393_, _23049_);
  not _31073_ (_26397_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _31074_ (_26398_, _26397_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _31075_ (_26399_, _26398_);
  or _31076_ (_26400_, _26399_, _23120_);
  not _31077_ (_26401_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _31078_ (_26402_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _26401_);
  not _31079_ (_26403_, _26402_);
  or _31080_ (_26404_, _26403_, _23205_);
  and _31081_ (_26405_, _26404_, _26400_);
  nor _31082_ (_26406_, _26402_, _26398_);
  or _31083_ (_26407_, _23269_, _26401_);
  nand _31084_ (_26408_, _26407_, _26406_);
  nand _31085_ (_26409_, _26408_, _26405_);
  and _31086_ (_26410_, _26409_, _26396_);
  and _31087_ (_26411_, _26410_, _23264_);
  or _31088_ (_26412_, _26394_, _23084_);
  or _31089_ (_26413_, _26399_, _23169_);
  or _31090_ (_26414_, _26403_, _23310_);
  and _31091_ (_26415_, _26414_, _26413_);
  or _31092_ (_26416_, _23301_, _26401_);
  nand _31093_ (_26417_, _26416_, _26406_);
  nand _31094_ (_26418_, _26417_, _26415_);
  and _31095_ (_26419_, _26418_, _26412_);
  and _31096_ (_26420_, _26419_, _23232_);
  nand _31097_ (_26421_, _26420_, _26411_);
  and _31098_ (_26422_, _26419_, _23563_);
  nand _31099_ (_26423_, _26418_, _26412_);
  or _31100_ (_26424_, _26423_, _23509_);
  and _31101_ (_26425_, _26410_, _23232_);
  and _31102_ (_26426_, _26425_, _26424_);
  nand _31103_ (_26427_, _26426_, _26422_);
  nand _31104_ (_26428_, _26427_, _26421_);
  nand _31105_ (_26429_, _26409_, _26396_);
  or _31106_ (_26430_, _26429_, _23199_);
  or _31107_ (_26431_, _26423_, _23150_);
  or _31108_ (_26432_, _26431_, _26430_);
  nand _31109_ (_26433_, _26431_, _26430_);
  and _31110_ (_26434_, _26433_, _26432_);
  and _31111_ (_26435_, _26434_, _26428_);
  and _31112_ (_26436_, _26410_, _23460_);
  and _31113_ (_26437_, _26436_, _26422_);
  or _31114_ (_26438_, _26429_, _23457_);
  or _31115_ (_26439_, _26438_, _26431_);
  and _31116_ (_26440_, _26419_, _23115_);
  or _31117_ (_26441_, _26440_, _26436_);
  and _31118_ (_26442_, _26441_, _26439_);
  nand _31119_ (_26443_, _26442_, _26437_);
  or _31120_ (_26444_, _26442_, _26437_);
  and _31121_ (_26445_, _26444_, _26443_);
  nand _31122_ (_26446_, _26445_, _26435_);
  not _31123_ (_26447_, _26438_);
  or _31124_ (_26448_, _26439_, _23079_);
  and _31125_ (_26449_, _26419_, _23959_);
  not _31126_ (_26450_, _26449_);
  nand _31127_ (_26451_, _26450_, _26439_);
  and _31128_ (_26452_, _26451_, _26448_);
  nand _31129_ (_26453_, _26452_, _26447_);
  or _31130_ (_26454_, _26449_, _26447_);
  nand _31131_ (_26455_, _26454_, _26453_);
  or _31132_ (_26456_, _26455_, _26446_);
  and _31133_ (_26457_, _26419_, _23491_);
  and _31134_ (_26458_, _26457_, _26411_);
  or _31135_ (_26459_, _26420_, _26411_);
  and _31136_ (_26460_, _26459_, _26421_);
  and _31137_ (_26461_, _26460_, _26458_);
  or _31138_ (_26462_, _26426_, _26422_);
  and _31139_ (_26463_, _26462_, _26427_);
  nand _31140_ (_26464_, _26463_, _26461_);
  not _31141_ (_26465_, _26464_);
  nand _31142_ (_26466_, _26434_, _26428_);
  or _31143_ (_26467_, _26434_, _26428_);
  and _31144_ (_26468_, _26467_, _26466_);
  nand _31145_ (_26469_, _26468_, _26465_);
  or _31146_ (_26470_, _26445_, _26435_);
  nand _31147_ (_26471_, _26470_, _26446_);
  or _31148_ (_26472_, _26471_, _26469_);
  and _31149_ (_26473_, _26446_, _26443_);
  nand _31150_ (_26474_, _26473_, _26455_);
  or _31151_ (_26475_, _26473_, _26455_);
  nand _31152_ (_26476_, _26475_, _26474_);
  or _31153_ (_26477_, _26476_, _26472_);
  and _31154_ (_26478_, _26477_, _26456_);
  nor _31155_ (_26479_, _26455_, _26443_);
  not _31156_ (_26480_, _26448_);
  and _31157_ (_26481_, _26452_, _26447_);
  or _31158_ (_26482_, _26423_, _23039_);
  or _31159_ (_26483_, _26429_, _23079_);
  or _31160_ (_26484_, _26483_, _26482_);
  nand _31161_ (_26485_, _26483_, _26482_);
  and _31162_ (_26486_, _26485_, _26484_);
  nand _31163_ (_26487_, _26486_, _26481_);
  or _31164_ (_26488_, _26486_, _26481_);
  and _31165_ (_26489_, _26488_, _26487_);
  nand _31166_ (_26490_, _26489_, _26480_);
  or _31167_ (_26491_, _26489_, _26480_);
  and _31168_ (_26492_, _26491_, _26490_);
  nand _31169_ (_26493_, _26492_, _26479_);
  or _31170_ (_26494_, _26492_, _26479_);
  nand _31171_ (_26495_, _26494_, _26493_);
  or _31172_ (_26496_, _26495_, _26478_);
  nand _31173_ (_26497_, _26495_, _26478_);
  and _31174_ (_26498_, _26497_, _26496_);
  nand _31175_ (_26499_, _26498_, _26395_);
  or _31176_ (_26500_, _26498_, _26395_);
  and _31177_ (_26501_, _26500_, _26499_);
  and _31178_ (_26502_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nand _31179_ (_26503_, _26476_, _26472_);
  and _31180_ (_26504_, _26503_, _26477_);
  nand _31181_ (_26505_, _26504_, _26502_);
  or _31182_ (_26506_, _26504_, _26502_);
  nand _31183_ (_26507_, _26506_, _26505_);
  and _31184_ (_26508_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nand _31185_ (_26509_, _26471_, _26469_);
  and _31186_ (_26510_, _26509_, _26472_);
  nand _31187_ (_26511_, _26510_, _26508_);
  or _31188_ (_26512_, _26510_, _26508_);
  nand _31189_ (_26513_, _26512_, _26511_);
  and _31190_ (_26514_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or _31191_ (_26515_, _26468_, _26465_);
  and _31192_ (_26516_, _26515_, _26469_);
  nand _31193_ (_26517_, _26516_, _26514_);
  and _31194_ (_26518_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or _31195_ (_26519_, _26463_, _26461_);
  and _31196_ (_26520_, _26519_, _26464_);
  nand _31197_ (_26521_, _26520_, _26518_);
  and _31198_ (_26522_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand _31199_ (_26523_, _26460_, _26458_);
  or _31200_ (_26524_, _26460_, _26458_);
  and _31201_ (_26525_, _26524_, _26523_);
  and _31202_ (_26526_, _26525_, _26522_);
  not _31203_ (_26527_, _26526_);
  or _31204_ (_26528_, _26520_, _26518_);
  nand _31205_ (_26529_, _26528_, _26521_);
  or _31206_ (_26530_, _26529_, _26527_);
  and _31207_ (_26531_, _26530_, _26521_);
  or _31208_ (_26532_, _26516_, _26514_);
  nand _31209_ (_26533_, _26532_, _26517_);
  or _31210_ (_26534_, _26533_, _26531_);
  and _31211_ (_26535_, _26534_, _26517_);
  or _31212_ (_26536_, _26535_, _26513_);
  and _31213_ (_26537_, _26536_, _26511_);
  or _31214_ (_26538_, _26537_, _26507_);
  nand _31215_ (_26539_, _26538_, _26505_);
  nand _31216_ (_26540_, _26539_, _26501_);
  nand _31217_ (_26541_, _26540_, _26499_);
  and _31218_ (_26542_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  nand _31219_ (_26543_, _26496_, _26493_);
  and _31220_ (_26544_, _26410_, _23487_);
  and _31221_ (_26545_, _26544_, _26450_);
  and _31222_ (_26546_, _26490_, _26487_);
  not _31223_ (_26547_, _26546_);
  nand _31224_ (_26548_, _26547_, _26545_);
  or _31225_ (_26549_, _26547_, _26545_);
  and _31226_ (_26550_, _26549_, _26548_);
  nand _31227_ (_26551_, _26550_, _26543_);
  or _31228_ (_26552_, _26550_, _26543_);
  and _31229_ (_26553_, _26552_, _26551_);
  nand _31230_ (_26554_, _26553_, _26542_);
  or _31231_ (_26555_, _26553_, _26542_);
  nand _31232_ (_26556_, _26555_, _26554_);
  not _31233_ (_26557_, _26556_);
  and _31234_ (_26558_, _26557_, _26541_);
  nor _31235_ (_26559_, _26557_, _26541_);
  nor _31236_ (_26560_, _26559_, _26558_);
  and _31237_ (_26561_, _26560_, _23531_);
  and _31238_ (_26562_, _26384_, _22995_);
  and _31239_ (_26563_, _23488_, _23456_);
  nand _31240_ (_26564_, _23534_, _23264_);
  nand _31241_ (_26565_, _24206_, _26564_);
  or _31242_ (_26566_, _26565_, _26563_);
  or _31243_ (_26567_, _26566_, _26562_);
  nor _31244_ (_26568_, _26567_, _26561_);
  and _31245_ (_26569_, _26568_, _26392_);
  nand _31246_ (_26570_, _26569_, _26382_);
  not _31247_ (_26571_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _31248_ (_26572_, \oc8051_top_1.oc8051_decoder1.state [1], _22735_);
  and _31249_ (_26573_, _26572_, _26571_);
  and _31250_ (_26574_, _24251_, _26573_);
  not _31251_ (_26575_, _26573_);
  and _31252_ (_26576_, _23816_, _23772_);
  nor _31253_ (_26577_, _26576_, _24251_);
  and _31254_ (_26578_, _23825_, _23805_);
  or _31255_ (_26579_, _23898_, _23807_);
  nor _31256_ (_26580_, _26579_, _26578_);
  and _31257_ (_26581_, _23818_, _23816_);
  and _31258_ (_26582_, _23903_, _23816_);
  nor _31259_ (_26583_, _26582_, _26581_);
  and _31260_ (_26584_, _23816_, _23810_);
  nor _31261_ (_26585_, _26584_, _23897_);
  and _31262_ (_26586_, _26585_, _26583_);
  and _31263_ (_26587_, _26586_, _26580_);
  and _31264_ (_26588_, _26587_, _26577_);
  nor _31265_ (_26589_, _26588_, _26575_);
  and _31266_ (_26590_, _23816_, _24278_);
  and _31267_ (_26591_, _26590_, _23903_);
  nor _31268_ (_26592_, _26591_, _26589_);
  and _31269_ (_26593_, _23802_, _23778_);
  and _31270_ (_26594_, _23800_, _23792_);
  nor _31271_ (_26595_, _26594_, _26593_);
  nor _31272_ (_26596_, _26595_, _24279_);
  nor _31273_ (_26597_, _26574_, _26596_);
  or _31274_ (_26598_, _26579_, _23897_);
  nand _31275_ (_26599_, _26598_, _26573_);
  or _31276_ (_26600_, _26583_, _26575_);
  and _31277_ (_26601_, \oc8051_top_1.oc8051_decoder1.state [0], _22735_);
  and _31278_ (_26602_, _26601_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _31279_ (_26603_, _23903_, _23792_);
  and _31280_ (_26605_, _26603_, _26602_);
  and _31281_ (_26606_, _26594_, _24278_);
  nor _31282_ (_26607_, _26606_, _26605_);
  not _31283_ (_26608_, _26591_);
  and _31284_ (_26609_, _26608_, _26607_);
  and _31285_ (_26610_, _26609_, _26600_);
  and _31286_ (_26611_, _26610_, _26599_);
  and _31287_ (_26612_, _26611_, _26597_);
  and _31288_ (_26613_, _26612_, _26592_);
  or _31289_ (_26614_, _26613_, _26574_);
  and _31290_ (_26615_, _26614_, _26570_);
  nor _31291_ (_26616_, _22737_, _23280_);
  and _31292_ (_26617_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _31293_ (_26618_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _31294_ (_26619_, _26618_, _26617_);
  and _31295_ (_26620_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _31296_ (_26622_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _31297_ (_26623_, _26622_, _26620_);
  and _31298_ (_26624_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _31299_ (_26625_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _31300_ (_26626_, _26625_, _26624_);
  and _31301_ (_26627_, _26626_, _26623_);
  and _31302_ (_26628_, _26627_, _26619_);
  nor _31303_ (_26629_, _26628_, _24471_);
  nor _31304_ (_26630_, _26629_, _26616_);
  not _31305_ (_26631_, _26630_);
  nand _31306_ (_26632_, _26582_, _24278_);
  and _31307_ (_26633_, _26632_, _26600_);
  and _31308_ (_26634_, _26607_, _26599_);
  nand _31309_ (_26635_, _26634_, _26633_);
  or _31310_ (_26636_, _26635_, _26631_);
  and _31311_ (_26637_, _26634_, _26633_);
  nor _31312_ (_26638_, _22737_, _23278_);
  or _31313_ (_26639_, _23623_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _31314_ (_26640_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _31315_ (_26641_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _31316_ (_26642_, _26641_, _26640_);
  and _31317_ (_26643_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _31318_ (_26644_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _31319_ (_26645_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _31320_ (_26646_, _26645_, _26644_);
  or _31321_ (_26647_, _26646_, _26643_);
  or _31322_ (_26648_, _26647_, _26642_);
  and _31323_ (_26649_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _31324_ (_26650_, _26649_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _31325_ (_26651_, _26650_, _26648_);
  and _31326_ (_26652_, _26651_, _22737_);
  and _31327_ (_26653_, _26652_, _26639_);
  nor _31328_ (_26654_, _26653_, _26638_);
  not _31329_ (_26655_, _26654_);
  or _31330_ (_26656_, _26655_, _26637_);
  and _31331_ (_26657_, _26656_, _26636_);
  and _31332_ (_26658_, _26657_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _31333_ (_26659_, _26657_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _31334_ (_26660_, _26635_, _26597_);
  nor _31335_ (_26662_, _26660_, _26592_);
  nand _31336_ (_26663_, _26662_, _26659_);
  nor _31337_ (_26664_, _26663_, _26658_);
  and _31338_ (_26665_, _26660_, _26592_);
  and _31339_ (_26666_, _26665_, _26631_);
  and _31340_ (_26667_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _31341_ (_26668_, _26667_, _26666_);
  or _31342_ (_26669_, _26668_, _26664_);
  or _31343_ (_26670_, _26669_, _26615_);
  nor _31344_ (_26671_, _26583_, _26601_);
  and _31345_ (_26672_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _31346_ (_26673_, _23911_, _23780_);
  nor _31347_ (_26674_, _24255_, _26673_);
  nor _31348_ (_26675_, _24244_, _23773_);
  and _31349_ (_26676_, _26675_, _26674_);
  nor _31350_ (_26677_, _26676_, _24279_);
  and _31351_ (_26678_, _26584_, _26573_);
  not _31352_ (_26679_, _22736_);
  nor _31353_ (_26680_, _26675_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _31354_ (_26681_, _26680_, _26679_);
  nor _31355_ (_26682_, _26681_, _26678_);
  not _31356_ (_26683_, _26682_);
  nor _31357_ (_26684_, _26683_, _26677_);
  nor _31358_ (_26686_, _26684_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _31359_ (_26687_, _26686_, _26672_);
  and _31360_ (_26688_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _31361_ (_26689_, _26688_);
  and _31362_ (_26690_, _23816_, _23806_);
  and _31363_ (_26691_, _23814_, _23772_);
  nor _31364_ (_26692_, _26691_, _26690_);
  and _31365_ (_26693_, _23788_, _23708_);
  and _31366_ (_26694_, _26693_, _23814_);
  nor _31367_ (_26695_, _26694_, _26603_);
  and _31368_ (_26696_, _26695_, _26692_);
  nor _31369_ (_26697_, _23910_, _23841_);
  and _31370_ (_26698_, _23810_, _23708_);
  nand _31371_ (_26699_, _26698_, _23814_);
  and _31372_ (_26700_, _26699_, _26697_);
  and _31373_ (_26701_, _23814_, _23784_);
  nor _31374_ (_26702_, _26701_, _23840_);
  not _31375_ (_26703_, _26702_);
  nor _31376_ (_26704_, _26703_, _24269_);
  and _31377_ (_26705_, _26704_, _26700_);
  and _31378_ (_26706_, _26705_, _26696_);
  nand _31379_ (_26707_, _26706_, _26674_);
  nand _31380_ (_26708_, _26707_, _24278_);
  and _31381_ (_26709_, _26678_, _23769_);
  nor _31382_ (_26710_, _26709_, _26671_);
  and _31383_ (_26711_, _26710_, _26678_);
  nor _31384_ (_26712_, _26711_, _26605_);
  nand _31385_ (_26713_, _26712_, _26708_);
  nand _31386_ (_26714_, _26713_, _22735_);
  and _31387_ (_26715_, _26714_, _26689_);
  not _31388_ (_26716_, _26715_);
  and _31389_ (_26717_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _31390_ (_26718_, _26717_);
  nor _31391_ (_26719_, _24274_, _23930_);
  and _31392_ (_26720_, _26719_, _24260_);
  and _31393_ (_26721_, _23838_, _23783_);
  not _31394_ (_26722_, _26721_);
  and _31395_ (_26723_, _23801_, _23803_);
  and _31396_ (_26724_, _23803_, _23772_);
  nor _31397_ (_26726_, _26724_, _26723_);
  and _31398_ (_26727_, _26726_, _26722_);
  and _31399_ (_26729_, _26727_, _26720_);
  and _31400_ (_26730_, _23926_, _23708_);
  and _31401_ (_26731_, _26730_, _23797_);
  and _31402_ (_26732_, _26731_, _23685_);
  nor _31403_ (_26733_, _26732_, _23845_);
  and _31404_ (_26734_, _23911_, _23792_);
  and _31405_ (_26735_, _23923_, _23791_);
  nor _31406_ (_26736_, _26735_, _26734_);
  and _31407_ (_26737_, _26736_, _26733_);
  and _31408_ (_26738_, _26737_, _26729_);
  or _31409_ (_26739_, _23819_, _23807_);
  nand _31410_ (_26740_, _26739_, _23685_);
  not _31411_ (_26741_, _23817_);
  and _31412_ (_26742_, _23844_, _23792_);
  nor _31413_ (_26743_, _26742_, _23793_);
  and _31414_ (_26744_, _26743_, _26741_);
  and _31415_ (_26745_, _26744_, _26740_);
  not _31416_ (_26747_, _23803_);
  nor _31417_ (_26748_, _23903_, _23812_);
  nor _31418_ (_26749_, _26748_, _26747_);
  or _31419_ (_26750_, _23911_, _23784_);
  nand _31420_ (_26751_, _26750_, _23803_);
  nand _31421_ (_26752_, _26751_, _26583_);
  nor _31422_ (_26753_, _26752_, _26749_);
  and _31423_ (_26754_, _26693_, _23803_);
  nor _31424_ (_26755_, _26754_, _26603_);
  and _31425_ (_26756_, _23892_, _23814_);
  and _31426_ (_26757_, _26730_, _23779_);
  nor _31427_ (_26758_, _26757_, _26756_);
  and _31428_ (_26759_, _26758_, _26755_);
  and _31429_ (_26760_, _23816_, _23805_);
  nor _31430_ (_26761_, _26760_, _23893_);
  and _31431_ (_26762_, _26761_, _24265_);
  and _31432_ (_26763_, _26762_, _26759_);
  and _31433_ (_26764_, _26763_, _26753_);
  and _31434_ (_26765_, _26764_, _26745_);
  nand _31435_ (_26766_, _26765_, _26738_);
  nand _31436_ (_26767_, _26766_, _24278_);
  nor _31437_ (_26768_, _26605_, _26678_);
  nand _31438_ (_26769_, _26768_, _26767_);
  nand _31439_ (_26770_, _26769_, _22735_);
  and _31440_ (_26772_, _26770_, _26718_);
  and _31441_ (_26773_, _26772_, _26716_);
  and _31442_ (_26775_, _26773_, _26687_);
  nand _31443_ (_26776_, _26775_, _25954_);
  nor _31444_ (_26777_, _26772_, _26715_);
  and _31445_ (_26778_, _26777_, _26687_);
  and _31446_ (_26779_, _24177_, _22867_);
  and _31447_ (_26780_, _26779_, _24188_);
  and _31448_ (_26781_, _26780_, _23577_);
  and _31449_ (_26782_, _26780_, _23880_);
  not _31450_ (_26783_, _26780_);
  and _31451_ (_26784_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _31452_ (_26786_, _26784_, _26782_);
  and _31453_ (_26787_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _31454_ (_26788_, _26783_, _23542_);
  nor _31455_ (_26789_, _26788_, _26787_);
  nand _31456_ (_26790_, _26780_, _24671_);
  or _31457_ (_26791_, _26780_, _22874_);
  and _31458_ (_26792_, _26791_, _26790_);
  and _31459_ (_26793_, _26792_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _31460_ (_26794_, _26793_, _26789_);
  and _31461_ (_26795_, _26794_, _26786_);
  and _31462_ (_26796_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _31463_ (_26797_, _26796_, _26781_);
  and _31464_ (_26798_, _26797_, _26795_);
  nor _31465_ (_26799_, _26797_, _26795_);
  nor _31466_ (_26800_, _26799_, _26798_);
  nor _31467_ (_26801_, _26800_, _22815_);
  nor _31468_ (_26802_, _26801_, _22857_);
  nor _31469_ (_26803_, _26802_, _26780_);
  nor _31470_ (_26804_, _26803_, _26781_);
  not _31471_ (_26805_, _26804_);
  nand _31472_ (_26806_, _26805_, _26778_);
  and _31473_ (_26807_, _26715_, _26687_);
  and _31474_ (_26808_, _26807_, _26772_);
  nand _31475_ (_26809_, _26808_, _25687_);
  not _31476_ (_26810_, _24473_);
  not _31477_ (_26811_, _26772_);
  and _31478_ (_26812_, _26807_, _26811_);
  nand _31479_ (_26813_, _26812_, _26810_);
  and _31480_ (_26814_, _26813_, _26809_);
  and _31481_ (_26815_, _26814_, _26806_);
  and _31482_ (_26816_, _26815_, _26776_);
  nor _31483_ (_26818_, _26816_, _22867_);
  and _31484_ (_26819_, _26816_, _22867_);
  nor _31485_ (_26820_, _26819_, _26818_);
  not _31486_ (_26821_, _26820_);
  and _31487_ (_00001_, _26775_, _25976_);
  not _31488_ (_00002_, _00001_);
  not _31489_ (_00003_, _26778_);
  nor _31490_ (_00004_, _26783_, _24082_);
  and _31491_ (_00005_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _31492_ (_00006_, _00005_, _00004_);
  and _31493_ (_00008_, _00006_, _26798_);
  nor _31494_ (_00009_, _00006_, _26798_);
  nor _31495_ (_00010_, _00009_, _00008_);
  nor _31496_ (_00011_, _00010_, _22815_);
  nor _31497_ (_00012_, _00011_, _22896_);
  nor _31498_ (_00013_, _00012_, _26780_);
  nor _31499_ (_00014_, _00013_, _00004_);
  nor _31500_ (_00015_, _00014_, _00003_);
  and _31501_ (_00016_, _26808_, _25855_);
  not _31502_ (_00017_, _00016_);
  or _31503_ (_00018_, _26772_, _26716_);
  nor _31504_ (_00020_, _00018_, _25577_);
  not _31505_ (_00021_, _26687_);
  and _31506_ (_00023_, _26715_, _00021_);
  nor _31507_ (_00024_, _00023_, _00020_);
  nand _31508_ (_00025_, _00024_, _00017_);
  nor _31509_ (_00026_, _00025_, _00015_);
  and _31510_ (_00027_, _00026_, _00002_);
  nor _31511_ (_00028_, _00027_, _22905_);
  and _31512_ (_00029_, _00027_, _22905_);
  nor _31513_ (_00030_, _00029_, _00028_);
  and _31514_ (_00031_, _26775_, _25995_);
  not _31515_ (_00033_, _26050_);
  and _31516_ (_00034_, _26812_, _00033_);
  nor _31517_ (_00035_, _00034_, _00031_);
  nor _31518_ (_00036_, _26783_, _24043_);
  and _31519_ (_00037_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _31520_ (_00038_, _00037_, _00036_);
  and _31521_ (_00039_, _00038_, _00008_);
  nor _31522_ (_00040_, _00038_, _00008_);
  nor _31523_ (_00041_, _00040_, _00039_);
  nor _31524_ (_00042_, _00041_, _22815_);
  nor _31525_ (_00043_, _00042_, _22927_);
  nor _31526_ (_00045_, _00043_, _26780_);
  nor _31527_ (_00046_, _00045_, _00036_);
  nor _31528_ (_00047_, _00046_, _00003_);
  nor _31529_ (_00048_, _26773_, _26687_);
  and _31530_ (_00049_, _00048_, _00018_);
  nor _31531_ (_00050_, _00049_, _00047_);
  and _31532_ (_00051_, _00050_, _00035_);
  nor _31533_ (_00052_, _00051_, _22936_);
  and _31534_ (_00053_, _00051_, _22936_);
  nor _31535_ (_00054_, _00053_, _00052_);
  nor _31536_ (_00055_, _00054_, _00030_);
  nor _31537_ (_00056_, _22737_, _23062_);
  and _31538_ (_00057_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _31539_ (_00058_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _31540_ (_00059_, _00058_, _00057_);
  and _31541_ (_00060_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _31542_ (_00061_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _31543_ (_00062_, _00061_, _00060_);
  and _31544_ (_00063_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _31545_ (_00064_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _31546_ (_00065_, _00064_, _00063_);
  and _31547_ (_00066_, _00065_, _00062_);
  and _31548_ (_00067_, _00066_, _00059_);
  nor _31549_ (_00068_, _00067_, _24471_);
  nor _31550_ (_00069_, _00068_, _00056_);
  not _31551_ (_00070_, _00069_);
  and _31552_ (_00071_, _00070_, _26812_);
  nor _31553_ (_00072_, _26783_, _24126_);
  and _31554_ (_00073_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _31555_ (_00075_, _00073_, _00072_);
  and _31556_ (_00076_, _00075_, _00039_);
  nor _31557_ (_00077_, _00075_, _00039_);
  nor _31558_ (_00078_, _00077_, _00076_);
  nor _31559_ (_00080_, _00078_, _22815_);
  nor _31560_ (_00081_, _00080_, _22960_);
  nor _31561_ (_00083_, _00081_, _26780_);
  nor _31562_ (_00084_, _00083_, _00072_);
  nor _31563_ (_00085_, _00084_, _00003_);
  and _31564_ (_00086_, _26775_, _26018_);
  or _31565_ (_00088_, _00048_, _00086_);
  or _31566_ (_00089_, _00088_, _00085_);
  nor _31567_ (_00090_, _00089_, _00071_);
  nor _31568_ (_00091_, _00090_, _22968_);
  and _31569_ (_00092_, _00090_, _22968_);
  nor _31570_ (_00093_, _00092_, _00091_);
  and _31571_ (_00094_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand _31572_ (_00095_, _00094_, _00076_);
  or _31573_ (_00096_, _00094_, _00076_);
  and _31574_ (_00097_, _00096_, _22854_);
  nand _31575_ (_00098_, _00097_, _00095_);
  nor _31576_ (_00099_, _26780_, _22826_);
  nand _31577_ (_00100_, _00099_, _00098_);
  and _31578_ (_00101_, _26780_, _23989_);
  not _31579_ (_00102_, _00101_);
  nand _31580_ (_00104_, _00102_, _00100_);
  not _31581_ (_00105_, _00104_);
  nand _31582_ (_00106_, _00105_, _26777_);
  nand _31583_ (_00107_, _25852_, _23989_);
  nand _31584_ (_00108_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand _31585_ (_00109_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _31586_ (_00110_, _00109_, _00108_);
  nand _31587_ (_00111_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand _31588_ (_00112_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _31589_ (_00113_, _00112_, _00111_);
  and _31590_ (_00114_, _00113_, _00110_);
  nand _31591_ (_00115_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand _31592_ (_00116_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _31593_ (_00117_, _00116_, _00115_);
  nand _31594_ (_00118_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand _31595_ (_00119_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _31596_ (_00120_, _00119_, _00118_);
  and _31597_ (_00121_, _00120_, _00117_);
  and _31598_ (_00122_, _00121_, _25872_);
  nand _31599_ (_00123_, _00122_, _00114_);
  and _31600_ (_00124_, _00123_, _00107_);
  nand _31601_ (_00125_, _00124_, _26773_);
  nor _31602_ (_00126_, _22737_, _23008_);
  and _31603_ (_00127_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _31604_ (_00128_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _31605_ (_00129_, _00128_, _00127_);
  and _31606_ (_00130_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _31607_ (_00131_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _31608_ (_00132_, _00131_, _00130_);
  and _31609_ (_00133_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _31610_ (_00134_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _31611_ (_00135_, _00134_, _00133_);
  and _31612_ (_00136_, _00135_, _00132_);
  and _31613_ (_00137_, _00136_, _00129_);
  nor _31614_ (_00138_, _00137_, _24471_);
  nor _31615_ (_00139_, _00138_, _00126_);
  or _31616_ (_00140_, _00139_, _00018_);
  and _31617_ (_00141_, _00140_, _26687_);
  and _31618_ (_00142_, _00141_, _00125_);
  nand _31619_ (_00143_, _00142_, _00106_);
  and _31620_ (_00144_, _00143_, _22844_);
  nor _31621_ (_00145_, _00143_, _22844_);
  nor _31622_ (_00146_, _00145_, _00144_);
  nor _31623_ (_00147_, _00146_, _00093_);
  and _31624_ (_00148_, _00147_, _00055_);
  and _31625_ (_00149_, _00148_, _26821_);
  nor _31626_ (_00150_, _25481_, _24180_);
  and _31627_ (_00151_, _00150_, _00149_);
  and _31628_ (_00152_, _00151_, _26671_);
  not _31629_ (_00153_, _00152_);
  and _31630_ (_00154_, _26775_, _25911_);
  not _31631_ (_00155_, _00154_);
  and _31632_ (_00156_, _26808_, _23664_);
  not _31633_ (_00157_, _26068_);
  and _31634_ (_00158_, _26812_, _00157_);
  nor _31635_ (_00159_, _00158_, _00156_);
  and _31636_ (_00160_, _26773_, _00021_);
  nor _31637_ (_00161_, _26793_, _26789_);
  nor _31638_ (_00162_, _00161_, _26794_);
  nor _31639_ (_00163_, _00162_, _22815_);
  nor _31640_ (_00164_, _00163_, _22911_);
  nor _31641_ (_00165_, _00164_, _26780_);
  nor _31642_ (_00166_, _00165_, _26788_);
  not _31643_ (_00167_, _00166_);
  and _31644_ (_00168_, _00167_, _26778_);
  nor _31645_ (_00169_, _00168_, _00160_);
  and _31646_ (_00170_, _00169_, _00159_);
  and _31647_ (_00171_, _00170_, _00155_);
  nor _31648_ (_00173_, _00171_, _22919_);
  and _31649_ (_00174_, _00171_, _22919_);
  nor _31650_ (_00175_, _00174_, _00173_);
  or _31651_ (_00176_, _26820_, _25113_);
  and _31652_ (_00177_, _26775_, _25891_);
  and _31653_ (_00178_, _26631_, _26812_);
  nor _31654_ (_00179_, _00178_, _00177_);
  nor _31655_ (_00180_, _26792_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _31656_ (_00181_, _00180_, _26793_);
  nor _31657_ (_00182_, _00181_, _22815_);
  nor _31658_ (_00183_, _00182_, _22875_);
  nor _31659_ (_00185_, _00183_, _26780_);
  not _31660_ (_00186_, _00185_);
  and _31661_ (_00187_, _00186_, _26790_);
  nor _31662_ (_00188_, _00187_, _00003_);
  and _31663_ (_00189_, _26808_, _23685_);
  nor _31664_ (_00190_, _00189_, _00188_);
  and _31665_ (_00191_, _00190_, _00179_);
  and _31666_ (_00192_, _00191_, _24175_);
  nor _31667_ (_00193_, _00191_, _24175_);
  or _31668_ (_00194_, _00193_, _00192_);
  and _31669_ (_00195_, _26775_, _25930_);
  not _31670_ (_00196_, _00195_);
  and _31671_ (_00197_, _26808_, _23643_);
  nor _31672_ (_00198_, _26794_, _26786_);
  nor _31673_ (_00199_, _00198_, _26795_);
  nor _31674_ (_00200_, _00199_, _22815_);
  nor _31675_ (_00201_, _00200_, _22942_);
  nor _31676_ (_00202_, _00201_, _26780_);
  nor _31677_ (_00204_, _00202_, _26782_);
  not _31678_ (_00205_, _00204_);
  and _31679_ (_00206_, _00205_, _26778_);
  nor _31680_ (_00207_, _22737_, _23226_);
  and _31681_ (_00208_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _31682_ (_00210_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _31683_ (_00211_, _00210_, _00208_);
  and _31684_ (_00213_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _31685_ (_00214_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _31686_ (_00216_, _00214_, _00213_);
  and _31687_ (_00217_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _31688_ (_00218_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _31689_ (_00219_, _00218_, _00217_);
  and _31690_ (_00220_, _00219_, _00216_);
  and _31691_ (_00221_, _00220_, _00211_);
  nor _31692_ (_00222_, _00221_, _24471_);
  nor _31693_ (_00223_, _00222_, _00207_);
  not _31694_ (_00224_, _00223_);
  and _31695_ (_00225_, _00224_, _26812_);
  or _31696_ (_00226_, _00225_, _00206_);
  nor _31697_ (_00227_, _00226_, _00197_);
  and _31698_ (_00228_, _00227_, _00196_);
  nor _31699_ (_00229_, _00228_, _22951_);
  and _31700_ (_00230_, _00228_, _22951_);
  nor _31701_ (_00231_, _00230_, _00229_);
  or _31702_ (_00232_, _00231_, _00194_);
  or _31703_ (_00233_, _00232_, _00176_);
  nor _31704_ (_00234_, _00233_, _00175_);
  and _31705_ (_00235_, _00234_, _00148_);
  and _31706_ (_00236_, _22844_, _22869_);
  and _31707_ (_00237_, _00236_, _00235_);
  and _31708_ (_00238_, _26698_, _23816_);
  and _31709_ (_00239_, _26582_, _23708_);
  or _31710_ (_00240_, _00239_, _26581_);
  and _31711_ (_00241_, _23380_, _23393_);
  nor _31712_ (_00242_, _23380_, _23393_);
  nor _31713_ (_00243_, _00242_, _00241_);
  not _31714_ (_00244_, _00243_);
  nor _31715_ (_00245_, _23376_, _23173_);
  and _31716_ (_00246_, _23376_, _23173_);
  nor _31717_ (_00247_, _00246_, _00245_);
  and _31718_ (_00248_, _23369_, _23316_);
  nor _31719_ (_00249_, _00248_, _23370_);
  nor _31720_ (_00250_, _23367_, _23319_);
  nor _31721_ (_00251_, _00250_, _23368_);
  nor _31722_ (_00252_, _26678_, _23321_);
  and _31723_ (_00253_, _00252_, _00251_);
  nand _31724_ (_00254_, _00253_, _00249_);
  nor _31725_ (_00255_, _00254_, _00247_);
  not _31726_ (_00256_, _26384_);
  nor _31727_ (_00257_, _23377_, _23168_);
  nor _31728_ (_00258_, _00257_, _23378_);
  and _31729_ (_00259_, _00258_, _00256_);
  and _31730_ (_00260_, _00259_, _00255_);
  nor _31731_ (_00261_, _23378_, _23164_);
  nor _31732_ (_00263_, _00261_, _23379_);
  and _31733_ (_00264_, _00263_, _26710_);
  and _31734_ (_00265_, _00264_, _00260_);
  and _31735_ (_00266_, _00265_, _00244_);
  not _31736_ (_00267_, _00266_);
  and _31737_ (_00268_, _26709_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not _31738_ (_00269_, _00268_);
  and _31739_ (_00271_, _26671_, _23478_);
  nor _31740_ (_00272_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _31741_ (_00273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _31742_ (_00274_, _00273_, _00272_);
  nor _31743_ (_00275_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _31744_ (_00277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _31745_ (_00278_, _00277_, _00275_);
  and _31746_ (_00279_, _00278_, _00274_);
  and _31747_ (_00281_, _00279_, _26711_);
  nor _31748_ (_00282_, _00281_, _00271_);
  and _31749_ (_00283_, _00282_, _00269_);
  and _31750_ (_00284_, _00283_, _00267_);
  or _31751_ (_00285_, _00284_, _00240_);
  nor _31752_ (_00286_, _00285_, _00238_);
  and _31753_ (_00287_, _26582_, _23707_);
  not _31754_ (_00288_, _00287_);
  and _31755_ (_00290_, _26584_, _23707_);
  nor _31756_ (_00292_, _00290_, _23897_);
  and _31757_ (_00293_, _00292_, _00288_);
  and _31758_ (_00294_, _00293_, _26580_);
  and _31759_ (_00295_, _00294_, _00284_);
  nor _31760_ (_00296_, _00295_, _00286_);
  not _31761_ (_00297_, _26603_);
  and _31762_ (_00298_, _26577_, _00297_);
  not _31763_ (_00300_, _00298_);
  nor _31764_ (_00301_, _00300_, _00296_);
  nor _31765_ (_00303_, _26605_, _26573_);
  nor _31766_ (_00304_, _00303_, _00301_);
  nor _31767_ (_00306_, _00304_, _26596_);
  and _31768_ (_00307_, _25478_, _24539_);
  and _31769_ (_00308_, _00307_, _25017_);
  not _31770_ (_00309_, _00308_);
  nor _31771_ (_00311_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _31772_ (_00312_, _00311_);
  nor _31773_ (_00313_, _00312_, _25683_);
  and _31774_ (_00314_, _00313_, _00309_);
  not _31775_ (_00315_, _00314_);
  and _31776_ (_00316_, _00315_, _26709_);
  not _31777_ (_00317_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _31778_ (_00318_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _22735_);
  and _31779_ (_00319_, _00318_, _00317_);
  not _31780_ (_00320_, _00319_);
  nor _31781_ (_00321_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _31782_ (_00322_, _00321_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _31783_ (_00323_, _24625_, _24004_);
  and _31784_ (_00324_, _00323_, _25681_);
  nor _31785_ (_00325_, _00324_, _00322_);
  and _31786_ (_00326_, _00325_, _00320_);
  nor _31787_ (_00327_, _22968_, _22936_);
  and _31788_ (_00328_, _00327_, _24539_);
  and _31789_ (_00329_, _00328_, _25123_);
  not _31790_ (_00330_, _00329_);
  and _31791_ (_00331_, _00330_, _00326_);
  not _31792_ (_00332_, _00331_);
  and _31793_ (_00333_, _00332_, _26711_);
  nor _31794_ (_00334_, _00333_, _00316_);
  not _31795_ (_00335_, _00334_);
  nor _31796_ (_00336_, _00335_, _00306_);
  not _31797_ (_00337_, _00336_);
  nor _31798_ (_00338_, _00337_, _00237_);
  and _31799_ (_00339_, _00338_, _00153_);
  nand _31800_ (_00340_, _26655_, _26606_);
  nand _31801_ (_00341_, _00340_, _00339_);
  or _31802_ (_00342_, _00341_, _26670_);
  or _31803_ (_00343_, _00339_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _31804_ (_00344_, _00343_, _22731_);
  and _31805_ (_26870_[0], _00344_, _00342_);
  or _31806_ (_00345_, _00339_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _31807_ (_00346_, _00345_, _22731_);
  nand _31808_ (_00347_, _26376_, _26184_);
  or _31809_ (_00348_, _26350_, _26348_);
  and _31810_ (_00349_, _00348_, _26351_);
  or _31811_ (_00350_, _00349_, _00347_);
  or _31812_ (_00351_, _26377_, _26345_);
  and _31813_ (_00352_, _00351_, _00350_);
  nand _31814_ (_00353_, _00352_, _23528_);
  and _31815_ (_00354_, _26553_, _26542_);
  nor _31816_ (_00355_, _26558_, _00354_);
  and _31817_ (_00356_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and _31818_ (_00357_, _26548_, _26484_);
  nand _31819_ (_00358_, _00357_, _26551_);
  nand _31820_ (_00359_, _00358_, _00356_);
  or _31821_ (_00360_, _00358_, _00356_);
  nand _31822_ (_00361_, _00360_, _00359_);
  nand _31823_ (_00362_, _00361_, _00355_);
  or _31824_ (_00363_, _00361_, _00355_);
  and _31825_ (_00364_, _00363_, _00362_);
  nand _31826_ (_00365_, _00364_, _23531_);
  nor _31827_ (_00366_, _23463_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _31828_ (_00367_, _00366_, _23264_);
  nor _31829_ (_00368_, _00366_, _23264_);
  nor _31830_ (_00369_, _00368_, _00367_);
  nor _31831_ (_00370_, _00369_, _23470_);
  not _31832_ (_00371_, _00370_);
  nand _31833_ (_00372_, _23534_, _23232_);
  and _31834_ (_00373_, _23484_, _23264_);
  not _31835_ (_00374_, _23535_);
  nor _31836_ (_00375_, _00374_, _23296_);
  nor _31837_ (_00376_, _00375_, _00373_);
  and _31838_ (_00377_, _00376_, _00372_);
  and _31839_ (_00378_, _00377_, _23527_);
  and _31840_ (_00379_, _00378_, _00371_);
  and _31841_ (_00380_, _00379_, _23518_);
  nor _31842_ (_00381_, _23324_, _23272_);
  or _31843_ (_00382_, _00381_, _23396_);
  and _31844_ (_00383_, _00382_, _23404_);
  nor _31845_ (_00384_, _00382_, _23404_);
  or _31846_ (_00385_, _00384_, _00383_);
  and _31847_ (_00386_, _00385_, _23390_);
  nor _31848_ (_00387_, _23366_, _23322_);
  nor _31849_ (_00388_, _00387_, _23367_);
  nor _31850_ (_00389_, _00388_, _22996_);
  nor _31851_ (_00390_, _00389_, _00386_);
  and _31852_ (_00391_, _00390_, _00380_);
  and _31853_ (_00392_, _00391_, _00365_);
  nand _31854_ (_00393_, _00392_, _00353_);
  and _31855_ (_00394_, _00393_, _26614_);
  and _31856_ (_00395_, _26665_, _00157_);
  and _31857_ (_00396_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _31858_ (_00397_, _00396_, _00395_);
  or _31859_ (_00398_, _26635_, _00157_);
  nor _31860_ (_00399_, _22737_, _23246_);
  and _31861_ (_00400_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _31862_ (_00401_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _31863_ (_00402_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _31864_ (_00403_, _00402_, _00401_);
  and _31865_ (_00404_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _31866_ (_00405_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _31867_ (_00406_, _00405_, _00404_);
  or _31868_ (_00407_, _00406_, _00403_);
  and _31869_ (_00408_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _31870_ (_00409_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _31871_ (_00410_, _00409_, _00408_);
  or _31872_ (_00411_, _00410_, _00407_);
  and _31873_ (_00412_, _00411_, _23623_);
  or _31874_ (_00413_, _00412_, _00400_);
  and _31875_ (_00414_, _00413_, _22737_);
  nor _31876_ (_00415_, _00414_, _00399_);
  not _31877_ (_00416_, _00415_);
  or _31878_ (_00417_, _00416_, _26637_);
  and _31879_ (_00418_, _00417_, _00398_);
  nand _31880_ (_00419_, _00418_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _31881_ (_00420_, _00418_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _31882_ (_00421_, _00420_, _00419_);
  or _31883_ (_00422_, _00421_, _26658_);
  and _31884_ (_00423_, _00421_, _26658_);
  not _31885_ (_00424_, _00423_);
  and _31886_ (_00425_, _00424_, _26662_);
  and _31887_ (_00426_, _00425_, _00422_);
  or _31888_ (_00427_, _00426_, _00397_);
  or _31889_ (_00428_, _00427_, _00394_);
  nand _31890_ (_00429_, _00416_, _26606_);
  nand _31891_ (_00430_, _00429_, _00339_);
  or _31892_ (_00431_, _00430_, _00428_);
  and _31893_ (_26870_[1], _00431_, _00346_);
  not _31894_ (_00432_, _26363_);
  and _31895_ (_00433_, _26362_, _26352_);
  nor _31896_ (_00434_, _00433_, _00432_);
  or _31897_ (_00435_, _00434_, _00347_);
  or _31898_ (_00436_, _26377_, _26358_);
  and _31899_ (_00437_, _00436_, _00435_);
  nand _31900_ (_00438_, _00437_, _23528_);
  and _31901_ (_00439_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  not _31902_ (_00440_, _26541_);
  or _31903_ (_00441_, _00361_, _26556_);
  or _31904_ (_00442_, _00441_, _00440_);
  nand _31905_ (_00443_, _00360_, _00354_);
  and _31906_ (_00444_, _00443_, _00359_);
  and _31907_ (_00445_, _00444_, _00442_);
  not _31908_ (_00446_, _00445_);
  nand _31909_ (_00447_, _00446_, _00439_);
  or _31910_ (_00448_, _00446_, _00439_);
  and _31911_ (_00449_, _00448_, _00447_);
  nand _31912_ (_00450_, _00449_, _23531_);
  nor _31913_ (_00451_, _00251_, _22996_);
  and _31914_ (_00452_, _23484_, _23232_);
  not _31915_ (_00453_, _00452_);
  nand _31916_ (_00454_, _23535_, _23264_);
  not _31917_ (_00455_, _23534_);
  or _31918_ (_00456_, _00455_, _23199_);
  and _31919_ (_00457_, _00456_, _00454_);
  and _31920_ (_00458_, _00457_, _00453_);
  and _31921_ (_00459_, _00458_, _23876_);
  not _31922_ (_00460_, _00459_);
  nor _31923_ (_00461_, _00460_, _00451_);
  nor _31924_ (_00462_, _23407_, _23405_);
  nor _31925_ (_00463_, _00462_, _23391_);
  and _31926_ (_00464_, _00463_, _23409_);
  and _31927_ (_00465_, _23462_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _31928_ (_00466_, _00368_, _23872_);
  nor _31929_ (_00467_, _00466_, _00465_);
  nor _31930_ (_00468_, _00467_, _23470_);
  nor _31931_ (_00469_, _00468_, _00464_);
  and _31932_ (_00470_, _00469_, _00461_);
  and _31933_ (_00471_, _00470_, _23868_);
  and _31934_ (_00472_, _00471_, _00450_);
  nand _31935_ (_00473_, _00472_, _00438_);
  and _31936_ (_00474_, _00473_, _26614_);
  and _31937_ (_00475_, _26665_, _00224_);
  and _31938_ (_00476_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _31939_ (_00477_, _00476_, _00475_);
  nand _31940_ (_00478_, _00424_, _00419_);
  or _31941_ (_00479_, _26635_, _00224_);
  nor _31942_ (_00480_, _22737_, _23228_);
  and _31943_ (_00481_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _31944_ (_00482_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _31945_ (_00483_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _31946_ (_00484_, _00483_, _00482_);
  and _31947_ (_00485_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _31948_ (_00486_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _31949_ (_00487_, _00486_, _00485_);
  and _31950_ (_00488_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _31951_ (_00489_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _31952_ (_00490_, _00489_, _00488_);
  and _31953_ (_00491_, _00490_, _00487_);
  and _31954_ (_00492_, _00491_, _00484_);
  nor _31955_ (_00493_, _00492_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _31956_ (_00494_, _00493_, _00481_);
  nor _31957_ (_00495_, _00494_, _25454_);
  nor _31958_ (_00496_, _00495_, _00480_);
  not _31959_ (_00497_, _00496_);
  or _31960_ (_00498_, _00497_, _26637_);
  nand _31961_ (_00499_, _00498_, _00479_);
  or _31962_ (_00500_, _00499_, _23213_);
  nand _31963_ (_00501_, _00499_, _23213_);
  and _31964_ (_00502_, _00501_, _00500_);
  or _31965_ (_00503_, _00502_, _00478_);
  and _31966_ (_00504_, _00502_, _00478_);
  not _31967_ (_00505_, _00504_);
  and _31968_ (_00506_, _00505_, _26662_);
  and _31969_ (_00507_, _00506_, _00503_);
  or _31970_ (_00508_, _00507_, _00477_);
  or _31971_ (_00509_, _00508_, _00474_);
  nand _31972_ (_00510_, _00497_, _26606_);
  nand _31973_ (_00511_, _00510_, _00339_);
  or _31974_ (_00512_, _00511_, _00509_);
  not _31975_ (_00513_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _31976_ (_00514_, _25694_, _00513_);
  and _31977_ (_00516_, _25694_, _00513_);
  nor _31978_ (_00517_, _00516_, _00514_);
  or _31979_ (_00518_, _00517_, _00339_);
  and _31980_ (_00519_, _00518_, _22731_);
  and _31981_ (_26870_[2], _00519_, _00512_);
  and _31982_ (_00520_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _31983_ (_00521_, _00520_, _00439_);
  not _31984_ (_00522_, _00521_);
  nor _31985_ (_00523_, _00522_, _00444_);
  nor _31986_ (_00524_, _00522_, _00441_);
  and _31987_ (_00525_, _00524_, _26541_);
  nor _31988_ (_00526_, _00525_, _00523_);
  not _31989_ (_00528_, _00520_);
  nand _31990_ (_00529_, _00528_, _00447_);
  and _31991_ (_00530_, _00529_, _00526_);
  nand _31992_ (_00531_, _00530_, _23531_);
  not _31993_ (_00532_, _26338_);
  or _31994_ (_00533_, _26377_, _00532_);
  or _31995_ (_00534_, _26364_, _26339_);
  and _31996_ (_00535_, _26363_, _26359_);
  nand _31997_ (_00536_, _00535_, _00534_);
  or _31998_ (_00537_, _00535_, _00534_);
  and _31999_ (_00538_, _00537_, _00536_);
  nand _32000_ (_00539_, _00538_, _26377_);
  nand _32001_ (_00540_, _00539_, _00533_);
  nand _32002_ (_00542_, _00540_, _23528_);
  nor _32003_ (_00543_, _00249_, _22996_);
  not _32004_ (_00544_, _00543_);
  not _32005_ (_00545_, _23463_);
  not _32006_ (_00546_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _32007_ (_00547_, _23462_, _00546_);
  nor _32008_ (_00548_, _00547_, _23563_);
  nor _32009_ (_00549_, _00548_, _23470_);
  and _32010_ (_00550_, _00549_, _00545_);
  not _32011_ (_00551_, _00550_);
  and _32012_ (_00552_, _23409_, _23402_);
  or _32013_ (_00553_, _00552_, _23391_);
  nor _32014_ (_00554_, _00553_, _23410_);
  not _32015_ (_00555_, _00554_);
  or _32016_ (_00556_, _00455_, _23150_);
  and _32017_ (_00557_, _23484_, _23563_);
  nand _32018_ (_00558_, _23535_, _23232_);
  not _32019_ (_00559_, _00558_);
  nor _32020_ (_00560_, _00559_, _00557_);
  and _32021_ (_00561_, _00560_, _00556_);
  and _32022_ (_00562_, _00561_, _23561_);
  not _32023_ (_00563_, _00562_);
  nor _32024_ (_00564_, _00563_, _23575_);
  and _32025_ (_00565_, _00564_, _00555_);
  and _32026_ (_00566_, _00565_, _00551_);
  and _32027_ (_00567_, _00566_, _00544_);
  and _32028_ (_00568_, _00567_, _00542_);
  nand _32029_ (_00569_, _00568_, _00531_);
  and _32030_ (_00570_, _00569_, _26614_);
  and _32031_ (_00571_, _26665_, _26810_);
  and _32032_ (_00572_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _32033_ (_00573_, _00572_, _00571_);
  nand _32034_ (_00574_, _00505_, _00500_);
  and _32035_ (_00575_, _26637_, _24473_);
  nor _32036_ (_00576_, _22737_, _23181_);
  and _32037_ (_00577_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _32038_ (_00578_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _32039_ (_00579_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _32040_ (_00580_, _00579_, _00578_);
  and _32041_ (_00581_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _32042_ (_00582_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or _32043_ (_00583_, _00582_, _00581_);
  or _32044_ (_00584_, _00583_, _00580_);
  and _32045_ (_00585_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _32046_ (_00586_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _32047_ (_00587_, _00586_, _00585_);
  or _32048_ (_00588_, _00587_, _00584_);
  and _32049_ (_00589_, _00588_, _23623_);
  or _32050_ (_00590_, _00589_, _00577_);
  and _32051_ (_00591_, _00590_, _22737_);
  nor _32052_ (_00592_, _00591_, _00576_);
  and _32053_ (_00593_, _00592_, _26635_);
  nor _32054_ (_00594_, _00593_, _00575_);
  and _32055_ (_00595_, _00594_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _32056_ (_00597_, _00594_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _32057_ (_00598_, _00597_, _00595_);
  nand _32058_ (_00599_, _00598_, _00574_);
  or _32059_ (_00600_, _00598_, _00574_);
  and _32060_ (_00601_, _00600_, _26662_);
  and _32061_ (_00602_, _00601_, _00599_);
  or _32062_ (_00603_, _00602_, _00573_);
  or _32063_ (_00604_, _00603_, _00570_);
  not _32064_ (_00605_, _00592_);
  nand _32065_ (_00606_, _00605_, _26606_);
  nand _32066_ (_00607_, _00606_, _00339_);
  or _32067_ (_00608_, _00607_, _00604_);
  and _32068_ (_00609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not _32069_ (_00610_, _00609_);
  nor _32070_ (_00611_, _00610_, _25694_);
  nor _32071_ (_00612_, _00514_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _32072_ (_00613_, _00612_, _00611_);
  or _32073_ (_00614_, _00613_, _00339_);
  and _32074_ (_00615_, _00614_, _22731_);
  and _32075_ (_26870_[3], _00615_, _00608_);
  nand _32076_ (_00616_, _26370_, _26368_);
  or _32077_ (_00617_, _26370_, _26368_);
  nand _32078_ (_00618_, _00617_, _00616_);
  nand _32079_ (_00619_, _00618_, _26377_);
  or _32080_ (_00620_, _26377_, _26326_);
  and _32081_ (_00621_, _00620_, _00619_);
  nand _32082_ (_00622_, _00621_, _23528_);
  or _32083_ (_00623_, _00525_, _00523_);
  and _32084_ (_00624_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  nand _32085_ (_00625_, _00624_, _00623_);
  or _32086_ (_00626_, _00624_, _00623_);
  and _32087_ (_00627_, _00626_, _00625_);
  nand _32088_ (_00628_, _00627_, _23531_);
  and _32089_ (_00629_, _00247_, _22995_);
  not _32090_ (_00630_, _00629_);
  nor _32091_ (_00631_, _23413_, _23173_);
  not _32092_ (_00632_, _00631_);
  nor _32093_ (_00633_, _23414_, _23391_);
  and _32094_ (_00634_, _00633_, _00632_);
  not _32095_ (_00635_, _00634_);
  and _32096_ (_00636_, _23484_, _23460_);
  not _32097_ (_00637_, _00636_);
  or _32098_ (_00638_, _00374_, _23199_);
  nand _32099_ (_00639_, _23534_, _23115_);
  and _32100_ (_00640_, _00639_, _00638_);
  and _32101_ (_00641_, _00640_, _00637_);
  nand _32102_ (_00642_, _00641_, _24075_);
  nor _32103_ (_00643_, _23464_, _23460_);
  not _32104_ (_00644_, _00643_);
  nor _32105_ (_00645_, _23465_, _23470_);
  and _32106_ (_00646_, _00645_, _00644_);
  not _32107_ (_00647_, _00646_);
  nand _32108_ (_00648_, _00647_, _24072_);
  or _32109_ (_00649_, _00648_, _00642_);
  nor _32110_ (_00650_, _00649_, _24079_);
  and _32111_ (_00651_, _00650_, _00635_);
  and _32112_ (_00652_, _00651_, _00630_);
  and _32113_ (_00653_, _00652_, _00628_);
  nand _32114_ (_00654_, _00653_, _00622_);
  and _32115_ (_00655_, _00654_, _26614_);
  not _32116_ (_00656_, _25577_);
  and _32117_ (_00658_, _26665_, _00656_);
  nor _32118_ (_00659_, _22737_, _23131_);
  and _32119_ (_00660_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _32120_ (_00661_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _32121_ (_00662_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _32122_ (_00663_, _00662_, _00661_);
  and _32123_ (_00664_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _32124_ (_00665_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _32125_ (_00666_, _00665_, _00664_);
  or _32126_ (_00667_, _00666_, _00663_);
  and _32127_ (_00668_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _32128_ (_00669_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _32129_ (_00670_, _00669_, _00668_);
  or _32130_ (_00671_, _00670_, _00667_);
  and _32131_ (_00672_, _00671_, _23623_);
  or _32132_ (_00673_, _00672_, _00660_);
  and _32133_ (_00675_, _00673_, _22737_);
  nor _32134_ (_00676_, _00675_, _00659_);
  not _32135_ (_00677_, _00676_);
  and _32136_ (_00678_, _00677_, _26606_);
  and _32137_ (_00679_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _32138_ (_00680_, _00679_, _00678_);
  or _32139_ (_00681_, _00680_, _00658_);
  and _32140_ (_00682_, _26637_, _25577_);
  and _32141_ (_00683_, _00676_, _26635_);
  nor _32142_ (_00684_, _00683_, _00682_);
  nand _32143_ (_00685_, _00684_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _32144_ (_00686_, _00684_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _32145_ (_00687_, _00686_, _00685_);
  nor _32146_ (_00688_, _00595_, _00574_);
  nor _32147_ (_00689_, _00688_, _00597_);
  or _32148_ (_00690_, _00689_, _00687_);
  nand _32149_ (_00691_, _00689_, _00687_);
  and _32150_ (_00692_, _00691_, _26662_);
  and _32151_ (_00693_, _00692_, _00690_);
  nor _32152_ (_00694_, _00693_, _00681_);
  nand _32153_ (_00695_, _00694_, _00339_);
  or _32154_ (_00696_, _00695_, _00655_);
  and _32155_ (_00697_, _00611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _32156_ (_00698_, _00611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _32157_ (_00699_, _00698_, _00697_);
  or _32158_ (_00700_, _00699_, _00339_);
  and _32159_ (_00701_, _00700_, _22731_);
  and _32160_ (_26870_[4], _00701_, _00696_);
  nand _32161_ (_00702_, _00347_, _26320_);
  and _32162_ (_00703_, _00616_, _26328_);
  nand _32163_ (_00704_, _00703_, _26371_);
  or _32164_ (_00705_, _00703_, _26371_);
  nand _32165_ (_00706_, _00705_, _00704_);
  nand _32166_ (_00707_, _00706_, _26377_);
  nand _32167_ (_00708_, _00707_, _00702_);
  nand _32168_ (_00709_, _00708_, _23528_);
  and _32169_ (_00710_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _32170_ (_00711_, _00710_, _00624_);
  nand _32171_ (_00712_, _00711_, _00623_);
  not _32172_ (_00713_, _00710_);
  nand _32173_ (_00714_, _00713_, _00625_);
  and _32174_ (_00715_, _00714_, _00712_);
  nand _32175_ (_00716_, _00715_, _23531_);
  nor _32176_ (_00717_, _23417_, _23414_);
  nor _32177_ (_00718_, _00717_, _23418_);
  and _32178_ (_00719_, _00718_, _23390_);
  not _32179_ (_00720_, _00719_);
  nor _32180_ (_00721_, _00258_, _22996_);
  nor _32181_ (_00722_, _23458_, _23039_);
  nor _32182_ (_00723_, _00722_, _23464_);
  and _32183_ (_00724_, _00723_, _23364_);
  and _32184_ (_00725_, _00724_, _23457_);
  not _32185_ (_00726_, _00724_);
  nor _32186_ (_00727_, _23465_, _23115_);
  and _32187_ (_00728_, _23465_, _23115_);
  nor _32188_ (_00729_, _00728_, _00727_);
  and _32189_ (_00730_, _00729_, _00726_);
  or _32190_ (_00731_, _00730_, _23470_);
  nor _32191_ (_00732_, _00731_, _00725_);
  and _32192_ (_00733_, _23484_, _23115_);
  not _32193_ (_00734_, _00733_);
  or _32194_ (_00735_, _00374_, _23150_);
  or _32195_ (_00736_, _00455_, _23079_);
  and _32196_ (_00737_, _00736_, _00735_);
  and _32197_ (_00738_, _00737_, _00734_);
  and _32198_ (_00739_, _00738_, _24039_);
  not _32199_ (_00740_, _00739_);
  nor _32200_ (_00741_, _00740_, _00732_);
  and _32201_ (_00742_, _00741_, _24032_);
  not _32202_ (_00743_, _00742_);
  nor _32203_ (_00744_, _00743_, _00721_);
  and _32204_ (_00745_, _00744_, _00720_);
  and _32205_ (_00746_, _00745_, _00716_);
  nand _32206_ (_00747_, _00746_, _00709_);
  and _32207_ (_00748_, _00747_, _26614_);
  and _32208_ (_00749_, _26665_, _00033_);
  not _32209_ (_00750_, _26089_);
  and _32210_ (_00751_, _26606_, _00750_);
  and _32211_ (_00752_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _32212_ (_00753_, _00752_, _00751_);
  or _32213_ (_00754_, _00753_, _00749_);
  nand _32214_ (_00755_, _00691_, _00685_);
  and _32215_ (_00756_, _26637_, _26050_);
  and _32216_ (_00757_, _26635_, _26089_);
  nor _32217_ (_00758_, _00757_, _00756_);
  and _32218_ (_00759_, _00758_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _32219_ (_00760_, _00758_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _32220_ (_00761_, _00760_, _00759_);
  or _32221_ (_00762_, _00761_, _00755_);
  and _32222_ (_00763_, _00761_, _00755_);
  not _32223_ (_00764_, _00763_);
  and _32224_ (_00765_, _00764_, _26662_);
  and _32225_ (_00766_, _00765_, _00762_);
  nor _32226_ (_00767_, _00766_, _00754_);
  nand _32227_ (_00768_, _00767_, _00339_);
  or _32228_ (_00769_, _00768_, _00748_);
  and _32229_ (_00770_, _00697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _32230_ (_00771_, _00697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _32231_ (_00772_, _00771_, _00770_);
  or _32232_ (_00773_, _00772_, _00339_);
  and _32233_ (_00774_, _00773_, _22731_);
  and _32234_ (_26870_[5], _00774_, _00769_);
  and _32235_ (_00775_, _26374_, _26313_);
  nor _32236_ (_00776_, _26374_, _26313_);
  or _32237_ (_00777_, _00776_, _00775_);
  and _32238_ (_00778_, _00777_, _26377_);
  nor _32239_ (_00779_, _26377_, _26306_);
  or _32240_ (_00780_, _00779_, _00778_);
  or _32241_ (_00781_, _00780_, _23529_);
  not _32242_ (_00782_, _23531_);
  and _32243_ (_00783_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not _32244_ (_00784_, _00783_);
  nor _32245_ (_00785_, _00784_, _00712_);
  and _32246_ (_00786_, _00784_, _00712_);
  or _32247_ (_00787_, _00786_, _00785_);
  or _32248_ (_00788_, _00787_, _00782_);
  nor _32249_ (_00789_, _00263_, _22996_);
  not _32250_ (_00790_, _00789_);
  nor _32251_ (_00791_, _23423_, _23418_);
  nor _32252_ (_00792_, _00791_, _23391_);
  and _32253_ (_00793_, _00792_, _23425_);
  and _32254_ (_00794_, _00726_, _23466_);
  and _32255_ (_00795_, _00726_, _00727_);
  nor _32256_ (_00796_, _00795_, _23079_);
  nor _32257_ (_00797_, _00796_, _00794_);
  nor _32258_ (_00798_, _00797_, _23470_);
  and _32259_ (_00799_, _23484_, _23959_);
  not _32260_ (_00800_, _00799_);
  or _32261_ (_00801_, _00455_, _23039_);
  nand _32262_ (_00802_, _23535_, _23115_);
  and _32263_ (_00803_, _00802_, _00801_);
  and _32264_ (_00804_, _00803_, _00800_);
  and _32265_ (_00805_, _00804_, _24122_);
  not _32266_ (_00806_, _00805_);
  nor _32267_ (_00807_, _00806_, _00798_);
  and _32268_ (_00808_, _00807_, _24115_);
  not _32269_ (_00809_, _00808_);
  nor _32270_ (_00810_, _00809_, _00793_);
  and _32271_ (_00811_, _00810_, _00790_);
  and _32272_ (_00812_, _00811_, _00788_);
  and _32273_ (_00813_, _00812_, _00781_);
  not _32274_ (_00814_, _00813_);
  and _32275_ (_00815_, _00814_, _26614_);
  not _32276_ (_00816_, _26108_);
  and _32277_ (_00817_, _26606_, _00816_);
  and _32278_ (_00818_, _26665_, _00070_);
  and _32279_ (_00819_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _32280_ (_00820_, _00819_, _00818_);
  or _32281_ (_00821_, _00820_, _00817_);
  or _32282_ (_00822_, _00763_, _00759_);
  and _32283_ (_00823_, _26637_, _00069_);
  and _32284_ (_00824_, _26635_, _26108_);
  nor _32285_ (_00825_, _00824_, _00823_);
  nand _32286_ (_00826_, _00825_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _32287_ (_00827_, _00825_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _32288_ (_00828_, _00827_, _00826_);
  or _32289_ (_00829_, _00828_, _00822_);
  nand _32290_ (_00830_, _00828_, _00822_);
  and _32291_ (_00831_, _00830_, _26662_);
  and _32292_ (_00832_, _00831_, _00829_);
  or _32293_ (_00833_, _00832_, _00821_);
  or _32294_ (_00834_, _00833_, _00815_);
  and _32295_ (_00835_, _00834_, _00339_);
  and _32296_ (_00836_, _00770_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _32297_ (_00837_, _00770_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _32298_ (_00838_, _00837_, _00836_);
  nor _32299_ (_00839_, _00838_, _00339_);
  or _32300_ (_00840_, _00839_, _00835_);
  and _32301_ (_26870_[6], _00840_, _22731_);
  nor _32302_ (_00841_, _00836_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _32303_ (_00842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _32304_ (_00843_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _32305_ (_00844_, _00843_, _00842_);
  and _32306_ (_00845_, _00844_, _00609_);
  not _32307_ (_00846_, _00845_);
  nor _32308_ (_00847_, _00846_, _25694_);
  nor _32309_ (_00848_, _00847_, _00841_);
  or _32310_ (_00849_, _00848_, _00339_);
  and _32311_ (_00850_, _00849_, _22731_);
  or _32312_ (_00851_, _26377_, _26298_);
  nor _32313_ (_00852_, _00775_, _26307_);
  nor _32314_ (_00853_, _00852_, _26311_);
  or _32315_ (_00854_, _00853_, _00347_);
  and _32316_ (_00855_, _00854_, _00851_);
  and _32317_ (_00856_, _00855_, _23528_);
  not _32318_ (_00857_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and _32319_ (_00858_, _00785_, _00857_);
  or _32320_ (_00859_, _26393_, _00857_);
  nor _32321_ (_00860_, _00859_, _00785_);
  or _32322_ (_00861_, _00860_, _00858_);
  and _32323_ (_00862_, _00861_, _23531_);
  and _32324_ (_00863_, _00243_, _22995_);
  nand _32325_ (_00864_, _23427_, _23393_);
  and _32326_ (_00865_, _00864_, _23429_);
  and _32327_ (_00866_, _00865_, _23390_);
  nor _32328_ (_00867_, _00724_, _23466_);
  nor _32329_ (_00868_, _00867_, _23487_);
  or _32330_ (_00869_, _23467_, _23470_);
  or _32331_ (_00870_, _00869_, _00868_);
  and _32332_ (_00871_, _23492_, _23456_);
  nor _32333_ (_00872_, _00374_, _23079_);
  and _32334_ (_00873_, _23484_, _23487_);
  and _32335_ (_00874_, _23441_, _23491_);
  or _32336_ (_00875_, _00874_, _00873_);
  or _32337_ (_00876_, _00875_, _00872_);
  nor _32338_ (_00877_, _00876_, _00871_);
  and _32339_ (_00878_, _00877_, _00870_);
  nand _32340_ (_00879_, _00878_, _23988_);
  or _32341_ (_00880_, _00879_, _00866_);
  or _32342_ (_00881_, _00880_, _00863_);
  or _32343_ (_00882_, _00881_, _00862_);
  or _32344_ (_00883_, _00882_, _00856_);
  and _32345_ (_00884_, _00883_, _26614_);
  not _32346_ (_00885_, _00139_);
  and _32347_ (_00886_, _26665_, _00885_);
  and _32348_ (_00887_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _32349_ (_00888_, _00887_, _00886_);
  nand _32350_ (_00889_, _00830_, _00826_);
  and _32351_ (_00890_, _26637_, _00139_);
  and _32352_ (_00891_, _26635_, _25475_);
  nor _32353_ (_00892_, _00891_, _00890_);
  and _32354_ (_00893_, _00892_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _32355_ (_00894_, _00892_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _32356_ (_00895_, _00894_, _00893_);
  nand _32357_ (_00896_, _00895_, _00889_);
  or _32358_ (_00897_, _00895_, _00889_);
  and _32359_ (_00898_, _00897_, _26662_);
  and _32360_ (_00899_, _00898_, _00896_);
  or _32361_ (_00900_, _00899_, _00888_);
  or _32362_ (_00901_, _00900_, _00884_);
  not _32363_ (_00902_, _25475_);
  nand _32364_ (_00903_, _26606_, _00902_);
  nand _32365_ (_00904_, _00903_, _00339_);
  or _32366_ (_00905_, _00904_, _00901_);
  and _32367_ (_26870_[7], _00905_, _00850_);
  and _32368_ (_00906_, _00847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _32369_ (_00907_, _00847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _32370_ (_00908_, _00907_, _00906_);
  or _32371_ (_00909_, _00908_, _00339_);
  and _32372_ (_00910_, _00909_, _22731_);
  and _32373_ (_00911_, _26570_, _26605_);
  and _32374_ (_00912_, _26606_, _26631_);
  nor _32375_ (_00913_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32376_ (_00914_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23275_);
  nor _32377_ (_00915_, _00914_, _00913_);
  not _32378_ (_00916_, _00915_);
  or _32379_ (_00917_, _00916_, _23430_);
  and _32380_ (_00918_, _00916_, _23430_);
  nor _32381_ (_00919_, _00918_, _23391_);
  and _32382_ (_00920_, _00919_, _00917_);
  nand _32383_ (_00921_, _26377_, _23528_);
  nor _32384_ (_00922_, _23975_, _23472_);
  not _32385_ (_00923_, _00922_);
  nor _32386_ (_00924_, _00923_, _23966_);
  nor _32387_ (_00925_, _00924_, _23301_);
  and _32388_ (_00926_, _00924_, _23301_);
  or _32389_ (_00927_, _00926_, _23953_);
  nor _32390_ (_00928_, _00927_, _00925_);
  and _32391_ (_00929_, _23484_, _23301_);
  and _32392_ (_00930_, _26457_, _23531_);
  and _32393_ (_00931_, _23488_, _23460_);
  nor _32394_ (_00932_, _23974_, _23296_);
  or _32395_ (_00933_, _00932_, _00931_);
  or _32396_ (_00934_, _00933_, _00930_);
  nor _32397_ (_00935_, _00934_, _00929_);
  not _32398_ (_00936_, _00935_);
  nor _32399_ (_00937_, _00936_, _00928_);
  nand _32400_ (_00938_, _00937_, _00921_);
  or _32401_ (_00939_, _00938_, _00920_);
  and _32402_ (_00940_, _00939_, _26574_);
  and _32403_ (_00941_, _26665_, _23765_);
  and _32404_ (_00942_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _32405_ (_00943_, _00942_, _00941_);
  or _32406_ (_00944_, _00943_, _00940_);
  or _32407_ (_00945_, _00944_, _00912_);
  or _32408_ (_00946_, _00945_, _00911_);
  not _32409_ (_00947_, _00339_);
  not _32410_ (_00948_, _00894_);
  and _32411_ (_00949_, _00948_, _00889_);
  or _32412_ (_00950_, _00949_, _00893_);
  and _32413_ (_00951_, _00950_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not _32414_ (_00952_, _00951_);
  or _32415_ (_00953_, _00950_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _32416_ (_00954_, _00953_, _00952_);
  or _32417_ (_00955_, _00954_, _00892_);
  nand _32418_ (_00956_, _00954_, _00892_);
  and _32419_ (_00957_, _00956_, _00955_);
  and _32420_ (_00958_, _00957_, _26662_);
  or _32421_ (_00959_, _00958_, _00947_);
  or _32422_ (_00960_, _00959_, _00946_);
  and _32423_ (_26870_[8], _00960_, _00910_);
  not _32424_ (_00961_, _00892_);
  nor _32425_ (_00962_, _00953_, _00961_);
  and _32426_ (_00963_, _00951_, _00961_);
  nor _32427_ (_00964_, _00963_, _00962_);
  nand _32428_ (_00965_, _00964_, _23243_);
  or _32429_ (_00966_, _00964_, _23243_);
  and _32430_ (_00967_, _00966_, _00965_);
  and _32431_ (_00968_, _00967_, _26662_);
  and _32432_ (_00969_, _00393_, _26605_);
  not _32433_ (_00970_, _26574_);
  nor _32434_ (_00971_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32435_ (_00973_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23243_);
  nor _32436_ (_00974_, _00973_, _00971_);
  not _32437_ (_00975_, _00974_);
  or _32438_ (_00976_, _00975_, _00917_);
  and _32439_ (_00977_, _00975_, _00917_);
  nor _32440_ (_00978_, _00977_, _23391_);
  and _32441_ (_00979_, _00978_, _00976_);
  not _32442_ (_00980_, _00979_);
  and _32443_ (_00981_, _26285_, _23528_);
  not _32444_ (_00982_, _00981_);
  and _32445_ (_00983_, _23484_, _23269_);
  nor _32446_ (_00984_, _23323_, _23039_);
  and _32447_ (_00986_, _00984_, _23964_);
  and _32448_ (_00987_, _00986_, _23364_);
  and _32449_ (_00988_, _23323_, _23039_);
  and _32450_ (_00989_, _00988_, _23957_);
  and _32451_ (_00990_, _00989_, _23456_);
  nor _32452_ (_00991_, _00990_, _00987_);
  nor _32453_ (_00992_, _00991_, _23305_);
  and _32454_ (_00993_, _00991_, _23305_);
  or _32455_ (_00995_, _00993_, _23953_);
  nor _32456_ (_00996_, _00995_, _00992_);
  and _32457_ (_00997_, _26410_, _23491_);
  not _32458_ (_00998_, _00997_);
  and _32459_ (_00999_, _00998_, _26424_);
  nor _32460_ (_01000_, _00999_, _26458_);
  and _32461_ (_01001_, _01000_, _23531_);
  and _32462_ (_01002_, _23488_, _23115_);
  and _32463_ (_01003_, _23506_, _23264_);
  or _32464_ (_01004_, _01003_, _01002_);
  or _32465_ (_01005_, _01004_, _01001_);
  or _32466_ (_01006_, _01005_, _00996_);
  nor _32467_ (_01007_, _01006_, _00983_);
  and _32468_ (_01008_, _01007_, _00982_);
  and _32469_ (_01009_, _01008_, _00980_);
  nor _32470_ (_01010_, _01009_, _00970_);
  and _32471_ (_01011_, _26665_, _23745_);
  and _32472_ (_01012_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _32473_ (_01013_, _26606_, _00157_);
  or _32474_ (_01014_, _01013_, _01012_);
  or _32475_ (_01015_, _01014_, _01011_);
  or _32476_ (_01016_, _01015_, _01010_);
  or _32477_ (_01017_, _01016_, _00969_);
  or _32478_ (_01018_, _01017_, _00968_);
  and _32479_ (_01019_, _01018_, _00339_);
  nor _32480_ (_01020_, _00906_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _32481_ (_01021_, _00906_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _32482_ (_01022_, _01021_, _01020_);
  nor _32483_ (_01023_, _01022_, _00339_);
  or _32484_ (_01024_, _01023_, _01019_);
  and _32485_ (_26870_[9], _01024_, _22731_);
  nor _32486_ (_01025_, _01021_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _32487_ (_01026_, _01021_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _32488_ (_01027_, _01026_, _01025_);
  or _32489_ (_01028_, _01027_, _00339_);
  and _32490_ (_01029_, _01028_, _22731_);
  and _32491_ (_01030_, _00473_, _26605_);
  nor _32492_ (_01031_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32493_ (_01032_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23215_);
  nor _32494_ (_01033_, _01032_, _01031_);
  not _32495_ (_01034_, _01033_);
  and _32496_ (_01035_, _01034_, _00976_);
  not _32497_ (_01036_, _01035_);
  or _32498_ (_01037_, _01034_, _00976_);
  and _32499_ (_01038_, _01037_, _23390_);
  and _32500_ (_01039_, _01038_, _01036_);
  not _32501_ (_01040_, _01039_);
  nor _32502_ (_01041_, _26525_, _26522_);
  nor _32503_ (_01042_, _01041_, _26526_);
  and _32504_ (_01043_, _01042_, _23531_);
  and _32505_ (_01044_, _23488_, _23959_);
  and _32506_ (_01045_, _23484_, _23237_);
  or _32507_ (_01046_, _01045_, _01044_);
  nor _32508_ (_01047_, _01046_, _01043_);
  and _32509_ (_01048_, _00990_, _23305_);
  and _32510_ (_01049_, _00986_, _23269_);
  and _32511_ (_01050_, _01049_, _23364_);
  nor _32512_ (_01051_, _01050_, _01048_);
  nor _32513_ (_01052_, _01051_, _23310_);
  and _32514_ (_01053_, _01051_, _23310_);
  or _32515_ (_01054_, _01053_, _23953_);
  nor _32516_ (_01055_, _01054_, _01052_);
  and _32517_ (_01056_, _23506_, _23232_);
  and _32518_ (_01057_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or _32519_ (_01058_, _01057_, _01056_);
  nor _32520_ (_01059_, _01058_, _01055_);
  and _32521_ (_01060_, _01059_, _01047_);
  and _32522_ (_01061_, _01060_, _01040_);
  nor _32523_ (_01062_, _01061_, _00970_);
  and _32524_ (_01063_, _26665_, _23724_);
  and _32525_ (_01064_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _32526_ (_01065_, _01064_, _01063_);
  or _32527_ (_01066_, _01065_, _01062_);
  or _32528_ (_01067_, _01066_, _01030_);
  and _32529_ (_01068_, _00962_, _23243_);
  and _32530_ (_01069_, _00963_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _32531_ (_01071_, _01069_, _01068_);
  nand _32532_ (_01072_, _01071_, _23215_);
  or _32533_ (_01073_, _01071_, _23215_);
  and _32534_ (_01074_, _01073_, _01072_);
  and _32535_ (_01075_, _01074_, _26662_);
  or _32536_ (_01076_, _01075_, _01067_);
  nand _32537_ (_01077_, _26606_, _00224_);
  nand _32538_ (_01078_, _01077_, _00339_);
  or _32539_ (_01079_, _01078_, _01076_);
  and _32540_ (_26870_[10], _01079_, _01029_);
  nor _32541_ (_01080_, _01026_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _32542_ (_01081_, _01026_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _32543_ (_01082_, _01081_, _01080_);
  or _32544_ (_01083_, _01082_, _00339_);
  and _32545_ (_01084_, _01083_, _22731_);
  and _32546_ (_01085_, _00569_, _26605_);
  nor _32547_ (_01086_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32548_ (_01087_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23177_);
  nor _32549_ (_01088_, _01087_, _01086_);
  not _32550_ (_01089_, _01088_);
  and _32551_ (_01090_, _01089_, _01037_);
  not _32552_ (_01091_, _01090_);
  or _32553_ (_01092_, _01089_, _01037_);
  and _32554_ (_01094_, _01092_, _23390_);
  and _32555_ (_01095_, _01094_, _01091_);
  not _32556_ (_01096_, _01095_);
  and _32557_ (_01097_, _26529_, _26527_);
  not _32558_ (_01098_, _01097_);
  and _32559_ (_01099_, _01098_, _26530_);
  and _32560_ (_01100_, _01099_, _23531_);
  not _32561_ (_01101_, _01100_);
  and _32562_ (_01102_, _01049_, _23237_);
  nor _32563_ (_01103_, _01102_, _23456_);
  nor _32564_ (_01104_, _23269_, _23237_);
  and _32565_ (_01105_, _01104_, _00989_);
  nor _32566_ (_01106_, _01105_, _23364_);
  or _32567_ (_01107_, _01106_, _01103_);
  and _32568_ (_01108_, _01107_, _23205_);
  nor _32569_ (_01109_, _01107_, _23205_);
  nor _32570_ (_01110_, _01109_, _01108_);
  and _32571_ (_01111_, _01110_, _23514_);
  and _32572_ (_01112_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _32573_ (_01113_, _23974_, _23199_);
  and _32574_ (_01114_, _23484_, _23371_);
  or _32575_ (_01115_, _01114_, _01113_);
  or _32576_ (_01116_, _01115_, _23489_);
  nor _32577_ (_01117_, _01116_, _01112_);
  not _32578_ (_01118_, _01117_);
  nor _32579_ (_01119_, _01118_, _01111_);
  and _32580_ (_01120_, _01119_, _01101_);
  and _32581_ (_01121_, _01120_, _01096_);
  nor _32582_ (_01122_, _01121_, _00970_);
  and _32583_ (_01123_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _32584_ (_01124_, _26606_, _26810_);
  or _32585_ (_01125_, _01124_, _01123_);
  or _32586_ (_01126_, _01125_, _01122_);
  or _32587_ (_01127_, _01126_, _01085_);
  and _32588_ (_01128_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _32589_ (_01129_, _01128_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _32590_ (_01130_, _01129_, _00949_);
  nor _32591_ (_01131_, _01130_, _00892_);
  or _32592_ (_01132_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _32593_ (_01133_, _01132_, _00953_);
  and _32594_ (_01134_, _01133_, _00892_);
  nor _32595_ (_01135_, _01134_, _01131_);
  or _32596_ (_01136_, _01135_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _32597_ (_01137_, _01135_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _32598_ (_01138_, _01137_, _01136_);
  and _32599_ (_01139_, _01138_, _26662_);
  or _32600_ (_01140_, _01139_, _01127_);
  and _32601_ (_01141_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _32602_ (_01142_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _32603_ (_01143_, _01142_, _01141_);
  and _32604_ (_01144_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _32605_ (_01145_, _01144_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _32606_ (_01146_, _01145_, _01143_);
  and _32607_ (_01147_, _01146_, _01129_);
  and _32608_ (_01148_, _01147_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _32609_ (_01149_, _01147_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _32610_ (_01150_, _01149_, _01148_);
  nand _32611_ (_01151_, _01150_, _26665_);
  nand _32612_ (_01152_, _01151_, _00339_);
  or _32613_ (_01153_, _01152_, _01140_);
  and _32614_ (_26870_[11], _01153_, _01084_);
  and _32615_ (_01154_, _00654_, _26605_);
  nor _32616_ (_01155_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32617_ (_01156_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23128_);
  nor _32618_ (_01157_, _01156_, _01155_);
  not _32619_ (_01158_, _01157_);
  and _32620_ (_01159_, _01158_, _01092_);
  not _32621_ (_01160_, _01159_);
  or _32622_ (_01161_, _01158_, _01092_);
  and _32623_ (_01162_, _01161_, _23390_);
  and _32624_ (_01163_, _01162_, _01160_);
  not _32625_ (_01164_, _01163_);
  and _32626_ (_01165_, _26533_, _26531_);
  not _32627_ (_01166_, _01165_);
  and _32628_ (_01167_, _01166_, _26534_);
  and _32629_ (_01168_, _01167_, _23531_);
  not _32630_ (_01169_, _01168_);
  and _32631_ (_01170_, _01105_, _23205_);
  and _32632_ (_01171_, _01170_, _23456_);
  and _32633_ (_01172_, _01102_, _23371_);
  and _32634_ (_01173_, _01172_, _23364_);
  nor _32635_ (_01174_, _01173_, _01171_);
  and _32636_ (_01175_, _01174_, _23169_);
  nor _32637_ (_01176_, _01174_, _23169_);
  nor _32638_ (_01177_, _01176_, _01175_);
  and _32639_ (_01178_, _01177_, _23514_);
  and _32640_ (_01179_, _23506_, _23364_);
  nor _32641_ (_01180_, _01179_, _23484_);
  or _32642_ (_01181_, _01180_, _23169_);
  or _32643_ (_01182_, _23974_, _23150_);
  or _32644_ (_01183_, _01182_, _23364_);
  and _32645_ (_01184_, _23488_, _23491_);
  and _32646_ (_01185_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _32647_ (_01186_, _01185_, _01184_);
  and _32648_ (_01187_, _01186_, _01183_);
  and _32649_ (_01188_, _01187_, _01181_);
  not _32650_ (_01189_, _01188_);
  nor _32651_ (_01190_, _01189_, _01178_);
  and _32652_ (_01191_, _01190_, _01169_);
  and _32653_ (_01192_, _01191_, _01164_);
  nor _32654_ (_01193_, _01192_, _00970_);
  and _32655_ (_01194_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _32656_ (_01195_, _26606_, _00656_);
  or _32657_ (_01197_, _01195_, _01194_);
  or _32658_ (_01198_, _01197_, _01193_);
  or _32659_ (_01199_, _01198_, _01154_);
  and _32660_ (_01200_, _01129_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _32661_ (_01201_, _01200_, _00950_);
  nor _32662_ (_01202_, _01201_, _00892_);
  nor _32663_ (_01203_, _01133_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _32664_ (_01204_, _01203_, _00892_);
  nor _32665_ (_01205_, _01204_, _01202_);
  nand _32666_ (_01206_, _01205_, _23128_);
  or _32667_ (_01207_, _01205_, _23128_);
  and _32668_ (_01208_, _01207_, _01206_);
  and _32669_ (_01209_, _01208_, _26662_);
  or _32670_ (_01210_, _01209_, _01199_);
  or _32671_ (_01211_, _01148_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _32672_ (_01212_, _01148_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not _32673_ (_01213_, _01212_);
  and _32674_ (_01214_, _01213_, _26665_);
  nand _32675_ (_01215_, _01214_, _01211_);
  nand _32676_ (_01216_, _01215_, _00339_);
  or _32677_ (_01217_, _01216_, _01210_);
  not _32678_ (_01218_, _25694_);
  and _32679_ (_01219_, _00845_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _32680_ (_01220_, _01219_, _01218_);
  not _32681_ (_01221_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand _32682_ (_01222_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _32683_ (_01223_, _01222_, _01221_);
  nand _32684_ (_01225_, _01223_, _01220_);
  nor _32685_ (_01226_, _01225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _32686_ (_01227_, _01225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _32687_ (_01228_, _01227_, _01226_);
  or _32688_ (_01229_, _01228_, _00339_);
  and _32689_ (_01230_, _01229_, _22731_);
  and _32690_ (_26870_[12], _01230_, _01217_);
  not _32691_ (_01231_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _32692_ (_01232_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _32693_ (_01233_, _01225_, _01232_);
  nand _32694_ (_01234_, _01233_, _01231_);
  or _32695_ (_01236_, _01233_, _01231_);
  and _32696_ (_01237_, _01236_, _01234_);
  or _32697_ (_01238_, _01237_, _00339_);
  and _32698_ (_01239_, _01238_, _22731_);
  and _32699_ (_01240_, _00747_, _26605_);
  nor _32700_ (_01241_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _32701_ (_01242_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23092_);
  nor _32702_ (_01243_, _01242_, _01241_);
  not _32703_ (_01244_, _01243_);
  and _32704_ (_01245_, _01244_, _01161_);
  not _32705_ (_01246_, _01245_);
  or _32706_ (_01247_, _01244_, _01161_);
  and _32707_ (_01248_, _01247_, _23390_);
  and _32708_ (_01249_, _01248_, _01246_);
  not _32709_ (_01250_, _01249_);
  and _32710_ (_01251_, _26535_, _26513_);
  not _32711_ (_01252_, _01251_);
  and _32712_ (_01253_, _01252_, _26536_);
  and _32713_ (_01255_, _01253_, _23531_);
  and _32714_ (_01256_, _01172_, _23156_);
  nor _32715_ (_01257_, _01256_, _23456_);
  and _32716_ (_01258_, _23205_, _23169_);
  and _32717_ (_01259_, _01258_, _01105_);
  nor _32718_ (_01260_, _01259_, _23364_);
  or _32719_ (_01261_, _01260_, _01257_);
  nor _32720_ (_01262_, _01261_, _23122_);
  and _32721_ (_01263_, _01261_, _23122_);
  nor _32722_ (_01264_, _01263_, _01262_);
  nor _32723_ (_01265_, _01264_, _23953_);
  and _32724_ (_01266_, _23364_, _23122_);
  nor _32725_ (_01267_, _23364_, _23457_);
  nor _32726_ (_01268_, _01267_, _01266_);
  nor _32727_ (_01269_, _01268_, _23974_);
  and _32728_ (_01270_, _23484_, _23122_);
  and _32729_ (_01271_, _23488_, _23264_);
  and _32730_ (_01272_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or _32731_ (_01273_, _01272_, _01271_);
  nor _32732_ (_01274_, _01273_, _01270_);
  not _32733_ (_01275_, _01274_);
  nor _32734_ (_01276_, _01275_, _01269_);
  not _32735_ (_01277_, _01276_);
  nor _32736_ (_01278_, _01277_, _01265_);
  not _32737_ (_01279_, _01278_);
  nor _32738_ (_01280_, _01279_, _01255_);
  and _32739_ (_01281_, _01280_, _01250_);
  nor _32740_ (_01282_, _01281_, _00970_);
  and _32741_ (_01283_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _32742_ (_01284_, _26606_, _00033_);
  or _32743_ (_01285_, _01284_, _01283_);
  or _32744_ (_01286_, _01285_, _01282_);
  or _32745_ (_01287_, _01286_, _01240_);
  nor _32746_ (_01288_, _00892_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not _32747_ (_01289_, _01202_);
  nand _32748_ (_01290_, _01203_, _23128_);
  and _32749_ (_01291_, _01290_, _01289_);
  or _32750_ (_01292_, _01291_, _01288_);
  nand _32751_ (_01293_, _01292_, _23092_);
  or _32752_ (_01294_, _01292_, _23092_);
  and _32753_ (_01295_, _01294_, _01293_);
  and _32754_ (_01296_, _01295_, _26662_);
  or _32755_ (_01297_, _01296_, _01287_);
  and _32756_ (_01298_, _01212_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _32757_ (_01299_, _01212_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _32758_ (_01300_, _01299_, _26665_);
  nor _32759_ (_01302_, _01300_, _01298_);
  or _32760_ (_01303_, _01302_, _00947_);
  or _32761_ (_01304_, _01303_, _01297_);
  and _32762_ (_26870_[13], _01304_, _01239_);
  or _32763_ (_01305_, _01298_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _32764_ (_01306_, _01298_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not _32765_ (_01308_, _01306_);
  and _32766_ (_01309_, _01308_, _26665_);
  and _32767_ (_01310_, _01309_, _01305_);
  not _32768_ (_01311_, _26605_);
  nor _32769_ (_01312_, _00813_, _01311_);
  nor _32770_ (_01313_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32771_ (_01314_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23057_);
  nor _32772_ (_01315_, _01314_, _01313_);
  not _32773_ (_01316_, _01315_);
  and _32774_ (_01317_, _01316_, _01247_);
  not _32775_ (_01318_, _01317_);
  or _32776_ (_01319_, _01316_, _01247_);
  and _32777_ (_01320_, _01319_, _23390_);
  and _32778_ (_01321_, _01320_, _01318_);
  not _32779_ (_01322_, _01321_);
  and _32780_ (_01323_, _26537_, _26507_);
  not _32781_ (_01324_, _01323_);
  and _32782_ (_01325_, _01324_, _26538_);
  and _32783_ (_01326_, _01325_, _23531_);
  and _32784_ (_01327_, _01259_, _24022_);
  and _32785_ (_01328_, _01256_, _23122_);
  and _32786_ (_01329_, _01328_, _23364_);
  nor _32787_ (_01330_, _01329_, _01327_);
  nor _32788_ (_01331_, _01330_, _23086_);
  and _32789_ (_01333_, _01330_, _23086_);
  nor _32790_ (_01335_, _01333_, _01331_);
  and _32791_ (_01337_, _01335_, _23514_);
  and _32792_ (_01338_, _23484_, _23084_);
  nor _32793_ (_01339_, _23364_, _23959_);
  not _32794_ (_01340_, _01339_);
  and _32795_ (_01341_, _23364_, _23086_);
  nor _32796_ (_01342_, _01341_, _23974_);
  and _32797_ (_01343_, _01342_, _01340_);
  and _32798_ (_01344_, _23488_, _23232_);
  and _32799_ (_01345_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or _32800_ (_01346_, _01345_, _01344_);
  or _32801_ (_01347_, _01346_, _01343_);
  nor _32802_ (_01348_, _01347_, _01338_);
  not _32803_ (_01349_, _01348_);
  nor _32804_ (_01350_, _01349_, _01337_);
  not _32805_ (_01351_, _01350_);
  nor _32806_ (_01352_, _01351_, _01326_);
  and _32807_ (_01353_, _01352_, _01322_);
  nor _32808_ (_01354_, _01353_, _00970_);
  and _32809_ (_01356_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _32810_ (_01357_, _26606_, _00070_);
  or _32811_ (_01358_, _01357_, _01356_);
  or _32812_ (_01359_, _01358_, _01354_);
  or _32813_ (_01360_, _01359_, _01312_);
  or _32814_ (_01361_, _01290_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _32815_ (_01362_, _01361_, _00961_);
  nand _32816_ (_01363_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _32817_ (_01364_, _01363_, _01201_);
  or _32818_ (_01365_, _01364_, _00892_);
  and _32819_ (_01366_, _01365_, _01362_);
  nand _32820_ (_01367_, _01366_, _23057_);
  or _32821_ (_01369_, _01366_, _23057_);
  and _32822_ (_01370_, _01369_, _01367_);
  and _32823_ (_01371_, _01370_, _26662_);
  or _32824_ (_01372_, _01371_, _01360_);
  or _32825_ (_01373_, _01372_, _01310_);
  or _32826_ (_01374_, _01373_, _00947_);
  not _32827_ (_01375_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _32828_ (_01376_, _01236_, _01375_);
  or _32829_ (_01377_, _01236_, _01375_);
  and _32830_ (_01378_, _01377_, _01376_);
  or _32831_ (_01380_, _01378_, _00339_);
  and _32832_ (_01381_, _01380_, _22731_);
  and _32833_ (_26870_[14], _01381_, _01374_);
  and _32834_ (_01382_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _22731_);
  and _32835_ (_01383_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not _32836_ (_01384_, _23615_);
  nor _32837_ (_01385_, _23639_, _01384_);
  nor _32838_ (_01386_, _23681_, _23660_);
  and _32839_ (_01387_, _01386_, _01385_);
  nor _32840_ (_01389_, _23765_, _23703_);
  not _32841_ (_01390_, _23724_);
  nor _32842_ (_01391_, _23745_, _01390_);
  and _32843_ (_01393_, _01391_, _01389_);
  and _32844_ (_01394_, _01393_, _01387_);
  not _32845_ (_01395_, _23660_);
  and _32846_ (_01396_, _01395_, _23615_);
  not _32847_ (_01397_, _23681_);
  nor _32848_ (_01398_, _01397_, _23639_);
  and _32849_ (_01399_, _01398_, _01396_);
  nor _32850_ (_01400_, _01399_, _01394_);
  and _32851_ (_01401_, _23745_, _01390_);
  not _32852_ (_01402_, _23765_);
  and _32853_ (_01403_, _01402_, _23703_);
  and _32854_ (_01405_, _01403_, _01401_);
  and _32855_ (_01406_, _01405_, _01387_);
  and _32856_ (_01408_, _23765_, _23703_);
  nor _32857_ (_01410_, _23745_, _23724_);
  and _32858_ (_01411_, _01410_, _01408_);
  and _32859_ (_01412_, _01411_, _01387_);
  nor _32860_ (_01413_, _01412_, _01406_);
  and _32861_ (_01414_, _01413_, _01400_);
  and _32862_ (_01415_, _01396_, _23639_);
  and _32863_ (_01416_, _01415_, _23681_);
  and _32864_ (_01417_, _23745_, _23724_);
  and _32865_ (_01418_, _01417_, _01389_);
  and _32866_ (_01419_, _01418_, _01416_);
  and _32867_ (_01420_, _01415_, _01397_);
  not _32868_ (_01422_, _01420_);
  and _32869_ (_01424_, _01408_, _01401_);
  and _32870_ (_01425_, _01410_, _23765_);
  nor _32871_ (_01427_, _01425_, _01424_);
  nor _32872_ (_01428_, _01427_, _01422_);
  nor _32873_ (_01429_, _01428_, _01419_);
  and _32874_ (_01430_, _01429_, _01414_);
  and _32875_ (_01431_, _01385_, _23660_);
  and _32876_ (_01432_, _01431_, _01397_);
  not _32877_ (_01433_, _01432_);
  and _32878_ (_01434_, _01417_, _01403_);
  nor _32879_ (_01435_, _01434_, _01424_);
  nor _32880_ (_01436_, _01435_, _01433_);
  not _32881_ (_01437_, _01436_);
  and _32882_ (_01438_, _01408_, _01391_);
  and _32883_ (_01439_, _01438_, _01387_);
  nor _32884_ (_01440_, _01402_, _23703_);
  and _32885_ (_01441_, _01440_, _01401_);
  and _32886_ (_01442_, _01441_, _01431_);
  nor _32887_ (_01443_, _01442_, _01439_);
  and _32888_ (_01444_, _01401_, _01389_);
  and _32889_ (_01445_, _01444_, _01387_);
  and _32890_ (_01446_, _01401_, _23765_);
  and _32891_ (_01447_, _01446_, _01387_);
  nor _32892_ (_01448_, _01447_, _01445_);
  and _32893_ (_01449_, _01448_, _01443_);
  and _32894_ (_01450_, _01449_, _01437_);
  and _32895_ (_01451_, _01450_, _01430_);
  and _32896_ (_01452_, _01391_, _23765_);
  not _32897_ (_01453_, _01452_);
  and _32898_ (_01454_, _01453_, _01435_);
  nor _32899_ (_01455_, _01454_, _23615_);
  not _32900_ (_01456_, _01455_);
  not _32901_ (_01457_, _01415_);
  and _32902_ (_01458_, _01403_, _01391_);
  nor _32903_ (_01459_, _01458_, _01441_);
  nor _32904_ (_01460_, _01459_, _01457_);
  and _32905_ (_01461_, _01416_, _01410_);
  nor _32906_ (_01462_, _01461_, _01460_);
  and _32907_ (_01463_, _01440_, _01391_);
  nor _32908_ (_01464_, _01458_, _01463_);
  nor _32909_ (_01465_, _01464_, _01433_);
  not _32910_ (_01466_, _01387_);
  and _32911_ (_01467_, _01402_, _23745_);
  and _32912_ (_01468_, _01467_, _23724_);
  nor _32913_ (_01469_, _01463_, _01468_);
  nor _32914_ (_01470_, _01469_, _01466_);
  nor _32915_ (_01471_, _01470_, _01465_);
  and _32916_ (_01472_, _01471_, _01462_);
  and _32917_ (_01473_, _01472_, _01456_);
  and _32918_ (_01474_, _01473_, _01451_);
  and _32919_ (_01475_, _01431_, _23681_);
  and _32920_ (_01476_, _01475_, _01444_);
  and _32921_ (_01477_, _01458_, _01387_);
  nor _32922_ (_01478_, _01477_, _01476_);
  nor _32923_ (_01479_, _01438_, _01418_);
  nor _32924_ (_01480_, _01479_, _01433_);
  not _32925_ (_01481_, _01405_);
  nor _32926_ (_01482_, _01432_, _01415_);
  nor _32927_ (_01483_, _01482_, _01481_);
  nor _32928_ (_01484_, _01483_, _01480_);
  and _32929_ (_01485_, _01484_, _01478_);
  not _32930_ (_01486_, _23703_);
  and _32931_ (_01487_, _23765_, _23724_);
  and _32932_ (_01488_, _01487_, _23745_);
  and _32933_ (_01489_, _01488_, _01486_);
  and _32934_ (_01490_, _01489_, _01416_);
  not _32935_ (_01491_, _01490_);
  and _32936_ (_01492_, _01438_, _01416_);
  and _32937_ (_01493_, _01475_, _01405_);
  nor _32938_ (_01494_, _01493_, _01492_);
  and _32939_ (_01496_, _01494_, _01491_);
  not _32940_ (_01497_, _01393_);
  nor _32941_ (_01498_, _01432_, _01384_);
  nor _32942_ (_01499_, _01498_, _01497_);
  not _32943_ (_01501_, _01424_);
  and _32944_ (_01502_, _01391_, _01486_);
  nor _32945_ (_01503_, _01502_, _01438_);
  and _32946_ (_01505_, _01503_, _01501_);
  and _32947_ (_01506_, _23660_, _23639_);
  and _32948_ (_01507_, _01506_, _23615_);
  not _32949_ (_01508_, _01507_);
  nor _32950_ (_01509_, _01508_, _01505_);
  nor _32951_ (_01510_, _01509_, _01499_);
  and _32952_ (_01511_, _01510_, _01496_);
  and _32953_ (_01512_, _01511_, _01485_);
  and _32954_ (_01513_, _01488_, _23703_);
  and _32955_ (_01514_, _01513_, _01416_);
  nor _32956_ (_01515_, _01514_, _01444_);
  nor _32957_ (_01516_, _01515_, _01482_);
  not _32958_ (_01517_, _01516_);
  and _32959_ (_01518_, _01434_, _01416_);
  and _32960_ (_01519_, _01438_, _01420_);
  nor _32961_ (_01520_, _01519_, _01518_);
  and _32962_ (_01521_, _01410_, _01402_);
  and _32963_ (_01522_, _01521_, _01432_);
  not _32964_ (_01523_, _01522_);
  and _32965_ (_01524_, _01410_, _01403_);
  and _32966_ (_01525_, _01524_, _01387_);
  and _32967_ (_01526_, _01440_, _01410_);
  and _32968_ (_01527_, _01526_, _01387_);
  or _32969_ (_01528_, _01527_, _01525_);
  or _32970_ (_01529_, _01424_, _01393_);
  and _32971_ (_01530_, _01529_, _01416_);
  nor _32972_ (_01531_, _01530_, _01528_);
  and _32973_ (_01532_, _01531_, _01523_);
  and _32974_ (_01533_, _01532_, _01520_);
  and _32975_ (_01534_, _01533_, _01517_);
  and _32976_ (_01535_, _01534_, _01512_);
  and _32977_ (_01536_, _01535_, _01474_);
  and _32978_ (_01537_, _01475_, _01441_);
  or _32979_ (_01538_, _01506_, _01384_);
  and _32980_ (_01539_, _01538_, _01438_);
  or _32981_ (_01540_, _01539_, _01412_);
  nor _32982_ (_01541_, _01540_, _01537_);
  and _32983_ (_01542_, _01541_, _01494_);
  and _32984_ (_01543_, _01542_, _01478_);
  nand _32985_ (_01544_, _01543_, _01533_);
  or _32986_ (_01545_, _01544_, _01536_);
  and _32987_ (_01546_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _32988_ (_01547_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _32989_ (_01548_, _01547_, _01546_);
  and _32990_ (_01549_, _01548_, _01545_);
  nor _32991_ (_01550_, _01548_, _01545_);
  nor _32992_ (_01551_, _01550_, _01549_);
  or _32993_ (_01552_, _01551_, _24471_);
  or _32994_ (_01553_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _32995_ (_01554_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _32996_ (_01555_, _01554_, _01553_);
  and _32997_ (_01556_, _01555_, _01552_);
  or _32998_ (_26871_[0], _01556_, _01383_);
  not _32999_ (_01557_, _01536_);
  and _33000_ (_01558_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _33001_ (_01559_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _33002_ (_01560_, _01559_, _01558_);
  and _33003_ (_01561_, _01560_, _01546_);
  nor _33004_ (_01562_, _01560_, _01546_);
  nor _33005_ (_01563_, _01562_, _01561_);
  nand _33006_ (_01564_, _01563_, _01557_);
  or _33007_ (_01565_, _01563_, _01557_);
  and _33008_ (_01566_, _01565_, _01564_);
  nand _33009_ (_01567_, _01566_, _01549_);
  or _33010_ (_01568_, _01566_, _01549_);
  and _33011_ (_01569_, _01568_, _01567_);
  or _33012_ (_01570_, _01569_, _24471_);
  or _33013_ (_01571_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _33014_ (_01572_, _01571_, _01554_);
  and _33015_ (_01573_, _01572_, _01570_);
  and _33016_ (_01574_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _33017_ (_26871_[1], _01574_, _01573_);
  and _33018_ (_01575_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nand _33019_ (_01576_, _01567_, _01564_);
  nor _33020_ (_01577_, _01561_, _01558_);
  not _33021_ (_01578_, _01577_);
  and _33022_ (_01579_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _33023_ (_01580_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _33024_ (_01581_, _01580_, _01579_);
  and _33025_ (_01582_, _01581_, _01578_);
  nor _33026_ (_01583_, _01581_, _01578_);
  nor _33027_ (_01584_, _01583_, _01582_);
  and _33028_ (_01585_, _01584_, _01576_);
  nor _33029_ (_01586_, _01584_, _01576_);
  nor _33030_ (_01587_, _01586_, _01585_);
  or _33031_ (_01588_, _01587_, _24471_);
  or _33032_ (_01589_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _33033_ (_01590_, _01589_, _01554_);
  and _33034_ (_01591_, _01590_, _01588_);
  or _33035_ (_26871_[2], _01591_, _01575_);
  nor _33036_ (_01592_, _01582_, _01579_);
  nor _33037_ (_01593_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _33038_ (_01594_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _33039_ (_01595_, _01594_, _01593_);
  and _33040_ (_01596_, _01595_, _01585_);
  nor _33041_ (_01597_, _01595_, _01585_);
  nor _33042_ (_01598_, _01597_, _01596_);
  or _33043_ (_01599_, _01598_, _24471_);
  or _33044_ (_01601_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _33045_ (_01602_, _01601_, _01554_);
  and _33046_ (_01603_, _01602_, _01599_);
  and _33047_ (_01605_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _33048_ (_26871_[3], _01605_, _01603_);
  and _33049_ (_01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _33050_ (_01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _33051_ (_01609_, _01608_, _01607_);
  nand _33052_ (_01610_, _01609_, _01593_);
  or _33053_ (_01611_, _01609_, _01593_);
  and _33054_ (_01612_, _01611_, _01610_);
  and _33055_ (_01613_, _01612_, _01596_);
  nor _33056_ (_01614_, _01612_, _01596_);
  nor _33057_ (_01615_, _01614_, _01613_);
  or _33058_ (_01616_, _01615_, _24471_);
  or _33059_ (_01617_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _33060_ (_01618_, _01617_, _01554_);
  and _33061_ (_01619_, _01618_, _01616_);
  and _33062_ (_01620_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _33063_ (_26871_[4], _01620_, _01619_);
  not _33064_ (_01621_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33065_ (_01622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _01621_);
  and _33066_ (_01623_, _01622_, _22731_);
  nand _33067_ (_01624_, _01608_, _01592_);
  and _33068_ (_01625_, _01624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not _33069_ (_01626_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _33070_ (_01627_, _01608_, _01626_);
  and _33071_ (_01628_, _01627_, _01592_);
  or _33072_ (_01629_, _01628_, _01625_);
  or _33073_ (_01630_, _01629_, _01613_);
  and _33074_ (_01631_, _01629_, _01612_);
  and _33075_ (_01632_, _01631_, _01596_);
  nor _33076_ (_01633_, _01632_, _24471_);
  and _33077_ (_01634_, _01633_, _01630_);
  nor _33078_ (_01635_, _24470_, _23090_);
  or _33079_ (_01636_, _01635_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33080_ (_01637_, _01636_, _01634_);
  and _33081_ (_26871_[5], _01637_, _01623_);
  not _33082_ (_01638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _33083_ (_01639_, _01628_, _01638_);
  and _33084_ (_01640_, _01627_, _01638_);
  and _33085_ (_01641_, _01640_, _01592_);
  nor _33086_ (_01642_, _01641_, _01639_);
  not _33087_ (_01643_, _01642_);
  and _33088_ (_01644_, _01643_, _01632_);
  nor _33089_ (_01645_, _01643_, _01632_);
  nor _33090_ (_01646_, _01645_, _01644_);
  or _33091_ (_01647_, _01646_, _24471_);
  or _33092_ (_01648_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _33093_ (_01649_, _01648_, _01554_);
  and _33094_ (_01650_, _01649_, _01647_);
  and _33095_ (_01651_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _33096_ (_26871_[6], _01651_, _01650_);
  and _33097_ (_01652_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _33098_ (_01653_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _33099_ (_01654_, _01640_, _01653_);
  and _33100_ (_01655_, _01654_, _01592_);
  nor _33101_ (_01656_, _01641_, _01653_);
  nor _33102_ (_01657_, _01656_, _01655_);
  not _33103_ (_01658_, _01657_);
  and _33104_ (_01659_, _01658_, _01644_);
  nor _33105_ (_01660_, _01658_, _01644_);
  nor _33106_ (_01661_, _01660_, _01659_);
  or _33107_ (_01663_, _01661_, _24471_);
  or _33108_ (_01664_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _33109_ (_01665_, _01664_, _01554_);
  and _33110_ (_01666_, _01665_, _01663_);
  or _33111_ (_26871_[7], _01666_, _01652_);
  not _33112_ (_01667_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _33113_ (_01668_, _01655_, _01667_);
  and _33114_ (_01669_, _01654_, _01667_);
  and _33115_ (_01670_, _01669_, _01592_);
  or _33116_ (_01671_, _01670_, _01668_);
  and _33117_ (_01672_, _01671_, _01659_);
  nor _33118_ (_01673_, _01671_, _01659_);
  nor _33119_ (_01674_, _01673_, _01672_);
  or _33120_ (_01675_, _01674_, _24471_);
  or _33121_ (_01676_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _33122_ (_01677_, _01676_, _01554_);
  and _33123_ (_01678_, _01677_, _01675_);
  and _33124_ (_01679_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _33125_ (_26871_[8], _01679_, _01678_);
  not _33126_ (_01680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _33127_ (_01681_, _01669_, _01680_);
  and _33128_ (_01682_, _01681_, _01592_);
  nor _33129_ (_01683_, _01670_, _01680_);
  nor _33130_ (_01684_, _01683_, _01682_);
  not _33131_ (_01685_, _01684_);
  and _33132_ (_01686_, _01685_, _01672_);
  or _33133_ (_01687_, _01685_, _01672_);
  nand _33134_ (_01689_, _01687_, _24470_);
  nor _33135_ (_01690_, _01689_, _01686_);
  nor _33136_ (_01691_, _24470_, _23243_);
  or _33137_ (_01692_, _01691_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33138_ (_01693_, _01692_, _01690_);
  or _33139_ (_01694_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _01621_);
  and _33140_ (_01695_, _01694_, _22731_);
  and _33141_ (_26871_[9], _01695_, _01693_);
  not _33142_ (_01696_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _33143_ (_01697_, _01682_, _01696_);
  and _33144_ (_01699_, _01681_, _01696_);
  and _33145_ (_01700_, _01699_, _01592_);
  nor _33146_ (_01701_, _01700_, _01697_);
  not _33147_ (_01702_, _01701_);
  and _33148_ (_01703_, _01702_, _01686_);
  nor _33149_ (_01704_, _01702_, _01686_);
  nor _33150_ (_01705_, _01704_, _01703_);
  or _33151_ (_01706_, _01705_, _24471_);
  or _33152_ (_01707_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _33153_ (_01708_, _01707_, _01554_);
  and _33154_ (_01709_, _01708_, _01706_);
  and _33155_ (_01710_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _33156_ (_26871_[10], _01710_, _01709_);
  and _33157_ (_01711_, _01699_, _01221_);
  and _33158_ (_01712_, _01711_, _01592_);
  nor _33159_ (_01713_, _01700_, _01221_);
  nor _33160_ (_01714_, _01713_, _01712_);
  not _33161_ (_01715_, _01714_);
  and _33162_ (_01716_, _01715_, _01703_);
  or _33163_ (_01717_, _01715_, _01703_);
  nand _33164_ (_01718_, _01717_, _24470_);
  nor _33165_ (_01719_, _01718_, _01716_);
  nor _33166_ (_01720_, _24470_, _23177_);
  or _33167_ (_01721_, _01720_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33168_ (_01722_, _01721_, _01719_);
  or _33169_ (_01723_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _01621_);
  and _33170_ (_01724_, _01723_, _22731_);
  and _33171_ (_26871_[11], _01724_, _01722_);
  nor _33172_ (_01725_, _01712_, _01232_);
  and _33173_ (_01726_, _01711_, _01232_);
  and _33174_ (_01727_, _01726_, _01592_);
  or _33175_ (_01728_, _01727_, _01725_);
  and _33176_ (_01730_, _01728_, _01716_);
  nor _33177_ (_01731_, _01728_, _01716_);
  nor _33178_ (_01732_, _01731_, _01730_);
  or _33179_ (_01733_, _01732_, _24471_);
  or _33180_ (_01734_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _33181_ (_01735_, _01734_, _01554_);
  and _33182_ (_01736_, _01735_, _01733_);
  and _33183_ (_01737_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _33184_ (_26871_[12], _01737_, _01736_);
  and _33185_ (_01738_, _01727_, _01231_);
  nor _33186_ (_01739_, _01727_, _01231_);
  nor _33187_ (_01740_, _01739_, _01738_);
  not _33188_ (_01741_, _01740_);
  and _33189_ (_01742_, _01741_, _01730_);
  nor _33190_ (_01743_, _01741_, _01730_);
  nor _33191_ (_01744_, _01743_, _01742_);
  or _33192_ (_01745_, _01744_, _24471_);
  or _33193_ (_01746_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _33194_ (_01747_, _01746_, _01554_);
  and _33195_ (_01748_, _01747_, _01745_);
  and _33196_ (_01749_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _33197_ (_26871_[13], _01749_, _01748_);
  nor _33198_ (_01750_, _01738_, _01375_);
  and _33199_ (_01751_, _01738_, _01375_);
  nor _33200_ (_01752_, _01751_, _01750_);
  not _33201_ (_01753_, _01752_);
  and _33202_ (_01754_, _01753_, _01742_);
  nor _33203_ (_01755_, _01753_, _01742_);
  nor _33204_ (_01756_, _01755_, _01754_);
  or _33205_ (_01757_, _01756_, _24471_);
  or _33206_ (_01758_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _33207_ (_01759_, _01758_, _01554_);
  and _33208_ (_01760_, _01759_, _01757_);
  and _33209_ (_01761_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _33210_ (_26871_[14], _01761_, _01760_);
  and _33211_ (_01762_, _25648_, _24051_);
  and _33212_ (_01763_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or _33213_ (_22617_, _01763_, _01762_);
  and _33214_ (_01764_, _26020_, _24134_);
  and _33215_ (_01765_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or _33216_ (_22618_, _01765_, _01764_);
  nor _33217_ (_01766_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor _33218_ (_01767_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _33219_ (_01768_, _01767_, _01766_);
  not _33220_ (_01769_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor _33221_ (_01770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _33222_ (_01771_, _01770_, _01769_);
  and _33223_ (_01772_, _01771_, _01768_);
  and _33224_ (_01773_, _01772_, _25010_);
  and _33225_ (_01774_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _33226_ (_01775_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _33227_ (_26875_[0], _01775_, _22731_);
  and _33228_ (_01776_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _33229_ (_01777_, _01776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _33230_ (_26875_[1], _01777_, _22731_);
  and _33231_ (_01778_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _33232_ (_01779_, _01778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _33233_ (_26875_[2], _01779_, _22731_);
  and _33234_ (_01780_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _33235_ (_01781_, _01780_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _33236_ (_26875_[3], _01781_, _22731_);
  and _33237_ (_01782_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _33238_ (_01783_, _01782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _33239_ (_26875_[4], _01783_, _22731_);
  and _33240_ (_01784_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _33241_ (_01785_, _01784_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _33242_ (_26875_[5], _01785_, _22731_);
  and _33243_ (_01786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22731_);
  and _33244_ (_01787_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _22731_);
  and _33245_ (_01788_, _01787_, _01773_);
  or _33246_ (_26875_[6], _01788_, _01786_);
  and _33247_ (_01789_, _01545_, _22737_);
  nand _33248_ (_01790_, _01789_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _33249_ (_01791_, _01789_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _33250_ (_01792_, _01791_, _01554_);
  and _33251_ (_26876_[0], _01792_, _01790_);
  and _33252_ (_01793_, _01545_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _33253_ (_01794_, _01536_, _23599_);
  nand _33254_ (_01795_, _01536_, _23599_);
  and _33255_ (_01796_, _01795_, _01794_);
  nand _33256_ (_01797_, _01796_, _01793_);
  or _33257_ (_01798_, _01796_, _01793_);
  and _33258_ (_01800_, _01798_, _01797_);
  or _33259_ (_01801_, _01800_, _25454_);
  or _33260_ (_01802_, _22737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _33261_ (_01803_, _01802_, _01554_);
  and _33262_ (_26876_[1], _01803_, _01801_);
  and _33263_ (_01804_, _26020_, _24051_);
  and _33264_ (_01805_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or _33265_ (_22619_, _01805_, _01804_);
  and _33266_ (_01806_, _26020_, _24089_);
  and _33267_ (_01807_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or _33268_ (_22621_, _01807_, _01806_);
  and _33269_ (_01808_, _24320_, _23583_);
  and _33270_ (_01809_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _33271_ (_22622_, _01809_, _01808_);
  and _33272_ (_01810_, _24301_, _24095_);
  and _33273_ (_01811_, _01810_, _24219_);
  not _33274_ (_01812_, _01810_);
  and _33275_ (_01813_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or _33276_ (_22623_, _01813_, _01811_);
  and _33277_ (_01814_, _25497_, _24174_);
  nor _33278_ (_01815_, _01814_, rst);
  and _33279_ (_01816_, _25607_, _24174_);
  not _33280_ (_01817_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _33281_ (_01818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _33282_ (_01819_, _01818_, _01817_);
  and _33283_ (_01820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _33284_ (_01821_, _01820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _33285_ (_01822_, _01821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _33286_ (_01823_, _01822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _33287_ (_01824_, _01823_, _01818_);
  and _33288_ (_01825_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _33289_ (_01826_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _33290_ (_01827_, _01826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _33291_ (_01828_, _01827_, _01819_);
  and _33292_ (_01829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _33293_ (_01830_, _01829_, _01828_);
  nor _33294_ (_01831_, _01830_, _01816_);
  and _33295_ (_22624_, _01831_, _01815_);
  and _33296_ (_01832_, _24476_, _24372_);
  and _33297_ (_01833_, _01832_, _24051_);
  not _33298_ (_01834_, _01832_);
  and _33299_ (_01835_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _33300_ (_22625_, _01835_, _01833_);
  not _33301_ (_01836_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and _33302_ (_01837_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _33303_ (_01838_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _33304_ (_01839_, _01838_, _01837_);
  and _33305_ (_26879_[0], _01839_, _22731_);
  and _33306_ (_01840_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _33307_ (_01841_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33308_ (_01842_, _01841_, _01840_);
  and _33309_ (_26879_[1], _01842_, _22731_);
  and _33310_ (_01843_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _33311_ (_01844_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33312_ (_01845_, _01844_, _01843_);
  and _33313_ (_26879_[2], _01845_, _22731_);
  and _33314_ (_01846_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _33315_ (_01847_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33316_ (_01848_, _01847_, _01846_);
  and _33317_ (_26879_[3], _01848_, _22731_);
  and _33318_ (_01849_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _33319_ (_01850_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33320_ (_01851_, _01850_, _01849_);
  and _33321_ (_26879_[4], _01851_, _22731_);
  and _33322_ (_01852_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _33323_ (_01853_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33324_ (_01854_, _01853_, _01852_);
  and _33325_ (_26879_[5], _01854_, _22731_);
  and _33326_ (_01855_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _33327_ (_01856_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33328_ (_01857_, _01856_, _01855_);
  and _33329_ (_26879_[6], _01857_, _22731_);
  not _33330_ (_01858_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _33331_ (_01859_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor _33332_ (_01860_, _01859_, _01858_);
  and _33333_ (_01861_, _01859_, _01858_);
  nor _33334_ (_01862_, _01861_, _01860_);
  and _33335_ (_26882_[0], _01862_, _22731_);
  nor _33336_ (_01863_, _01860_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _33337_ (_01864_, _01860_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _33338_ (_01865_, _01864_, _01863_);
  nor _33339_ (_26882_[1], _01865_, rst);
  and _33340_ (_01866_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _33341_ (_01867_, _01866_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _33342_ (_01868_, _01866_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _33343_ (_01869_, _01868_, _01867_);
  or _33344_ (_01870_, _01869_, _01859_);
  and _33345_ (_26882_[2], _01870_, _22731_);
  and _33346_ (_01871_, _01832_, _24089_);
  and _33347_ (_01872_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _33348_ (_27066_, _01872_, _01871_);
  and _33349_ (_01873_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _33350_ (_01874_, _25694_, _25696_);
  or _33351_ (_01875_, _01874_, _01873_);
  and _33352_ (_26884_[0], _01875_, _22731_);
  and _33353_ (_01876_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _33354_ (_01877_, _25694_, _25700_);
  or _33355_ (_01878_, _01877_, _01876_);
  and _33356_ (_26884_[1], _01878_, _22731_);
  and _33357_ (_01879_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _33358_ (_01880_, _25694_, _25705_);
  or _33359_ (_01881_, _01880_, _01879_);
  and _33360_ (_26884_[2], _01881_, _22731_);
  and _33361_ (_01882_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _33362_ (_01883_, _25694_, _25711_);
  or _33363_ (_01884_, _01883_, _01882_);
  and _33364_ (_26884_[3], _01884_, _22731_);
  and _33365_ (_01885_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _33366_ (_01886_, _25694_, _25715_);
  or _33367_ (_01887_, _01886_, _01885_);
  and _33368_ (_26884_[4], _01887_, _22731_);
  and _33369_ (_01888_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _33370_ (_01889_, _25694_, _25720_);
  or _33371_ (_01890_, _01889_, _01888_);
  and _33372_ (_26884_[5], _01890_, _22731_);
  and _33373_ (_01891_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _33374_ (_01892_, _25694_, _25724_);
  or _33375_ (_01893_, _01892_, _01891_);
  and _33376_ (_26884_[6], _01893_, _22731_);
  and _33377_ (_01894_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _33378_ (_01895_, _25694_, _25729_);
  or _33379_ (_01896_, _01895_, _01894_);
  and _33380_ (_26884_[7], _01896_, _22731_);
  and _33381_ (_01897_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _33382_ (_01898_, _25694_, _25735_);
  or _33383_ (_01899_, _01898_, _01897_);
  and _33384_ (_26884_[8], _01899_, _22731_);
  and _33385_ (_01900_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _33386_ (_01901_, _25694_, _25739_);
  or _33387_ (_01902_, _01901_, _01900_);
  and _33388_ (_26884_[9], _01902_, _22731_);
  and _33389_ (_01903_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _33390_ (_01904_, _25694_, _25744_);
  or _33391_ (_01905_, _01904_, _01903_);
  and _33392_ (_26884_[10], _01905_, _22731_);
  and _33393_ (_01906_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _33394_ (_01907_, _25694_, _25750_);
  or _33395_ (_01908_, _01907_, _01906_);
  and _33396_ (_26884_[11], _01908_, _22731_);
  and _33397_ (_01909_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _33398_ (_01910_, _25694_, _25754_);
  or _33399_ (_01911_, _01910_, _01909_);
  and _33400_ (_26884_[12], _01911_, _22731_);
  and _33401_ (_01912_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _33402_ (_01913_, _25694_, _25758_);
  or _33403_ (_01914_, _01913_, _01912_);
  and _33404_ (_26884_[13], _01914_, _22731_);
  and _33405_ (_01915_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _33406_ (_01916_, _25694_, _25763_);
  or _33407_ (_01917_, _01916_, _01915_);
  and _33408_ (_26884_[14], _01917_, _22731_);
  and _33409_ (_01918_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _33410_ (_01919_, _25694_, _25767_);
  or _33411_ (_01920_, _01919_, _01918_);
  and _33412_ (_26884_[15], _01920_, _22731_);
  and _33413_ (_01921_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _33414_ (_01922_, _25694_, _25771_);
  or _33415_ (_01923_, _01922_, _01921_);
  and _33416_ (_26884_[16], _01923_, _22731_);
  and _33417_ (_01924_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _33418_ (_01926_, _25694_, _25776_);
  or _33419_ (_01927_, _01926_, _01924_);
  and _33420_ (_26884_[17], _01927_, _22731_);
  and _33421_ (_01928_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _33422_ (_01929_, _25694_, _25780_);
  or _33423_ (_01930_, _01929_, _01928_);
  and _33424_ (_26884_[18], _01930_, _22731_);
  and _33425_ (_01931_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _33426_ (_01932_, _25694_, _25784_);
  or _33427_ (_01933_, _01932_, _01931_);
  and _33428_ (_26884_[19], _01933_, _22731_);
  and _33429_ (_01934_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _33430_ (_01935_, _25694_, _25788_);
  or _33431_ (_01936_, _01935_, _01934_);
  and _33432_ (_26884_[20], _01936_, _22731_);
  and _33433_ (_01937_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _33434_ (_01938_, _25694_, _25792_);
  or _33435_ (_01939_, _01938_, _01937_);
  and _33436_ (_26884_[21], _01939_, _22731_);
  and _33437_ (_01940_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _33438_ (_01941_, _25694_, _25796_);
  or _33439_ (_01942_, _01941_, _01940_);
  and _33440_ (_26884_[22], _01942_, _22731_);
  and _33441_ (_01943_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _33442_ (_01944_, _25694_, _25800_);
  or _33443_ (_01945_, _01944_, _01943_);
  and _33444_ (_26884_[23], _01945_, _22731_);
  and _33445_ (_01946_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _33446_ (_01947_, _25694_, _25804_);
  or _33447_ (_01948_, _01947_, _01946_);
  and _33448_ (_26884_[24], _01948_, _22731_);
  and _33449_ (_01949_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _33450_ (_01950_, _25694_, _25808_);
  or _33451_ (_01951_, _01950_, _01949_);
  and _33452_ (_26884_[25], _01951_, _22731_);
  and _33453_ (_01952_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _33454_ (_01953_, _25694_, _25812_);
  or _33455_ (_01954_, _01953_, _01952_);
  and _33456_ (_26884_[26], _01954_, _22731_);
  and _33457_ (_01955_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _33458_ (_01956_, _25694_, _25816_);
  or _33459_ (_01957_, _01956_, _01955_);
  and _33460_ (_26884_[27], _01957_, _22731_);
  and _33461_ (_01958_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _33462_ (_01959_, _25694_, _25820_);
  or _33463_ (_01960_, _01959_, _01958_);
  and _33464_ (_26884_[28], _01960_, _22731_);
  and _33465_ (_01961_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _33466_ (_01962_, _25694_, _25825_);
  or _33467_ (_01963_, _01962_, _01961_);
  and _33468_ (_26884_[29], _01963_, _22731_);
  and _33469_ (_01964_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _33470_ (_01965_, _25694_, _25829_);
  or _33471_ (_01966_, _01965_, _01964_);
  and _33472_ (_26884_[30], _01966_, _22731_);
  and _33473_ (_01967_, _24257_, _23780_);
  and _33474_ (_01968_, _23926_, _23780_);
  or _33475_ (_01969_, _26673_, _24244_);
  or _33476_ (_01970_, _01969_, _01968_);
  or _33477_ (_01971_, _01970_, _01967_);
  or _33478_ (_01972_, _01971_, _26749_);
  and _33479_ (_01973_, _23844_, _23687_);
  or _33480_ (_01974_, _23912_, _23790_);
  or _33481_ (_01975_, _01974_, _01973_);
  or _33482_ (_01976_, _23836_, _23773_);
  or _33483_ (_01977_, _01976_, _24267_);
  and _33484_ (_01978_, _23827_, _23687_);
  and _33485_ (_01979_, _26693_, _23687_);
  or _33486_ (_01980_, _01979_, _23898_);
  or _33487_ (_01981_, _01980_, _01978_);
  or _33488_ (_01982_, _01981_, _01977_);
  or _33489_ (_01983_, _01982_, _01975_);
  or _33490_ (_01984_, _24269_, _23916_);
  and _33491_ (_01985_, _23911_, _23816_);
  and _33492_ (_01986_, _23814_, _23789_);
  and _33493_ (_01987_, _23825_, _23788_);
  or _33494_ (_01988_, _01987_, _01986_);
  or _33495_ (_01989_, _01988_, _01985_);
  and _33496_ (_01990_, _23781_, _23786_);
  and _33497_ (_01991_, _01990_, _23707_);
  and _33498_ (_01992_, _01991_, _23803_);
  and _33499_ (_01993_, _23911_, _23814_);
  or _33500_ (_01994_, _01993_, _23830_);
  or _33501_ (_01995_, _01994_, _01992_);
  or _33502_ (_01996_, _01995_, _01989_);
  or _33503_ (_01997_, _01996_, _01984_);
  or _33504_ (_01998_, _01997_, _01983_);
  or _33505_ (_01999_, _01998_, _01972_);
  and _33506_ (_02000_, _01999_, _22737_);
  and _33507_ (_02001_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _33508_ (_02002_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _33509_ (_02003_, _26601_, _02002_);
  nor _33510_ (_02004_, _24246_, _23708_);
  and _33511_ (_02005_, _23816_, _23788_);
  nor _33512_ (_02006_, _02005_, _24246_);
  nand _33513_ (_02007_, _23788_, _23779_);
  and _33514_ (_02008_, _02007_, _02006_);
  nor _33515_ (_02009_, _02008_, _02004_);
  and _33516_ (_02010_, _02009_, _02003_);
  or _33517_ (_02011_, _02010_, _26681_);
  or _33518_ (_02012_, _02011_, _02001_);
  or _33519_ (_02013_, _02012_, _02000_);
  and _33520_ (_26849_[1], _02013_, _22731_);
  and _33521_ (_02014_, _23830_, _23791_);
  and _33522_ (_02015_, _26594_, _23707_);
  or _33523_ (_02016_, _02015_, _24251_);
  or _33524_ (_02017_, _02016_, _02014_);
  and _33525_ (_02018_, _23803_, _23789_);
  and _33526_ (_02019_, _01991_, _23814_);
  and _33527_ (_02020_, _01991_, _23824_);
  and _33528_ (_02021_, _26593_, _23707_);
  or _33529_ (_02022_, _02021_, _02020_);
  or _33530_ (_02023_, _02022_, _02019_);
  or _33531_ (_02024_, _02023_, _02018_);
  and _33532_ (_02025_, _23926_, _23687_);
  or _33533_ (_02026_, _02025_, _23910_);
  or _33534_ (_02027_, _24273_, _24258_);
  or _33535_ (_02028_, _02027_, _02026_);
  or _33536_ (_02029_, _02028_, _02024_);
  or _33537_ (_02031_, _01984_, _24250_);
  or _33538_ (_02032_, _02031_, _02029_);
  or _33539_ (_02033_, _02032_, _02017_);
  or _33540_ (_02034_, _02033_, _01983_);
  and _33541_ (_02035_, _02034_, _22737_);
  and _33542_ (_02036_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _33543_ (_02037_, _02036_, _02011_);
  or _33544_ (_02038_, _02037_, _02035_);
  and _33545_ (_26849_[0], _02038_, _22731_);
  and _33546_ (_02039_, _24097_, _23944_);
  and _33547_ (_02040_, _02039_, _24159_);
  not _33548_ (_02041_, _02040_);
  and _33549_ (_02043_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _33550_ (_02044_, _02040_, _23996_);
  or _33551_ (_22626_, _02044_, _02043_);
  nand _33552_ (_26842_[0], _02009_, _23855_);
  and _33553_ (_02045_, _24301_, _24159_);
  and _33554_ (_02046_, _02045_, _23583_);
  not _33555_ (_02047_, _02045_);
  and _33556_ (_02048_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _33557_ (_27232_, _02048_, _02046_);
  nor _33558_ (_02049_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _33559_ (_02050_, _02049_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not _33560_ (_02051_, _02050_);
  or _33561_ (_02053_, _02051_, _26570_);
  or _33562_ (_02054_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _33563_ (_02055_, _02054_, _22731_);
  and _33564_ (_26888_[0], _02055_, _02053_);
  or _33565_ (_02056_, _02051_, _00393_);
  or _33566_ (_02057_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _33567_ (_02058_, _02057_, _22731_);
  and _33568_ (_26888_[1], _02058_, _02056_);
  or _33569_ (_02059_, _02051_, _00473_);
  or _33570_ (_02060_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _33571_ (_02061_, _02060_, _22731_);
  and _33572_ (_26888_[2], _02061_, _02059_);
  or _33573_ (_02062_, _02051_, _00569_);
  or _33574_ (_02063_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _33575_ (_02064_, _02063_, _22731_);
  and _33576_ (_26888_[3], _02064_, _02062_);
  and _33577_ (_02065_, _24236_, _24006_);
  and _33578_ (_02066_, _02065_, _24219_);
  not _33579_ (_02067_, _02065_);
  and _33580_ (_02068_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or _33581_ (_22627_, _02068_, _02066_);
  and _33582_ (_02069_, _02045_, _24089_);
  and _33583_ (_02070_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _33584_ (_22628_, _02070_, _02069_);
  and _33585_ (_02071_, _24553_, _24174_);
  or _33586_ (_02072_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _33587_ (_02073_, _02072_, _22731_);
  not _33588_ (_02074_, _02071_);
  or _33589_ (_02075_, _02074_, _23880_);
  and _33590_ (_22629_, _02075_, _02073_);
  and _33591_ (_02076_, _01832_, _24134_);
  and _33592_ (_02077_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _33593_ (_22630_, _02077_, _02076_);
  nor _33594_ (_02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _33595_ (_02079_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _33596_ (_02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _22731_);
  and _33597_ (_02082_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _33598_ (_22631_, _02082_, _02079_);
  and _33599_ (_02083_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _33600_ (_02084_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _33601_ (_22632_, _02084_, _02083_);
  and _33602_ (_02085_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _33603_ (_02086_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _33604_ (_22633_, _02086_, _02085_);
  and _33605_ (_02087_, _01832_, _23996_);
  and _33606_ (_02088_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _33607_ (_22634_, _02088_, _02087_);
  and _33608_ (_02089_, _02045_, _24051_);
  and _33609_ (_02090_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _33610_ (_22635_, _02090_, _02089_);
  and _33611_ (_02091_, _25648_, _23548_);
  and _33612_ (_02092_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or _33613_ (_22636_, _02092_, _02091_);
  and _33614_ (_02093_, _24476_, _24146_);
  and _33615_ (_02094_, _02093_, _23583_);
  not _33616_ (_02095_, _02093_);
  and _33617_ (_02096_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _33618_ (_27037_, _02096_, _02094_);
  and _33619_ (_02097_, _02093_, _24051_);
  and _33620_ (_02098_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _33621_ (_22637_, _02098_, _02097_);
  and _33622_ (_02100_, _02093_, _24089_);
  and _33623_ (_02101_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _33624_ (_22638_, _02101_, _02100_);
  and _33625_ (_22639_, _01786_, _24747_);
  and _33626_ (_02102_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _33627_ (_02103_, _02102_, _24841_);
  and _33628_ (_22640_, _02103_, _22731_);
  or _33629_ (_02104_, _24844_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _33630_ (_02105_, _02104_, _22731_);
  not _33631_ (_02106_, _24763_);
  or _33632_ (_02107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _33633_ (_02108_, _02107_, _02106_);
  nor _33634_ (_02109_, _24915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _33635_ (_02110_, _02109_, _24919_);
  and _33636_ (_02111_, _02110_, _02108_);
  or _33637_ (_02112_, _02111_, _24757_);
  and _33638_ (_02113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _24750_);
  nand _33639_ (_02114_, _24777_, _24763_);
  nand _33640_ (_02115_, _02114_, _24758_);
  nand _33641_ (_02116_, _02115_, _02113_);
  nand _33642_ (_02117_, _02116_, _02112_);
  and _33643_ (_02118_, _02117_, _24809_);
  and _33644_ (_02119_, _24805_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  not _33645_ (_02120_, _24802_);
  and _33646_ (_02121_, _02107_, _02120_);
  or _33647_ (_02122_, _24931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _33648_ (_02123_, _24930_, _24802_);
  and _33649_ (_02124_, _02123_, _02122_);
  or _33650_ (_02125_, _02124_, _02121_);
  and _33651_ (_02126_, _02125_, _24797_);
  and _33652_ (_02127_, _24802_, _24790_);
  or _33653_ (_02129_, _02127_, _24795_);
  and _33654_ (_02130_, _02129_, _02113_);
  or _33655_ (_02131_, _02130_, _02126_);
  and _33656_ (_02132_, _02131_, _24806_);
  or _33657_ (_02133_, _02132_, _02119_);
  and _33658_ (_02134_, _02133_, _24781_);
  or _33659_ (_02135_, _02134_, _02118_);
  or _33660_ (_02136_, _02135_, _24747_);
  and _33661_ (_22641_, _02136_, _02105_);
  and _33662_ (_02137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _33663_ (_02138_, _02137_, _24777_);
  or _33664_ (_02139_, _24848_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _33665_ (_02140_, _02139_, _24846_);
  or _33666_ (_02141_, _02140_, _02138_);
  and _33667_ (_02142_, _02141_, _24763_);
  or _33668_ (_02143_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _24750_);
  and _33669_ (_02144_, _02143_, _02106_);
  or _33670_ (_02145_, _02144_, _02142_);
  and _33671_ (_02146_, _02145_, _25006_);
  and _33672_ (_02147_, _02143_, _02120_);
  or _33673_ (_02148_, _24870_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _33674_ (_02149_, _24869_, _24802_);
  and _33675_ (_02150_, _02149_, _02148_);
  or _33676_ (_02152_, _02150_, _02147_);
  and _33677_ (_02153_, _02152_, _24943_);
  or _33678_ (_02154_, _02153_, _02146_);
  and _33679_ (_02155_, _02154_, _24844_);
  and _33680_ (_02156_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _33681_ (_02157_, _02156_, _24805_);
  and _33682_ (_02158_, _02157_, _24781_);
  nand _33683_ (_02159_, _24757_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _33684_ (_02160_, _02159_, _24781_);
  or _33685_ (_02161_, _02160_, _24747_);
  or _33686_ (_02162_, _02161_, _02158_);
  and _33687_ (_02163_, _02162_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _33688_ (_02164_, _02163_, _02155_);
  and _33689_ (_22642_, _02164_, _22731_);
  and _33690_ (_02166_, _24621_, _24607_);
  nand _33691_ (_02167_, _02166_, _23504_);
  or _33692_ (_02168_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _33693_ (_02169_, _02168_, _24630_);
  and _33694_ (_02170_, _02169_, _02167_);
  nor _33695_ (_02171_, _24630_, _24043_);
  or _33696_ (_02172_, _02171_, _02170_);
  and _33697_ (_22643_, _02172_, _22731_);
  and _33698_ (_02173_, _24636_, _24544_);
  and _33699_ (_02174_, _02173_, _23504_);
  nor _33700_ (_02175_, _02173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _33701_ (_02176_, _02175_, _02174_);
  nand _33702_ (_02177_, _02176_, _24557_);
  nand _33703_ (_02178_, _24554_, _24082_);
  and _33704_ (_02179_, _02178_, _22731_);
  and _33705_ (_22644_, _02179_, _02177_);
  and _33706_ (_02180_, _24451_, _23996_);
  and _33707_ (_02181_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _33708_ (_22645_, _02181_, _02180_);
  and _33709_ (_02182_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _33710_ (_02183_, _02040_, _23887_);
  or _33711_ (_27028_, _02183_, _02182_);
  and _33712_ (_02184_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and _33713_ (_02185_, _02040_, _23583_);
  or _33714_ (_27029_, _02185_, _02184_);
  and _33715_ (_02186_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and _33716_ (_02187_, _02040_, _23548_);
  or _33717_ (_22646_, _02187_, _02186_);
  and _33718_ (_02188_, _01832_, _24219_);
  and _33719_ (_02189_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _33720_ (_22647_, _02189_, _02188_);
  and _33721_ (_02190_, _02093_, _23996_);
  and _33722_ (_02191_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _33723_ (_22648_, _02191_, _02190_);
  nand _33724_ (_02192_, _01816_, _23989_);
  not _33725_ (_02193_, _01814_);
  or _33726_ (_02194_, _02193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _33727_ (_02195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _33728_ (_02196_, _02195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _33729_ (_02197_, _02195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _33730_ (_02198_, _02197_, _02196_);
  not _33731_ (_02199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _33732_ (_02200_, _02199_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _33733_ (_02201_, t0_i);
  and _33734_ (_02202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _02201_);
  and _33735_ (_02203_, _02202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  or _33736_ (_02204_, _02203_, _02200_);
  and _33737_ (_02205_, _02204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _33738_ (_02206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _33739_ (_02207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _33740_ (_02208_, _02207_, _02206_);
  and _33741_ (_02209_, _02208_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _33742_ (_02210_, _02209_, _02205_);
  and _33743_ (_02211_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _33744_ (_02212_, _02211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _33745_ (_02213_, _02212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _33746_ (_02214_, _02213_, _02198_);
  nand _33747_ (_02215_, _02196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _33748_ (_02216_, _02212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand _33749_ (_02217_, _02216_, _02215_);
  and _33750_ (_02218_, _02217_, _02214_);
  nor _33751_ (_02219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _33752_ (_02220_, _02219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _33753_ (_02221_, _02216_);
  and _33754_ (_02222_, _02221_, _01829_);
  or _33755_ (_02223_, _02222_, _02220_);
  and _33756_ (_02224_, _02223_, _02213_);
  or _33757_ (_02225_, _02224_, _02218_);
  or _33758_ (_02226_, _02225_, _01814_);
  and _33759_ (_02227_, _02226_, _02194_);
  or _33760_ (_02228_, _02227_, _01816_);
  and _33761_ (_02229_, _02228_, _22731_);
  and _33762_ (_22649_, _02229_, _02192_);
  and _33763_ (_02230_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _33764_ (_02231_, _02040_, _24051_);
  or _33765_ (_22650_, _02231_, _02230_);
  and _33766_ (_02232_, _24476_, _24140_);
  and _33767_ (_02233_, _02232_, _24051_);
  not _33768_ (_02234_, _02232_);
  and _33769_ (_02235_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or _33770_ (_22651_, _02235_, _02233_);
  not _33771_ (_02236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _33772_ (_02237_, _02236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not _33773_ (_02238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _33774_ (_02239_, t1_i);
  and _33775_ (_02240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _02239_);
  nor _33776_ (_02241_, _02240_, _02238_);
  not _33777_ (_02242_, _02241_);
  not _33778_ (_02243_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _33779_ (_02244_, _02243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nor _33780_ (_02245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _33781_ (_02246_, _02245_);
  and _33782_ (_02247_, _02246_, _02244_);
  and _33783_ (_02248_, _02247_, _02242_);
  not _33784_ (_02249_, _02248_);
  and _33785_ (_02250_, _02249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _33786_ (_02251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _33787_ (_02252_, _02251_, _02248_);
  and _33788_ (_02253_, _02252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _33789_ (_02254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not _33790_ (_02255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _33791_ (_02256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _33792_ (_02257_, _02256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand _33793_ (_02258_, _02257_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _33794_ (_02259_, _02258_, _02255_);
  and _33795_ (_02260_, _02259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _33796_ (_02262_, _02260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _33797_ (_02263_, _02262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _33798_ (_02264_, _02263_, _02254_);
  and _33799_ (_02265_, _02264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _33800_ (_02266_, _02265_, _02253_);
  and _33801_ (_02267_, _02266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _33802_ (_02268_, _02267_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _33803_ (_02269_, _02268_, _02250_);
  and _33804_ (_02270_, _02269_, _02237_);
  nor _33805_ (_02271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _33806_ (_02272_, _02259_, _02254_);
  and _33807_ (_02273_, _02272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _33808_ (_02274_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _33809_ (_02275_, _02274_, _02251_);
  and _33810_ (_02276_, _02275_, _02248_);
  and _33811_ (_02277_, _02276_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _33812_ (_02278_, _02277_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _33813_ (_02279_, _02278_, _02250_);
  and _33814_ (_02280_, _02279_, _02271_);
  and _33815_ (_02281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _33816_ (_02282_, _02281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _33817_ (_02283_, _02236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _33818_ (_02284_, _02262_, _02248_);
  and _33819_ (_02285_, _02284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or _33820_ (_02286_, _02285_, _02250_);
  and _33821_ (_02287_, _02286_, _02283_);
  or _33822_ (_02288_, _02287_, _02282_);
  or _33823_ (_02289_, _02288_, _02280_);
  nor _33824_ (_02290_, _02289_, _02270_);
  and _33825_ (_02291_, _25556_, _24174_);
  and _33826_ (_02292_, _02291_, _24179_);
  nor _33827_ (_02293_, _02292_, _02290_);
  and _33828_ (_02294_, _25602_, _24174_);
  nor _33829_ (_02295_, _02294_, rst);
  and _33830_ (_22652_, _02295_, _02293_);
  and _33831_ (_02296_, _02232_, _23996_);
  and _33832_ (_02297_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or _33833_ (_27021_, _02297_, _02296_);
  and _33834_ (_02298_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _33835_ (_02299_, _01814_, _23989_);
  not _33836_ (_02300_, _01816_);
  not _33837_ (_02301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _33838_ (_02302_, _01823_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _33839_ (_02303_, _02302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _33840_ (_02304_, _02209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _33841_ (_02305_, _02304_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _33842_ (_02306_, _02305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _33843_ (_02307_, _02306_, _02303_);
  nand _33844_ (_02308_, _02307_, _02205_);
  nor _33845_ (_02309_, _02308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _33846_ (_02310_, _02309_, _02301_);
  and _33847_ (_02311_, _02309_, _02301_);
  or _33848_ (_02312_, _02311_, _02310_);
  and _33849_ (_02313_, _02312_, _02198_);
  or _33850_ (_02314_, _01826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not _33851_ (_02315_, _01827_);
  and _33852_ (_02316_, _01829_, _02315_);
  and _33853_ (_02317_, _02316_, _02314_);
  and _33854_ (_02318_, _02210_, _02303_);
  or _33855_ (_02319_, _02318_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not _33856_ (_02320_, _02219_);
  and _33857_ (_02321_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _33858_ (_02322_, _02210_, _02321_);
  nor _33859_ (_02323_, _02322_, _02320_);
  and _33860_ (_02324_, _02323_, _02319_);
  or _33861_ (_02325_, _02324_, _02317_);
  or _33862_ (_02326_, _02325_, _02313_);
  or _33863_ (_02328_, _02326_, _01814_);
  and _33864_ (_02329_, _02328_, _02300_);
  and _33865_ (_02330_, _02329_, _02299_);
  or _33866_ (_02331_, _02330_, _02298_);
  and _33867_ (_22653_, _02331_, _22731_);
  and _33868_ (_02332_, _02232_, _24134_);
  and _33869_ (_02333_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or _33870_ (_27020_, _02333_, _02332_);
  and _33871_ (_02334_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _33872_ (_02335_, _02040_, _24089_);
  or _33873_ (_22654_, _02335_, _02334_);
  and _33874_ (_02336_, _02093_, _23548_);
  and _33875_ (_02337_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _33876_ (_22655_, _02337_, _02336_);
  and _33877_ (_02338_, _02039_, _24297_);
  not _33878_ (_02339_, _02338_);
  and _33879_ (_02340_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and _33880_ (_02341_, _02338_, _24134_);
  or _33881_ (_22656_, _02341_, _02340_);
  and _33882_ (_02343_, _02093_, _24219_);
  and _33883_ (_02344_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _33884_ (_22657_, _02344_, _02343_);
  and _33885_ (_02345_, _02232_, _24219_);
  and _33886_ (_02346_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or _33887_ (_22658_, _02346_, _02345_);
  and _33888_ (_02347_, _24017_, _23583_);
  and _33889_ (_02348_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or _33890_ (_22659_, _02348_, _02347_);
  or _33891_ (_02349_, _02019_, _26756_);
  or _33892_ (_02350_, _02349_, _23840_);
  or _33893_ (_02351_, _02021_, _02015_);
  and _33894_ (_02352_, _26760_, _23708_);
  or _33895_ (_02353_, _02352_, _23841_);
  or _33896_ (_02354_, _02353_, _02351_);
  or _33897_ (_02355_, _02354_, _02350_);
  and _33898_ (_02356_, _02355_, _22737_);
  and _33899_ (_02357_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _33900_ (_02358_, _26675_);
  and _33901_ (_02359_, _02358_, _02003_);
  and _33902_ (_02360_, _02351_, _26573_);
  or _33903_ (_02361_, _02360_, _02359_);
  or _33904_ (_02362_, _02361_, _02357_);
  or _33905_ (_02363_, _02362_, _02356_);
  and _33906_ (_26848_[1], _02363_, _22731_);
  and _33907_ (_02364_, _24365_, _24297_);
  and _33908_ (_02365_, _02364_, _23583_);
  not _33909_ (_02366_, _02364_);
  and _33910_ (_02367_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _33911_ (_27208_, _02367_, _02365_);
  and _33912_ (_02368_, _24408_, _24159_);
  and _33913_ (_02369_, _02368_, _24051_);
  not _33914_ (_02370_, _02368_);
  and _33915_ (_02371_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or _33916_ (_27152_, _02371_, _02369_);
  and _33917_ (_02372_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and _33918_ (_02373_, _02338_, _23996_);
  or _33919_ (_22660_, _02373_, _02372_);
  and _33920_ (_02374_, _26743_, _26736_);
  and _33921_ (_02375_, _26698_, _23779_);
  or _33922_ (_02376_, _01992_, _26760_);
  or _33923_ (_02377_, _02376_, _02375_);
  or _33924_ (_02378_, _23805_, _23800_);
  and _33925_ (_02379_, _02378_, _23803_);
  or _33926_ (_02380_, _02379_, _26724_);
  or _33927_ (_02381_, _02380_, _02377_);
  nor _33928_ (_02382_, _02381_, _02015_);
  nand _33929_ (_02383_, _02382_, _02374_);
  or _33930_ (_02384_, _02022_, _26721_);
  or _33931_ (_02385_, _23841_, _23839_);
  and _33932_ (_02386_, _23772_, _23824_);
  or _33933_ (_02387_, _02386_, _02385_);
  or _33934_ (_02388_, _02387_, _02384_);
  or _33935_ (_02389_, _26691_, _23830_);
  or _33936_ (_02390_, _02389_, _23828_);
  or _33937_ (_02391_, _02390_, _02388_);
  or _33938_ (_02392_, _02391_, _02350_);
  or _33939_ (_02393_, _02392_, _02383_);
  and _33940_ (_02394_, _02393_, _22737_);
  and _33941_ (_02395_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _33942_ (_02396_, _26595_, _23708_);
  and _33943_ (_02397_, _02396_, _26573_);
  and _33944_ (_02398_, _26581_, _26573_);
  or _33945_ (_02399_, _02398_, _02359_);
  or _33946_ (_02400_, _02399_, _02397_);
  or _33947_ (_02401_, _02400_, _02395_);
  or _33948_ (_02402_, _02401_, _02394_);
  and _33949_ (_26853_, _02402_, _22731_);
  and _33950_ (_02403_, _02368_, _23583_);
  and _33951_ (_02404_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or _33952_ (_22661_, _02404_, _02403_);
  and _33953_ (_02405_, _02368_, _23548_);
  and _33954_ (_02406_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or _33955_ (_22662_, _02406_, _02405_);
  and _33956_ (_02407_, _02045_, _23887_);
  and _33957_ (_02408_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _33958_ (_22663_, _02408_, _02407_);
  and _33959_ (_02409_, _02368_, _24219_);
  and _33960_ (_02410_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or _33961_ (_22664_, _02410_, _02409_);
  and _33962_ (_02411_, _02065_, _23548_);
  and _33963_ (_02412_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or _33964_ (_22665_, _02412_, _02411_);
  and _33965_ (_02413_, _24408_, _24297_);
  and _33966_ (_02414_, _02413_, _24134_);
  not _33967_ (_02415_, _02413_);
  and _33968_ (_02416_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _33969_ (_22666_, _02416_, _02414_);
  and _33970_ (_02417_, _02413_, _24089_);
  and _33971_ (_02418_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _33972_ (_27149_, _02418_, _02417_);
  and _33973_ (_02419_, _02413_, _23887_);
  and _33974_ (_02420_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _33975_ (_27148_, _02420_, _02419_);
  and _33976_ (_02421_, _24497_, _24134_);
  and _33977_ (_02422_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or _33978_ (_27245_, _02422_, _02421_);
  or _33979_ (_02423_, _02386_, _02021_);
  or _33980_ (_02424_, _02423_, _02389_);
  or _33981_ (_02425_, _02424_, _02383_);
  and _33982_ (_02426_, _02425_, _22737_);
  and _33983_ (_02427_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _33984_ (_02428_, _02427_, _02400_);
  or _33985_ (_02429_, _02428_, _02426_);
  and _33986_ (_26848_[0], _02429_, _22731_);
  and _33987_ (_02430_, _24497_, _24051_);
  and _33988_ (_02431_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or _33989_ (_22667_, _02431_, _02430_);
  and _33990_ (_02432_, _25413_, _24016_);
  and _33991_ (_02433_, _02432_, _23996_);
  not _33992_ (_02434_, _02432_);
  and _33993_ (_02435_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  or _33994_ (_22668_, _02435_, _02433_);
  and _33995_ (_02436_, _02413_, _23548_);
  and _33996_ (_02437_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _33997_ (_22669_, _02437_, _02436_);
  and _33998_ (_02438_, _24188_, _22868_);
  and _33999_ (_02439_, _02438_, _24533_);
  and _34000_ (_02440_, _02439_, _22731_);
  and _34001_ (_02441_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _34002_ (_02442_, _02273_, _02253_);
  and _34003_ (_02443_, _02442_, _02271_);
  and _34004_ (_02444_, _02266_, _02237_);
  nor _34005_ (_02445_, _02444_, _02443_);
  and _34006_ (_02446_, _02445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _34007_ (_02447_, _02445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _34008_ (_02448_, _02447_, _02446_);
  nor _34009_ (_02449_, _02448_, _02292_);
  not _34010_ (_02450_, _24126_);
  and _34011_ (_02451_, _02292_, _02450_);
  or _34012_ (_02452_, _02451_, _02449_);
  and _34013_ (_02453_, _02452_, _02295_);
  or _34014_ (_22670_, _02453_, _02441_);
  and _34015_ (_02455_, _24408_, _24016_);
  and _34016_ (_02456_, _02455_, _24134_);
  not _34017_ (_02458_, _02455_);
  and _34018_ (_02459_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _34019_ (_22671_, _02459_, _02456_);
  and _34020_ (_02460_, _02455_, _24089_);
  and _34021_ (_02461_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _34022_ (_22672_, _02461_, _02460_);
  and _34023_ (_02462_, _02232_, _23583_);
  and _34024_ (_02463_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or _34025_ (_22673_, _02463_, _02462_);
  and _34026_ (_02465_, _02232_, _23887_);
  and _34027_ (_02467_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or _34028_ (_22674_, _02467_, _02465_);
  and _34029_ (_02468_, _02232_, _23548_);
  and _34030_ (_02469_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or _34031_ (_27019_, _02469_, _02468_);
  and _34032_ (_02470_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and _34033_ (_02471_, _02338_, _23887_);
  or _34034_ (_22675_, _02471_, _02470_);
  and _34035_ (_02472_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and _34036_ (_02473_, _02338_, _23548_);
  or _34037_ (_27025_, _02473_, _02472_);
  nand _34038_ (_02474_, _26406_, _23531_);
  or _34039_ (_02475_, _23531_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _34040_ (_02476_, _02475_, _22731_);
  and _34041_ (_22676_, _02476_, _02474_);
  and _34042_ (_02478_, _24899_, _24496_);
  and _34043_ (_02479_, _02478_, _24134_);
  not _34044_ (_02480_, _02478_);
  and _34045_ (_02481_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _34046_ (_22677_, _02481_, _02479_);
  and _34047_ (_02483_, _02455_, _23887_);
  and _34048_ (_02484_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _34049_ (_22678_, _02484_, _02483_);
  and _34050_ (_02485_, _02478_, _23996_);
  and _34051_ (_02486_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or _34052_ (_22679_, _02486_, _02485_);
  and _34053_ (_02488_, _24349_, _24006_);
  and _34054_ (_02489_, _02488_, _24089_);
  not _34055_ (_02490_, _02488_);
  and _34056_ (_02491_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or _34057_ (_22680_, _02491_, _02489_);
  and _34058_ (_02492_, _02364_, _24089_);
  and _34059_ (_02494_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _34060_ (_22681_, _02494_, _02492_);
  nand _34061_ (_02495_, _24299_, _22847_);
  and _34062_ (_02497_, _02495_, _24003_);
  and _34063_ (_02498_, _02497_, _24159_);
  and _34064_ (_02499_, _02498_, _24089_);
  not _34065_ (_02500_, _02498_);
  and _34066_ (_02501_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or _34067_ (_22682_, _02501_, _02499_);
  and _34068_ (_02502_, _24496_, _23941_);
  and _34069_ (_02503_, _02502_, _24219_);
  not _34070_ (_02504_, _02502_);
  and _34071_ (_02505_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _34072_ (_27248_, _02505_, _02503_);
  and _34073_ (_02507_, _02455_, _23548_);
  and _34074_ (_02508_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _34075_ (_27145_, _02508_, _02507_);
  and _34076_ (_02509_, _02498_, _23583_);
  and _34077_ (_02511_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _34078_ (_22683_, _02511_, _02509_);
  and _34079_ (_02512_, _24004_, _22977_);
  and _34080_ (_02513_, _02512_, _24146_);
  not _34081_ (_02514_, _02513_);
  and _34082_ (_02515_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and _34083_ (_02516_, _02513_, _24089_);
  or _34084_ (_22684_, _02516_, _02515_);
  and _34085_ (_02517_, _24408_, _24236_);
  and _34086_ (_02518_, _02517_, _23996_);
  not _34087_ (_02519_, _02517_);
  and _34088_ (_02520_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or _34089_ (_27143_, _02520_, _02518_);
  and _34090_ (_02521_, _02517_, _24051_);
  and _34091_ (_02522_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or _34092_ (_22685_, _02522_, _02521_);
  and _34093_ (_02523_, _02517_, _23583_);
  and _34094_ (_02524_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or _34095_ (_22686_, _02524_, _02523_);
  and _34096_ (_02525_, _24889_, _23583_);
  and _34097_ (_02526_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _34098_ (_22687_, _02526_, _02525_);
  and _34099_ (_02527_, _24698_, _24543_);
  and _34100_ (_02528_, _02527_, _24594_);
  nand _34101_ (_02530_, _02528_, _23504_);
  or _34102_ (_02531_, _02528_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _34103_ (_02532_, _25227_, _24628_);
  not _34104_ (_02534_, _02532_);
  and _34105_ (_02535_, _02534_, _02531_);
  and _34106_ (_02536_, _02535_, _02530_);
  nor _34107_ (_02537_, _02534_, _24126_);
  or _34108_ (_02539_, _02537_, _02536_);
  and _34109_ (_22690_, _02539_, _22731_);
  and _34110_ (_02540_, _02527_, _24607_);
  nand _34111_ (_02541_, _02540_, _23504_);
  or _34112_ (_02542_, _02540_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _34113_ (_02543_, _02542_, _02534_);
  and _34114_ (_02544_, _02543_, _02541_);
  nor _34115_ (_02545_, _02534_, _24043_);
  or _34116_ (_02546_, _02545_, _02544_);
  and _34117_ (_22691_, _02546_, _22731_);
  and _34118_ (_02548_, _24638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _34119_ (_02549_, _02548_, _24637_);
  and _34120_ (_02550_, _02549_, _02527_);
  not _34121_ (_02551_, _02527_);
  or _34122_ (_02552_, _02551_, _24643_);
  and _34123_ (_02553_, _02552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _34124_ (_02555_, _02553_, _02532_);
  or _34125_ (_02556_, _02555_, _02550_);
  nand _34126_ (_02557_, _02532_, _24082_);
  and _34127_ (_02558_, _02557_, _22731_);
  and _34128_ (_22692_, _02558_, _02556_);
  and _34129_ (_02560_, _02527_, _24533_);
  nand _34130_ (_02561_, _02560_, _23504_);
  or _34131_ (_02562_, _02560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _34132_ (_02563_, _02562_, _02534_);
  and _34133_ (_02564_, _02563_, _02561_);
  and _34134_ (_02565_, _02532_, _23577_);
  or _34135_ (_02566_, _02565_, _02564_);
  and _34136_ (_22693_, _02566_, _22731_);
  nor _34137_ (_02568_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _34138_ (_02569_, _02568_);
  nor _34139_ (_02570_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _34140_ (_02571_, _02570_, _02569_);
  and _34141_ (_02572_, _02571_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _34142_ (_02573_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _34143_ (_02574_, _02571_, _02573_);
  or _34144_ (_02576_, _02574_, _02572_);
  or _34145_ (_02577_, _02576_, _02527_);
  not _34146_ (_02578_, _24562_);
  nor _34147_ (_02580_, _02578_, _23504_);
  or _34148_ (_02581_, _24562_, _02573_);
  nand _34149_ (_02582_, _02581_, _02527_);
  or _34150_ (_02583_, _02582_, _02580_);
  and _34151_ (_02584_, _02583_, _02577_);
  or _34152_ (_02585_, _02584_, _02532_);
  or _34153_ (_02586_, _02534_, _23880_);
  and _34154_ (_02587_, _02586_, _22731_);
  and _34155_ (_22694_, _02587_, _02585_);
  or _34156_ (_02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _34157_ (_02589_, _02588_, _02527_);
  and _34158_ (_02590_, _24177_, _24531_);
  not _34159_ (_02591_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _34160_ (_02592_, _24177_, _02591_);
  nand _34161_ (_02593_, _02592_, _02527_);
  or _34162_ (_02594_, _02593_, _02590_);
  and _34163_ (_02595_, _02594_, _02589_);
  or _34164_ (_02596_, _02595_, _02532_);
  nand _34165_ (_02597_, _02532_, _23542_);
  and _34166_ (_02598_, _02597_, _22731_);
  and _34167_ (_22695_, _02598_, _02596_);
  and _34168_ (_02599_, _24577_, _24531_);
  not _34169_ (_02600_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _34170_ (_02601_, _24577_, _02600_);
  nand _34171_ (_02602_, _02601_, _02527_);
  or _34172_ (_02603_, _02602_, _02599_);
  not _34173_ (_02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _34174_ (_02605_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _34175_ (_02606_, _02605_, _02568_);
  and _34176_ (_02607_, _02606_, _02570_);
  or _34177_ (_02608_, _02607_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _34178_ (_02609_, _02608_, _02527_);
  and _34179_ (_02610_, _02609_, _02603_);
  or _34180_ (_02611_, _02610_, _02532_);
  nand _34181_ (_02612_, _02532_, _24210_);
  and _34182_ (_02613_, _02612_, _22731_);
  and _34183_ (_22696_, _02613_, _02611_);
  nand _34184_ (_02614_, _02294_, _23989_);
  nor _34185_ (_02615_, _02283_, _02237_);
  and _34186_ (_02616_, _25557_, _24174_);
  or _34187_ (_02617_, _02616_, _02615_);
  and _34188_ (_02618_, _02617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or _34189_ (_02619_, _02284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _34190_ (_02620_, _02263_, _02248_);
  nor _34191_ (_02621_, _02620_, _02615_);
  and _34192_ (_02622_, _02621_, _02619_);
  and _34193_ (_02623_, _02620_, _02283_);
  and _34194_ (_02624_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _34195_ (_02625_, _02624_, _02622_);
  nor _34196_ (_02626_, _02625_, _02616_);
  or _34197_ (_02627_, _02626_, _02618_);
  or _34198_ (_02628_, _02627_, _02294_);
  and _34199_ (_02629_, _02628_, _22731_);
  and _34200_ (_22697_, _02629_, _02614_);
  or _34201_ (_02630_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _34202_ (_02631_, _02630_, _22731_);
  nand _34203_ (_02632_, _02071_, _24126_);
  and _34204_ (_22698_, _02632_, _02631_);
  or _34205_ (_02633_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _34206_ (_02634_, _02633_, _22731_);
  nand _34207_ (_02635_, _02071_, _24043_);
  and _34208_ (_22699_, _02635_, _02634_);
  or _34209_ (_02636_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _34210_ (_02637_, _02636_, _22731_);
  or _34211_ (_02638_, _02074_, _23577_);
  and _34212_ (_22700_, _02638_, _02637_);
  or _34213_ (_02639_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _34214_ (_02640_, _02639_, _22731_);
  nand _34215_ (_02641_, _02071_, _23542_);
  and _34216_ (_22701_, _02641_, _02640_);
  nand _34217_ (_02642_, _02071_, _24210_);
  or _34218_ (_02643_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _34219_ (_02644_, _02643_, _22731_);
  and _34220_ (_22702_, _02644_, _02642_);
  not _34221_ (_02645_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _34222_ (_02646_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _34223_ (_02647_, _02646_, _02568_);
  and _34224_ (_02648_, _02569_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _34225_ (_02649_, _02648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _34226_ (_02650_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _34227_ (_02651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _34228_ (_02652_, _02651_, _02650_);
  and _34229_ (_02653_, _02652_, _02649_);
  nor _34230_ (_02654_, _02653_, _02647_);
  nor _34231_ (_02655_, _02654_, _02645_);
  and _34232_ (_02656_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _34233_ (_02657_, _02656_, _02655_);
  and _34234_ (_02658_, _25227_, _24182_);
  nor _34235_ (_02659_, _02658_, _02657_);
  not _34236_ (_02660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _34237_ (_02661_, _02660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _34238_ (_02662_, _02661_, _02569_);
  and _34239_ (_02663_, _02662_, _02658_);
  or _34240_ (_02664_, _02663_, _02659_);
  and _34241_ (_22703_, _02664_, _22731_);
  and _34242_ (_02665_, _02658_, _02569_);
  nand _34243_ (_02666_, _02665_, _23989_);
  and _34244_ (_02668_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  not _34245_ (_02669_, _02654_);
  and _34246_ (_02670_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _34247_ (_02671_, _02670_, _02668_);
  or _34248_ (_02672_, _02671_, _02658_);
  and _34249_ (_02673_, _02672_, _22731_);
  and _34250_ (_22704_, _02673_, _02666_);
  not _34251_ (_02674_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _34252_ (_02675_, _02658_, _02660_);
  and _34253_ (_02676_, _02675_, _02674_);
  and _34254_ (_02677_, _02676_, _25554_);
  and _34255_ (_02678_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _34256_ (_02679_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _34257_ (_02680_, _02679_, _02678_);
  nor _34258_ (_02681_, _02680_, _02658_);
  and _34259_ (_02682_, _02665_, _02450_);
  or _34260_ (_02683_, _02682_, _02681_);
  or _34261_ (_02684_, _02683_, _02677_);
  and _34262_ (_22705_, _02684_, _22731_);
  and _34263_ (_02685_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _34264_ (_02686_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _34265_ (_02687_, _02686_, _02685_);
  nor _34266_ (_02688_, _02687_, _02658_);
  not _34267_ (_02689_, _24043_);
  and _34268_ (_02690_, _02665_, _02689_);
  and _34269_ (_02691_, _02658_, _02568_);
  and _34270_ (_02692_, _02691_, _02450_);
  or _34271_ (_02693_, _02692_, _02690_);
  or _34272_ (_02694_, _02693_, _02688_);
  and _34273_ (_22706_, _02694_, _22731_);
  and _34274_ (_02695_, _02676_, _02689_);
  and _34275_ (_02696_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _34276_ (_02697_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _34277_ (_02698_, _02697_, _02696_);
  nor _34278_ (_02699_, _02698_, _02658_);
  not _34279_ (_02700_, _24082_);
  and _34280_ (_02701_, _02665_, _02700_);
  or _34281_ (_02702_, _02701_, _02699_);
  or _34282_ (_02703_, _02702_, _02695_);
  and _34283_ (_22707_, _02703_, _22731_);
  and _34284_ (_02704_, _02665_, _23577_);
  and _34285_ (_02705_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _34286_ (_02706_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _34287_ (_02707_, _02706_, _02705_);
  nor _34288_ (_02708_, _02707_, _02658_);
  and _34289_ (_02709_, _02691_, _02700_);
  or _34290_ (_02710_, _02709_, _02708_);
  or _34291_ (_02711_, _02710_, _02704_);
  and _34292_ (_22708_, _02711_, _22731_);
  and _34293_ (_02712_, _02676_, _23577_);
  and _34294_ (_02713_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _34295_ (_02714_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _34296_ (_02715_, _02714_, _02713_);
  nor _34297_ (_02716_, _02715_, _02658_);
  and _34298_ (_02717_, _02665_, _23880_);
  or _34299_ (_02718_, _02717_, _02716_);
  or _34300_ (_02720_, _02718_, _02712_);
  and _34301_ (_22709_, _02720_, _22731_);
  and _34302_ (_02722_, _02676_, _23880_);
  and _34303_ (_02723_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _34304_ (_02724_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _34305_ (_02726_, _02724_, _02723_);
  nor _34306_ (_02727_, _02726_, _02658_);
  not _34307_ (_02728_, _23542_);
  and _34308_ (_02729_, _02665_, _02728_);
  or _34309_ (_02730_, _02729_, _02727_);
  or _34310_ (_02731_, _02730_, _02722_);
  and _34311_ (_22710_, _02731_, _22731_);
  and _34312_ (_02732_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _34313_ (_02733_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _34314_ (_02734_, _02733_, _02732_);
  nor _34315_ (_02735_, _02734_, _02658_);
  and _34316_ (_02737_, _02665_, _24671_);
  or _34317_ (_02738_, _02737_, _02735_);
  and _34318_ (_02739_, _02691_, _02728_);
  or _34319_ (_02740_, _02739_, _02738_);
  and _34320_ (_22711_, _02740_, _22731_);
  or _34321_ (_02742_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _34322_ (_02743_, _02647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _34323_ (_02744_, _02743_, _02653_);
  and _34324_ (_02745_, _02744_, _02742_);
  nor _34325_ (_02746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor _34326_ (_02748_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _34327_ (_02749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _34328_ (_02750_, _02749_, _02748_);
  and _34329_ (_02752_, _02750_, _02746_);
  nor _34330_ (_02753_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _34331_ (_02754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _34332_ (_02755_, _02754_, _02753_);
  and _34333_ (_02756_, _02755_, _02647_);
  and _34334_ (_02757_, _02756_, _02752_);
  and _34335_ (_02758_, _02757_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _34336_ (_02759_, _02758_, _02745_);
  nor _34337_ (_02760_, _02759_, _02658_);
  and _34338_ (_02761_, _02691_, _24671_);
  or _34339_ (_02762_, _02761_, _02760_);
  and _34340_ (_22712_, _02762_, _22731_);
  and _34341_ (_02764_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and _34342_ (_02765_, _02338_, _24089_);
  or _34343_ (_22713_, _02765_, _02764_);
  and _34344_ (_02767_, _25413_, _24349_);
  and _34345_ (_02768_, _02767_, _23996_);
  not _34346_ (_02769_, _02767_);
  and _34347_ (_02771_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _34348_ (_27175_, _02771_, _02768_);
  and _34349_ (_02772_, _02488_, _23887_);
  and _34350_ (_02774_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or _34351_ (_22714_, _02774_, _02772_);
  and _34352_ (_02775_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and _34353_ (_02776_, _02338_, _23583_);
  or _34354_ (_27026_, _02776_, _02775_);
  and _34355_ (_02777_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _34356_ (_02778_, _02777_, _02569_);
  not _34357_ (_02779_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _34358_ (_02780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _02779_);
  not _34359_ (_02782_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _34360_ (_02783_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _02782_);
  and _34361_ (_02784_, _02783_, _02780_);
  and _34362_ (_02785_, _02784_, _02778_);
  not _34363_ (_02786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _34364_ (_02787_, _02786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _34365_ (_02789_, _02568_, _02600_);
  and _34366_ (_02790_, _02789_, _02787_);
  and _34367_ (_02792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _34368_ (_02793_, _02792_, _02569_);
  nor _34369_ (_02794_, _02793_, _02790_);
  nor _34370_ (_02795_, _02794_, _02778_);
  or _34371_ (_02796_, _02795_, _02785_);
  and _34372_ (_02798_, _02568_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _34373_ (_02799_, _02798_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or _34374_ (_02800_, _02799_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _34375_ (_02801_, _02800_, _02796_);
  nor _34376_ (_02802_, _02799_, _02785_);
  or _34377_ (_02803_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _34378_ (_02804_, _02803_, _02080_);
  and _34379_ (_02806_, _02804_, _02801_);
  or _34380_ (_22715_, _02806_, _02079_);
  and _34381_ (_22716_, t0_i, _22731_);
  and _34382_ (_02807_, _02498_, _23996_);
  and _34383_ (_02809_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _34384_ (_22717_, _02809_, _02807_);
  not _34385_ (_02810_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not _34386_ (_02811_, _02802_);
  nor _34387_ (_02812_, _02811_, _02795_);
  nor _34388_ (_02813_, _02812_, _02810_);
  or _34389_ (_02814_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _34390_ (_02815_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _02810_);
  or _34391_ (_02816_, _02815_, _02802_);
  and _34392_ (_02817_, _02816_, _22731_);
  and _34393_ (_22718_, _02817_, _02814_);
  and _34394_ (_02818_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _34395_ (_02819_, _02811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not _34396_ (_02820_, _02778_);
  nor _34397_ (_02821_, _02784_, _02820_);
  and _34398_ (_02823_, _02821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor _34399_ (_02824_, _02778_, _02790_);
  or _34400_ (_02825_, _02824_, _02823_);
  nor _34401_ (_02826_, _02793_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor _34402_ (_02827_, _02826_, _02799_);
  and _34403_ (_02829_, _02827_, _02825_);
  or _34404_ (_02830_, _02829_, _02819_);
  and _34405_ (_02831_, _02830_, _02080_);
  or _34406_ (_22719_, _02831_, _02818_);
  and _34407_ (_02832_, _02488_, _23548_);
  and _34408_ (_02833_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or _34409_ (_22720_, _02833_, _02832_);
  and _34410_ (_02834_, _02498_, _24134_);
  and _34411_ (_02835_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _34412_ (_22721_, _02835_, _02834_);
  and _34413_ (_02836_, _02039_, _24016_);
  not _34414_ (_02837_, _02836_);
  and _34415_ (_02838_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and _34416_ (_02839_, _02836_, _24134_);
  or _34417_ (_27024_, _02839_, _02838_);
  not _34418_ (_02840_, _02812_);
  or _34419_ (_02841_, _02840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _34420_ (_02842_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _34421_ (_02844_, _02842_, _02080_);
  and _34422_ (_02845_, _02844_, _02841_);
  or _34423_ (_22722_, _02845_, _02085_);
  and _34424_ (_02846_, _02478_, _23583_);
  and _34425_ (_02847_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or _34426_ (_27247_, _02847_, _02846_);
  and _34427_ (_02848_, _02517_, _23887_);
  and _34428_ (_02849_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or _34429_ (_22723_, _02849_, _02848_);
  and _34430_ (_02851_, _02432_, _24051_);
  and _34431_ (_02852_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  or _34432_ (_22724_, _02852_, _02851_);
  and _34433_ (_02854_, _02784_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _34434_ (_02855_, _02854_, _02794_);
  or _34435_ (_02856_, _02855_, _02812_);
  and _34436_ (_02857_, _02856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _34437_ (_02858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _02810_);
  nand _34438_ (_02859_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _34439_ (_02860_, _02859_, _02802_);
  or _34440_ (_02861_, _02860_, _02858_);
  or _34441_ (_02862_, _02861_, _02857_);
  and _34442_ (_22725_, _02862_, _22731_);
  nor _34443_ (_02863_, _02793_, _02778_);
  or _34444_ (_02865_, _02863_, _02810_);
  or _34445_ (_02866_, _02865_, _02782_);
  and _34446_ (_02867_, _02778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _34447_ (_02868_, _02867_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _34448_ (_02869_, _02868_, _22731_);
  and _34449_ (_22726_, _02869_, _02866_);
  nand _34450_ (_02870_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22731_);
  nor _34451_ (_02871_, _02870_, _02813_);
  or _34452_ (_02872_, _02855_, _02811_);
  and _34453_ (_02873_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _34454_ (_02874_, _02873_, _02872_);
  or _34455_ (_22727_, _02874_, _02871_);
  and _34456_ (_02875_, _02865_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _34457_ (_02876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _34458_ (_02877_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _34459_ (_02879_, _02877_, _02876_);
  and _34460_ (_02880_, _02879_, _02867_);
  or _34461_ (_02881_, _02880_, _02875_);
  and _34462_ (_22728_, _02881_, _22731_);
  and _34463_ (_02882_, _02497_, _24297_);
  and _34464_ (_02883_, _02882_, _24134_);
  not _34465_ (_02884_, _02882_);
  and _34466_ (_02885_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _34467_ (_22729_, _02885_, _02883_);
  or _34468_ (_02886_, _02649_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _34469_ (_02887_, _02649_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _34470_ (_02888_, _02887_, rst);
  nand _34471_ (_02889_, _02888_, _02886_);
  nor _34472_ (_22730_, _02889_, _02658_);
  and _34473_ (_02890_, _24408_, _24349_);
  and _34474_ (_02891_, _02890_, _23996_);
  not _34475_ (_02892_, _02890_);
  and _34476_ (_02893_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or _34477_ (_22739_, _02893_, _02891_);
  and _34478_ (_02894_, _02478_, _24089_);
  and _34479_ (_02895_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or _34480_ (_22743_, _02895_, _02894_);
  and _34481_ (_02896_, _02876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _34482_ (_02897_, _02896_, _02779_);
  and _34483_ (_02898_, _02867_, _02897_);
  or _34484_ (_02899_, _02898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not _34485_ (_02900_, rxd_i);
  nand _34486_ (_02901_, _02898_, _02900_);
  and _34487_ (_02902_, _02901_, _22731_);
  and _34488_ (_22748_, _02902_, _02899_);
  and _34489_ (_02903_, _02882_, _24051_);
  and _34490_ (_02904_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _34491_ (_26986_, _02904_, _02903_);
  or _34492_ (_02905_, _02887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _34493_ (_02906_, _02887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _34494_ (_02907_, _02906_, rst);
  nand _34495_ (_02908_, _02907_, _02905_);
  nor _34496_ (_22754_, _02908_, _02658_);
  nor _34497_ (_02909_, _02906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _34498_ (_02910_, _02906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _34499_ (_02911_, _02910_, _02909_);
  nand _34500_ (_02912_, _02911_, _22731_);
  nor _34501_ (_22756_, _02912_, _02658_);
  or _34502_ (_02913_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _34503_ (_02914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _02810_);
  or _34504_ (_02915_, _02914_, _02802_);
  and _34505_ (_02916_, _02915_, _22731_);
  and _34506_ (_22765_, _02916_, _02913_);
  and _34507_ (_02917_, _02882_, _24089_);
  and _34508_ (_02918_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _34509_ (_22770_, _02918_, _02917_);
  and _34510_ (_02919_, _02478_, _24051_);
  and _34511_ (_02920_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _34512_ (_22787_, _02920_, _02919_);
  and _34513_ (_02921_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  and _34514_ (_02922_, _02836_, _23996_);
  or _34515_ (_22798_, _02922_, _02921_);
  and _34516_ (_02923_, _02865_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor _34517_ (_02925_, _02896_, _02820_);
  or _34518_ (_02926_, _02925_, _02923_);
  and _34519_ (_02927_, _02876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _34520_ (_02928_, _02927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _34521_ (_02929_, _02928_, _22731_);
  and _34522_ (_22807_, _02929_, _02926_);
  and _34523_ (_02930_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _34524_ (_22819_, _02930_, _02818_);
  and _34525_ (_02931_, _02498_, _24219_);
  and _34526_ (_02932_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _34527_ (_27007_, _02932_, _02931_);
  and _34528_ (_02934_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _34529_ (_02935_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _34530_ (_22842_, _02935_, _02934_);
  and _34531_ (_02936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _34532_ (_02937_, _02936_, _02858_);
  and _34533_ (_22848_, _02937_, _22731_);
  and _34534_ (_02938_, _02890_, _24134_);
  and _34535_ (_02939_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or _34536_ (_22860_, _02939_, _02938_);
  and _34537_ (_02940_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _34538_ (_02941_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _34539_ (_22870_, _02941_, _02940_);
  and _34540_ (_02942_, _02882_, _23996_);
  and _34541_ (_02943_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _34542_ (_22873_, _02943_, _02942_);
  and _34543_ (_02944_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and _34544_ (_02945_, _02836_, _23887_);
  or _34545_ (_22879_, _02945_, _02944_);
  or _34546_ (_02946_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _34547_ (_02947_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _02810_);
  or _34548_ (_02948_, _02947_, _02802_);
  and _34549_ (_02949_, _02948_, _22731_);
  and _34550_ (_22883_, _02949_, _02946_);
  or _34551_ (_02950_, _02840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _34552_ (_02951_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _34553_ (_02952_, _02951_, _02080_);
  and _34554_ (_02953_, _02952_, _02950_);
  or _34555_ (_22889_, _02953_, _02083_);
  or _34556_ (_02954_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _34557_ (_02955_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _02810_);
  or _34558_ (_02956_, _02955_, _02802_);
  and _34559_ (_02957_, _02956_, _22731_);
  and _34560_ (_22892_, _02957_, _02954_);
  or _34561_ (_02958_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _34562_ (_02959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _02810_);
  or _34563_ (_02960_, _02959_, _02802_);
  and _34564_ (_02961_, _02960_, _22731_);
  and _34565_ (_22895_, _02961_, _02958_);
  and _34566_ (_02962_, _02890_, _24089_);
  and _34567_ (_02963_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or _34568_ (_22915_, _02963_, _02962_);
  and _34569_ (_02964_, _24476_, _24236_);
  and _34570_ (_02965_, _02964_, _23996_);
  not _34571_ (_02966_, _02964_);
  and _34572_ (_02967_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _34573_ (_27187_, _02967_, _02965_);
  and _34574_ (_02968_, _02890_, _23887_);
  and _34575_ (_02969_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or _34576_ (_22929_, _02969_, _02968_);
  and _34577_ (_02970_, _24301_, _24016_);
  and _34578_ (_02971_, _02970_, _23583_);
  not _34579_ (_02972_, _02970_);
  and _34580_ (_02973_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or _34581_ (_22939_, _02973_, _02971_);
  and _34582_ (_02974_, _24497_, _23583_);
  and _34583_ (_02975_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or _34584_ (_22944_, _02975_, _02974_);
  and _34585_ (_02976_, _02882_, _24219_);
  and _34586_ (_02977_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _34587_ (_22955_, _02977_, _02976_);
  and _34588_ (_02978_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and _34589_ (_02979_, _02836_, _24089_);
  or _34590_ (_22959_, _02979_, _02978_);
  and _34591_ (_02980_, _02497_, _24016_);
  and _34592_ (_02981_, _02980_, _23996_);
  not _34593_ (_02982_, _02980_);
  and _34594_ (_02983_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _34595_ (_23014_, _02983_, _02981_);
  and _34596_ (_02984_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and _34597_ (_02985_, _02836_, _23583_);
  or _34598_ (_23021_, _02985_, _02984_);
  and _34599_ (_02986_, _02882_, _23548_);
  and _34600_ (_02987_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _34601_ (_23046_, _02987_, _02986_);
  and _34602_ (_02988_, _02882_, _23887_);
  and _34603_ (_02989_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _34604_ (_23077_, _02989_, _02988_);
  and _34605_ (_02990_, _24899_, _23945_);
  and _34606_ (_02991_, _02990_, _24089_);
  not _34607_ (_02992_, _02990_);
  and _34608_ (_02993_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or _34609_ (_27055_, _02993_, _02991_);
  and _34610_ (_02994_, _02970_, _23887_);
  and _34611_ (_02995_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or _34612_ (_23102_, _02995_, _02994_);
  and _34613_ (_02996_, _24301_, _24140_);
  and _34614_ (_02997_, _02996_, _23583_);
  not _34615_ (_02998_, _02996_);
  and _34616_ (_02999_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  or _34617_ (_23110_, _02999_, _02997_);
  and _34618_ (_03001_, _24372_, _24301_);
  and _34619_ (_03002_, _03001_, _23548_);
  not _34620_ (_03003_, _03001_);
  and _34621_ (_03004_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _34622_ (_23135_, _03004_, _03002_);
  and _34623_ (_03005_, _02980_, _23583_);
  and _34624_ (_03006_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _34625_ (_23153_, _03006_, _03005_);
  and _34626_ (_03007_, _02980_, _23887_);
  and _34627_ (_03008_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _34628_ (_23165_, _03008_, _03007_);
  nor _34629_ (_26867_[2], _00223_, rst);
  and _34630_ (_03009_, _24518_, _24219_);
  and _34631_ (_03010_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or _34632_ (_23171_, _03010_, _03009_);
  and _34633_ (_03011_, _02512_, _24372_);
  not _34634_ (_03013_, _03011_);
  and _34635_ (_03014_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and _34636_ (_03015_, _03011_, _24219_);
  or _34637_ (_23180_, _03015_, _03014_);
  nor _34638_ (_26877_[4], _00676_, rst);
  and _34639_ (_03016_, _02990_, _23548_);
  and _34640_ (_03017_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or _34641_ (_23200_, _03017_, _03016_);
  and _34642_ (_03018_, _02980_, _24051_);
  and _34643_ (_03019_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _34644_ (_26971_, _03019_, _03018_);
  and _34645_ (_03020_, _02497_, _24236_);
  and _34646_ (_03021_, _03020_, _23996_);
  not _34647_ (_03022_, _03020_);
  and _34648_ (_03023_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _34649_ (_26952_, _03023_, _03021_);
  and _34650_ (_03024_, _03020_, _24134_);
  and _34651_ (_03025_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _34652_ (_23303_, _03025_, _03024_);
  and _34653_ (_03026_, _24474_, _23945_);
  and _34654_ (_03028_, _03026_, _24051_);
  not _34655_ (_03029_, _03026_);
  and _34656_ (_03030_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _34657_ (_23307_, _03030_, _03028_);
  and _34658_ (_03031_, _24237_, _24051_);
  and _34659_ (_03032_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _34660_ (_23315_, _03032_, _03031_);
  and _34661_ (_03033_, _25413_, _24372_);
  and _34662_ (_03034_, _03033_, _24089_);
  not _34663_ (_03035_, _03033_);
  and _34664_ (_03036_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or _34665_ (_23326_, _03036_, _03034_);
  and _34666_ (_03037_, _03026_, _23996_);
  and _34667_ (_03038_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _34668_ (_23332_, _03038_, _03037_);
  and _34669_ (_03039_, _02980_, _24219_);
  and _34670_ (_03040_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _34671_ (_23339_, _03040_, _03039_);
  and _34672_ (_03041_, _03026_, _24134_);
  and _34673_ (_03042_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _34674_ (_27052_, _03042_, _03041_);
  and _34675_ (_03043_, _24496_, _24236_);
  and _34676_ (_03044_, _03043_, _24051_);
  not _34677_ (_03045_, _03043_);
  and _34678_ (_03046_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or _34679_ (_23365_, _03046_, _03044_);
  nor _34680_ (_26877_[3], _00592_, rst);
  and _34681_ (_03048_, _02497_, _24349_);
  and _34682_ (_03049_, _03048_, _23996_);
  not _34683_ (_03050_, _03048_);
  and _34684_ (_03052_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _34685_ (_26933_, _03052_, _03049_);
  and _34686_ (_03054_, _24442_, _24089_);
  and _34687_ (_03055_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or _34688_ (_23384_, _03055_, _03054_);
  and _34689_ (_03057_, _03048_, _24134_);
  and _34690_ (_03058_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _34691_ (_23389_, _03058_, _03057_);
  and _34692_ (_03059_, _03048_, _24051_);
  and _34693_ (_03060_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _34694_ (_23394_, _03060_, _03059_);
  and _34695_ (_03061_, _03026_, _23583_);
  and _34696_ (_03062_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _34697_ (_23428_, _03062_, _03061_);
  and _34698_ (_03065_, _03020_, _24219_);
  and _34699_ (_03066_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _34700_ (_23431_, _03066_, _03065_);
  and _34701_ (_03067_, _03020_, _23887_);
  and _34702_ (_03068_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _34703_ (_23435_, _03068_, _03067_);
  and _34704_ (_03070_, _02432_, _24134_);
  and _34705_ (_03071_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or _34706_ (_23502_, _03071_, _03070_);
  and _34707_ (_03072_, _24497_, _23887_);
  and _34708_ (_03073_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or _34709_ (_27244_, _03073_, _03072_);
  nor _34710_ (_03074_, _00287_, _26581_);
  nor _34711_ (_03075_, _03074_, _26601_);
  nor _34712_ (_03077_, _00239_, _23893_);
  and _34713_ (_03078_, _03077_, _23902_);
  and _34714_ (_03080_, _03078_, _23931_);
  and _34715_ (_03081_, _03080_, _02374_);
  nor _34716_ (_03082_, _03081_, _24279_);
  nor _34717_ (_03083_, _03082_, _03075_);
  nor _34718_ (_26892_, _03083_, rst);
  and _34719_ (_03084_, _24298_, _24173_);
  and _34720_ (_03085_, _03084_, _25024_);
  and _34721_ (_03086_, _03085_, _22978_);
  nand _34722_ (_03087_, _03086_, _23989_);
  or _34723_ (_03088_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _34724_ (_03089_, _03088_, _22731_);
  and _34725_ (_26854_[7], _03089_, _03087_);
  and _34726_ (_03090_, _03084_, _26779_);
  not _34727_ (_03091_, _03090_);
  nor _34728_ (_03093_, _03091_, _23989_);
  and _34729_ (_03094_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _34730_ (_03096_, _03094_, _22979_);
  or _34731_ (_03097_, _03096_, _03093_);
  or _34732_ (_03098_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _34733_ (_03100_, _03098_, _22731_);
  and _34734_ (_26855_[7], _03100_, _03097_);
  nor _34735_ (_03101_, _03090_, _03085_);
  and _34736_ (_03102_, _03084_, _24627_);
  not _34737_ (_03104_, _03102_);
  and _34738_ (_03105_, _03104_, _03101_);
  nor _34739_ (_03106_, _03105_, _22979_);
  not _34740_ (_03107_, _03106_);
  and _34741_ (_03108_, _03107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _34742_ (_03109_, _03104_, _23989_);
  not _34743_ (_03110_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _34744_ (_03111_, _03101_, _03110_);
  or _34745_ (_03113_, _03111_, _03109_);
  and _34746_ (_03114_, _03113_, _22978_);
  or _34747_ (_03115_, _03114_, _03108_);
  and _34748_ (_26856_[7], _03115_, _22731_);
  and _34749_ (_03118_, _03084_, _24187_);
  and _34750_ (_03119_, _03118_, _22978_);
  and _34751_ (_03120_, _03119_, _25554_);
  nor _34752_ (_03121_, _03118_, _03102_);
  and _34753_ (_03122_, _03121_, _03101_);
  or _34754_ (_03124_, _03122_, _22979_);
  or _34755_ (_03126_, _03124_, _03106_);
  and _34756_ (_03127_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _34757_ (_03128_, _03127_, _03120_);
  and _34758_ (_26857_[7], _03128_, _22731_);
  nand _34759_ (_03129_, _03121_, _03091_);
  and _34760_ (_03131_, _03129_, _22978_);
  and _34761_ (_03132_, _25226_, _24298_);
  and _34762_ (_03133_, _03132_, _25024_);
  not _34763_ (_03134_, _03133_);
  and _34764_ (_03135_, _03134_, _03121_);
  and _34765_ (_03136_, _03135_, _03091_);
  or _34766_ (_03137_, _03085_, _22979_);
  or _34767_ (_03138_, _03137_, _03136_);
  or _34768_ (_03139_, _03138_, _03131_);
  and _34769_ (_03140_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nand _34770_ (_03141_, _03133_, _22978_);
  nor _34771_ (_03142_, _03141_, _23989_);
  or _34772_ (_03143_, _03142_, _03140_);
  and _34773_ (_26858_[7], _03143_, _22731_);
  and _34774_ (_03144_, _03132_, _26779_);
  and _34775_ (_03145_, _03144_, _22978_);
  and _34776_ (_03146_, _03145_, _25554_);
  nor _34777_ (_03147_, _03144_, _03133_);
  and _34778_ (_03148_, _03147_, _03122_);
  or _34779_ (_03149_, _03137_, _03090_);
  nor _34780_ (_03150_, _03149_, _03148_);
  nand _34781_ (_03151_, _03150_, _03135_);
  and _34782_ (_03152_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or _34783_ (_03153_, _03152_, _03146_);
  and _34784_ (_26859_[7], _03153_, _22731_);
  and _34785_ (_03155_, _03132_, _24627_);
  not _34786_ (_03157_, _03155_);
  and _34787_ (_03158_, _03157_, _03148_);
  or _34788_ (_03159_, _03158_, _22979_);
  nor _34789_ (_03161_, _03148_, _22979_);
  or _34790_ (_03162_, _03161_, _03159_);
  and _34791_ (_03164_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand _34792_ (_03165_, _03155_, _22978_);
  nor _34793_ (_03166_, _03165_, _23989_);
  or _34794_ (_03167_, _03166_, _03164_);
  and _34795_ (_26860_[7], _03167_, _22731_);
  and _34796_ (_03168_, _03132_, _24187_);
  and _34797_ (_03169_, _03168_, _25554_);
  and _34798_ (_03170_, _03168_, _22978_);
  not _34799_ (_03171_, _03170_);
  and _34800_ (_03172_, _03171_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or _34801_ (_03173_, _03172_, _03169_);
  or _34802_ (_03174_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _34803_ (_03175_, _03174_, _22731_);
  and _34804_ (_26861_[7], _03175_, _03173_);
  nor _34805_ (_26877_[2], _00496_, rst);
  and _34806_ (_03176_, _03020_, _23548_);
  and _34807_ (_03178_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _34808_ (_26951_, _03178_, _03176_);
  and _34809_ (_03180_, _02497_, _23941_);
  and _34810_ (_03181_, _03180_, _23996_);
  not _34811_ (_03182_, _03180_);
  and _34812_ (_03183_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _34813_ (_23678_, _03183_, _03181_);
  and _34814_ (_03184_, _03048_, _24219_);
  and _34815_ (_03185_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or _34816_ (_23725_, _03185_, _03184_);
  and _34817_ (_03186_, _24056_, _23945_);
  and _34818_ (_03187_, _03186_, _23583_);
  not _34819_ (_03188_, _03186_);
  and _34820_ (_03189_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or _34821_ (_27051_, _03189_, _03187_);
  nor _34822_ (_26877_[1], _00415_, rst);
  and _34823_ (_03190_, _03048_, _23583_);
  and _34824_ (_03191_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _34825_ (_23849_, _03191_, _03190_);
  and _34826_ (_03192_, _24330_, _23996_);
  and _34827_ (_03193_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _34828_ (_23852_, _03193_, _03192_);
  and _34829_ (_03194_, _03048_, _23887_);
  and _34830_ (_03195_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _34831_ (_23866_, _03195_, _03194_);
  nor _34832_ (_26877_[0], _26654_, rst);
  and _34833_ (_03197_, _03180_, _23548_);
  and _34834_ (_03198_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _34835_ (_23942_, _03198_, _03197_);
  and _34836_ (_03199_, _03180_, _24219_);
  and _34837_ (_03200_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _34838_ (_23956_, _03200_, _03199_);
  and _34839_ (_03201_, _03186_, _24219_);
  and _34840_ (_03202_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or _34841_ (_23961_, _03202_, _03201_);
  and _34842_ (_03203_, _03186_, _24134_);
  and _34843_ (_03204_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or _34844_ (_24007_, _03204_, _03203_);
  and _34845_ (_03205_, _03180_, _23583_);
  and _34846_ (_03207_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _34847_ (_24010_, _03207_, _03205_);
  and _34848_ (_03208_, _03180_, _24051_);
  and _34849_ (_03209_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _34850_ (_24012_, _03209_, _03208_);
  and _34851_ (_03210_, _03180_, _24089_);
  and _34852_ (_03211_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _34853_ (_24046_, _03211_, _03210_);
  and _34854_ (_03212_, _03186_, _24051_);
  and _34855_ (_03213_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or _34856_ (_24049_, _03213_, _03212_);
  and _34857_ (_03214_, _03186_, _23996_);
  and _34858_ (_03215_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or _34859_ (_24084_, _03215_, _03214_);
  and _34860_ (_03217_, _02497_, _24899_);
  and _34861_ (_03218_, _03217_, _23887_);
  not _34862_ (_03219_, _03217_);
  and _34863_ (_03220_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _34864_ (_24090_, _03220_, _03218_);
  and _34865_ (_03221_, _02512_, _24319_);
  not _34866_ (_03222_, _03221_);
  and _34867_ (_03224_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  and _34868_ (_03225_, _03221_, _23583_);
  or _34869_ (_24103_, _03225_, _03224_);
  and _34870_ (_03226_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  and _34871_ (_03227_, _03221_, _23887_);
  or _34872_ (_24128_, _03227_, _03226_);
  and _34873_ (_03228_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and _34874_ (_03229_, _03221_, _23548_);
  or _34875_ (_24135_, _03229_, _03228_);
  and _34876_ (_03230_, _03217_, _24134_);
  and _34877_ (_03231_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _34878_ (_24138_, _03231_, _03230_);
  and _34879_ (_03232_, _03217_, _24051_);
  and _34880_ (_03233_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _34881_ (_24168_, _03233_, _03232_);
  and _34882_ (_03234_, _03217_, _24089_);
  and _34883_ (_03235_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _34884_ (_27312_, _03235_, _03234_);
  and _34885_ (_03236_, _24408_, _24095_);
  and _34886_ (_03237_, _03236_, _23996_);
  not _34887_ (_03238_, _03236_);
  and _34888_ (_03239_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _34889_ (_24183_, _03239_, _03237_);
  and _34890_ (_03241_, _25413_, _23941_);
  and _34891_ (_03242_, _03241_, _24051_);
  not _34892_ (_03243_, _03241_);
  and _34893_ (_03244_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  or _34894_ (_24191_, _03244_, _03242_);
  and _34895_ (_03245_, _25413_, _24899_);
  and _34896_ (_03246_, _03245_, _23996_);
  not _34897_ (_03247_, _03245_);
  and _34898_ (_03248_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or _34899_ (_24195_, _03248_, _03246_);
  and _34900_ (_03249_, _03245_, _23548_);
  and _34901_ (_03250_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  or _34902_ (_24199_, _03250_, _03249_);
  and _34903_ (_03251_, _02497_, _24474_);
  and _34904_ (_03252_, _03251_, _24089_);
  not _34905_ (_03253_, _03251_);
  and _34906_ (_03254_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _34907_ (_24202_, _03254_, _03252_);
  and _34908_ (_03255_, _25413_, _24474_);
  and _34909_ (_03256_, _03255_, _23583_);
  not _34910_ (_03257_, _03255_);
  and _34911_ (_03258_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _34912_ (_24205_, _03258_, _03256_);
  and _34913_ (_03259_, _03251_, _23583_);
  and _34914_ (_03260_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _34915_ (_24211_, _03260_, _03259_);
  and _34916_ (_03261_, _03236_, _24089_);
  and _34917_ (_03263_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _34918_ (_24213_, _03263_, _03261_);
  and _34919_ (_03264_, _03236_, _24134_);
  and _34920_ (_03265_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _34921_ (_24215_, _03265_, _03264_);
  and _34922_ (_03266_, _03251_, _23887_);
  and _34923_ (_03267_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _34924_ (_27290_, _03267_, _03266_);
  and _34925_ (_03269_, _25413_, _24056_);
  and _34926_ (_03270_, _03269_, _24219_);
  not _34927_ (_03271_, _03269_);
  and _34928_ (_03272_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or _34929_ (_24222_, _03272_, _03270_);
  and _34930_ (_03273_, _03251_, _23548_);
  and _34931_ (_03274_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _34932_ (_27289_, _03274_, _03273_);
  and _34933_ (_03275_, _25413_, _24223_);
  and _34934_ (_03276_, _03275_, _24089_);
  not _34935_ (_03277_, _03275_);
  and _34936_ (_03278_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _34937_ (_24227_, _03278_, _03276_);
  and _34938_ (_03279_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  and _34939_ (_03280_, _02513_, _23996_);
  or _34940_ (_24235_, _03280_, _03279_);
  and _34941_ (_03281_, _25413_, _24319_);
  and _34942_ (_03282_, _03281_, _24219_);
  not _34943_ (_03283_, _03281_);
  and _34944_ (_03284_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or _34945_ (_24241_, _03284_, _03282_);
  and _34946_ (_03285_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  and _34947_ (_03286_, _03221_, _24134_);
  or _34948_ (_24242_, _03286_, _03285_);
  and _34949_ (_03287_, _25413_, _24095_);
  and _34950_ (_03288_, _03287_, _24134_);
  not _34951_ (_03289_, _03287_);
  and _34952_ (_03290_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or _34953_ (_24252_, _03290_, _03288_);
  and _34954_ (_03291_, _03251_, _23996_);
  and _34955_ (_03292_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _34956_ (_24256_, _03292_, _03291_);
  and _34957_ (_03293_, _03287_, _23887_);
  and _34958_ (_03294_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or _34959_ (_24280_, _03294_, _03293_);
  and _34960_ (_03295_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  and _34961_ (_03296_, _03221_, _24051_);
  or _34962_ (_24282_, _03296_, _03295_);
  and _34963_ (_03298_, _03251_, _24134_);
  and _34964_ (_03299_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or _34965_ (_24285_, _03299_, _03298_);
  and _34966_ (_03301_, _03251_, _24051_);
  and _34967_ (_03302_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _34968_ (_24288_, _03302_, _03301_);
  and _34969_ (_03303_, _03033_, _24051_);
  and _34970_ (_03304_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or _34971_ (_27162_, _03304_, _03303_);
  and _34972_ (_03305_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  and _34973_ (_03306_, _03221_, _24089_);
  or _34974_ (_24316_, _03306_, _03305_);
  and _34975_ (_03307_, _23944_, _22847_);
  and _34976_ (_03308_, _24003_, _03307_);
  and _34977_ (_03309_, _03308_, _24223_);
  and _34978_ (_03310_, _03309_, _24219_);
  not _34979_ (_03311_, _03309_);
  and _34980_ (_03312_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or _34981_ (_26962_, _03312_, _03310_);
  and _34982_ (_03313_, _25413_, _24297_);
  and _34983_ (_03314_, _03313_, _23583_);
  not _34984_ (_03315_, _03313_);
  and _34985_ (_03316_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or _34986_ (_27177_, _03316_, _03314_);
  and _34987_ (_03317_, _03313_, _24219_);
  and _34988_ (_03318_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or _34989_ (_24326_, _03318_, _03317_);
  and _34990_ (_03319_, _02512_, _22974_);
  not _34991_ (_03320_, _03319_);
  and _34992_ (_03322_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _34993_ (_03323_, _03319_, _23583_);
  or _34994_ (_24329_, _03323_, _03322_);
  and _34995_ (_03324_, _02497_, _24056_);
  and _34996_ (_03325_, _03324_, _24134_);
  not _34997_ (_03326_, _03324_);
  and _34998_ (_03327_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _34999_ (_24335_, _03327_, _03325_);
  and _35000_ (_03328_, _03324_, _24051_);
  and _35001_ (_03329_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _35002_ (_24338_, _03329_, _03328_);
  and _35003_ (_03330_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _35004_ (_03331_, _03319_, _24089_);
  or _35005_ (_24344_, _03331_, _03330_);
  and _35006_ (_03332_, _24518_, _23887_);
  and _35007_ (_03333_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or _35008_ (_24346_, _03333_, _03332_);
  and _35009_ (_03334_, _03324_, _23996_);
  and _35010_ (_03335_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _35011_ (_24356_, _03335_, _03334_);
  and _35012_ (_03337_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _35013_ (_03338_, _03319_, _24134_);
  or _35014_ (_24359_, _03338_, _03337_);
  and _35015_ (_03340_, _02488_, _24219_);
  and _35016_ (_03341_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or _35017_ (_24363_, _03341_, _03340_);
  and _35018_ (_03343_, _02497_, _24223_);
  and _35019_ (_03344_, _03343_, _23996_);
  not _35020_ (_03346_, _03343_);
  and _35021_ (_03347_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _35022_ (_24366_, _03347_, _03344_);
  and _35023_ (_03348_, _03324_, _24219_);
  and _35024_ (_03349_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _35025_ (_27258_, _03349_, _03348_);
  and _35026_ (_03350_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and _35027_ (_03351_, _03319_, _23996_);
  or _35028_ (_24370_, _03351_, _03350_);
  and _35029_ (_03353_, _02767_, _24089_);
  and _35030_ (_03354_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or _35031_ (_24390_, _03354_, _03353_);
  and _35032_ (_03355_, _24159_, _24141_);
  and _35033_ (_03356_, _03355_, _23548_);
  not _35034_ (_03357_, _03355_);
  and _35035_ (_03358_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _35036_ (_24419_, _03358_, _03356_);
  and _35037_ (_03360_, _25413_, _24236_);
  and _35038_ (_03361_, _03360_, _24134_);
  not _35039_ (_03362_, _03360_);
  and _35040_ (_03363_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or _35041_ (_24423_, _03363_, _03361_);
  and _35042_ (_03364_, _03313_, _23996_);
  and _35043_ (_03365_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or _35044_ (_24429_, _03365_, _03364_);
  and _35045_ (_03366_, _03360_, _24089_);
  and _35046_ (_03367_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _35047_ (_24432_, _03367_, _03366_);
  and _35048_ (_03368_, _03324_, _23887_);
  and _35049_ (_03369_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _35050_ (_24435_, _03369_, _03368_);
  and _35051_ (_26840_[2], _23639_, _22731_);
  and _35052_ (_03370_, _24408_, _22974_);
  and _35053_ (_03371_, _03370_, _24219_);
  not _35054_ (_03372_, _03370_);
  and _35055_ (_03373_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _35056_ (_27117_, _03373_, _03371_);
  and _35057_ (_03374_, _03370_, _23887_);
  and _35058_ (_03375_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _35059_ (_24445_, _03375_, _03374_);
  and _35060_ (_03376_, _03343_, _23887_);
  and _35061_ (_03377_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _35062_ (_27243_, _03377_, _03376_);
  and _35063_ (_03378_, _03343_, _23548_);
  and _35064_ (_03379_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _35065_ (_24456_, _03379_, _03378_);
  and _35066_ (_03380_, _03343_, _24219_);
  and _35067_ (_03381_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _35068_ (_24463_, _03381_, _03380_);
  and _35069_ (_03382_, _03287_, _23996_);
  and _35070_ (_03383_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or _35071_ (_24466_, _03383_, _03382_);
  and _35072_ (_03384_, _03355_, _24089_);
  and _35073_ (_03385_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _35074_ (_24475_, _03385_, _03384_);
  and _35075_ (_03386_, _03370_, _24051_);
  and _35076_ (_03387_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _35077_ (_24477_, _03387_, _03386_);
  and _35078_ (_03388_, _02432_, _23548_);
  and _35079_ (_03390_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  or _35080_ (_24483_, _03390_, _03388_);
  and _35081_ (_03391_, _03370_, _24134_);
  and _35082_ (_03392_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _35083_ (_24488_, _03392_, _03391_);
  and _35084_ (_03393_, _02767_, _24051_);
  and _35085_ (_03394_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _35086_ (_24498_, _03394_, _03393_);
  and _35087_ (_03396_, _03343_, _24051_);
  and _35088_ (_03397_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _35089_ (_24501_, _03397_, _03396_);
  and _35090_ (_03398_, _03343_, _24089_);
  and _35091_ (_03400_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _35092_ (_24506_, _03400_, _03398_);
  and _35093_ (_03402_, _03343_, _23583_);
  and _35094_ (_03403_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _35095_ (_24524_, _03403_, _03402_);
  not _35096_ (_03404_, _03086_);
  and _35097_ (_03405_, _03404_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _35098_ (_03406_, _03086_, _24671_);
  or _35099_ (_03407_, _03406_, _03405_);
  and _35100_ (_26854_[0], _03407_, _22731_);
  nand _35101_ (_03408_, _03086_, _23542_);
  or _35102_ (_03409_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _35103_ (_03410_, _03409_, _22731_);
  and _35104_ (_26854_[1], _03410_, _03408_);
  or _35105_ (_03411_, _03404_, _23880_);
  or _35106_ (_03412_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _35107_ (_03413_, _03412_, _22731_);
  and _35108_ (_26854_[2], _03413_, _03411_);
  or _35109_ (_03414_, _03404_, _23577_);
  or _35110_ (_03416_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _35111_ (_03417_, _03416_, _22731_);
  and _35112_ (_26854_[3], _03417_, _03414_);
  nand _35113_ (_03419_, _03086_, _24082_);
  or _35114_ (_03420_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _35115_ (_03421_, _03420_, _22731_);
  and _35116_ (_26854_[4], _03421_, _03419_);
  nand _35117_ (_03423_, _03086_, _24043_);
  or _35118_ (_03424_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _35119_ (_03425_, _03424_, _22731_);
  and _35120_ (_26854_[5], _03425_, _03423_);
  nand _35121_ (_03428_, _03086_, _24126_);
  or _35122_ (_03429_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _35123_ (_03430_, _03429_, _22731_);
  and _35124_ (_26854_[6], _03430_, _03428_);
  and _35125_ (_03431_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _35126_ (_03432_, _03090_, _24671_);
  or _35127_ (_03433_, _03432_, _22979_);
  or _35128_ (_03434_, _03433_, _03431_);
  or _35129_ (_03435_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _35130_ (_03436_, _03435_, _22731_);
  and _35131_ (_26855_[0], _03436_, _03434_);
  nor _35132_ (_03437_, _03091_, _23542_);
  and _35133_ (_03438_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _35134_ (_03439_, _03438_, _22979_);
  or _35135_ (_03441_, _03439_, _03437_);
  or _35136_ (_03442_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _35137_ (_03444_, _03442_, _22731_);
  and _35138_ (_26855_[1], _03444_, _03441_);
  and _35139_ (_03445_, _03090_, _23880_);
  and _35140_ (_03446_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _35141_ (_03447_, _03446_, _22979_);
  or _35142_ (_03448_, _03447_, _03445_);
  or _35143_ (_03449_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _35144_ (_03450_, _03449_, _22731_);
  and _35145_ (_26855_[2], _03450_, _03448_);
  and _35146_ (_03451_, _03090_, _23577_);
  and _35147_ (_03452_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _35148_ (_03453_, _03452_, _22979_);
  or _35149_ (_03454_, _03453_, _03451_);
  or _35150_ (_03455_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _35151_ (_03457_, _03455_, _22731_);
  and _35152_ (_26855_[3], _03457_, _03454_);
  nor _35153_ (_03458_, _03091_, _24082_);
  and _35154_ (_03459_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _35155_ (_03460_, _03459_, _22979_);
  or _35156_ (_03461_, _03460_, _03458_);
  or _35157_ (_03462_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _35158_ (_03463_, _03462_, _22731_);
  and _35159_ (_26855_[4], _03463_, _03461_);
  nor _35160_ (_03464_, _03091_, _24043_);
  and _35161_ (_03465_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _35162_ (_03466_, _03465_, _22979_);
  or _35163_ (_03468_, _03466_, _03464_);
  or _35164_ (_03469_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _35165_ (_03470_, _03469_, _22731_);
  and _35166_ (_26855_[5], _03470_, _03468_);
  nor _35167_ (_03471_, _03091_, _24126_);
  and _35168_ (_03473_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _35169_ (_03474_, _03473_, _22979_);
  or _35170_ (_03476_, _03474_, _03471_);
  or _35171_ (_03478_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _35172_ (_03479_, _03478_, _22731_);
  and _35173_ (_26855_[6], _03479_, _03476_);
  and _35174_ (_03481_, _03107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand _35175_ (_03482_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _35176_ (_03484_, _03482_, _03101_);
  nor _35177_ (_03485_, _24210_, _22979_);
  and _35178_ (_03487_, _03485_, _03102_);
  or _35179_ (_03488_, _03487_, _03484_);
  or _35180_ (_03489_, _03488_, _03481_);
  and _35181_ (_26856_[0], _03489_, _22731_);
  or _35182_ (_03490_, _03101_, _22979_);
  nand _35183_ (_03491_, _03490_, _03106_);
  and _35184_ (_03492_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nand _35185_ (_03493_, _03102_, _22978_);
  nor _35186_ (_03494_, _03493_, _23542_);
  or _35187_ (_03495_, _03494_, _03492_);
  and _35188_ (_26856_[1], _03495_, _22731_);
  and _35189_ (_03496_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _35190_ (_03497_, _23880_, _22978_);
  and _35191_ (_03499_, _03497_, _03102_);
  or _35192_ (_03500_, _03499_, _03496_);
  and _35193_ (_26856_[2], _03500_, _22731_);
  and _35194_ (_03501_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _35195_ (_03502_, _23577_, _22978_);
  and _35196_ (_03503_, _03502_, _03102_);
  or _35197_ (_03504_, _03503_, _03501_);
  and _35198_ (_26856_[3], _03504_, _22731_);
  and _35199_ (_03505_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _35200_ (_03506_, _24082_, _22979_);
  and _35201_ (_03508_, _03506_, _03102_);
  or _35202_ (_03510_, _03508_, _03505_);
  and _35203_ (_26856_[4], _03510_, _22731_);
  and _35204_ (_03512_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _35205_ (_03513_, _24043_, _22979_);
  and _35206_ (_03514_, _03513_, _03102_);
  or _35207_ (_03515_, _03514_, _03512_);
  and _35208_ (_26856_[5], _03515_, _22731_);
  and _35209_ (_03516_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _35210_ (_03517_, _24126_, _22979_);
  and _35211_ (_03518_, _03517_, _03102_);
  or _35212_ (_03520_, _03518_, _03516_);
  and _35213_ (_26856_[6], _03520_, _22731_);
  and _35214_ (_03521_, _03119_, _24671_);
  and _35215_ (_03522_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _35216_ (_03523_, _03522_, _03521_);
  and _35217_ (_26857_[0], _03523_, _22731_);
  and _35218_ (_03524_, _03119_, _02728_);
  and _35219_ (_03525_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _35220_ (_03526_, _03525_, _03524_);
  and _35221_ (_26857_[1], _03526_, _22731_);
  and _35222_ (_03527_, _03119_, _23880_);
  and _35223_ (_03528_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or _35224_ (_03530_, _03528_, _03527_);
  and _35225_ (_26857_[2], _03530_, _22731_);
  and _35226_ (_03531_, _03119_, _23577_);
  and _35227_ (_03532_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _35228_ (_03534_, _03532_, _03531_);
  and _35229_ (_26857_[3], _03534_, _22731_);
  and _35230_ (_03535_, _03119_, _02700_);
  and _35231_ (_03536_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or _35232_ (_03537_, _03536_, _03535_);
  and _35233_ (_26857_[4], _03537_, _22731_);
  and _35234_ (_03538_, _03119_, _02689_);
  and _35235_ (_03540_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _35236_ (_03541_, _03540_, _03538_);
  and _35237_ (_26857_[5], _03541_, _22731_);
  and _35238_ (_03542_, _03119_, _02450_);
  and _35239_ (_03543_, _03124_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nand _35240_ (_03544_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _35241_ (_03545_, _03544_, _03105_);
  or _35242_ (_03546_, _03545_, _03543_);
  or _35243_ (_03547_, _03546_, _03542_);
  and _35244_ (_26857_[6], _03547_, _22731_);
  and _35245_ (_03549_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _35246_ (_03550_, _03485_, _03133_);
  or _35247_ (_03551_, _03550_, _03549_);
  and _35248_ (_26858_[0], _03551_, _22731_);
  and _35249_ (_03552_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _35250_ (_03554_, _23542_, _22979_);
  and _35251_ (_03555_, _03554_, _03133_);
  or _35252_ (_03556_, _03555_, _03552_);
  and _35253_ (_26858_[1], _03556_, _22731_);
  and _35254_ (_03557_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _35255_ (_03558_, _03497_, _03133_);
  or _35256_ (_03559_, _03558_, _03557_);
  and _35257_ (_26858_[2], _03559_, _22731_);
  and _35258_ (_03561_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _35259_ (_03562_, _03502_, _03133_);
  or _35260_ (_03563_, _03562_, _03561_);
  and _35261_ (_26858_[3], _03563_, _22731_);
  and _35262_ (_03564_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _35263_ (_03565_, _03506_, _03133_);
  or _35264_ (_03566_, _03565_, _03564_);
  and _35265_ (_26858_[4], _03566_, _22731_);
  and _35266_ (_03567_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _35267_ (_03568_, _03513_, _03133_);
  or _35268_ (_03569_, _03568_, _03567_);
  and _35269_ (_26858_[5], _03569_, _22731_);
  and _35270_ (_03570_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _35271_ (_03571_, _03517_, _03133_);
  or _35272_ (_03572_, _03571_, _03570_);
  and _35273_ (_26858_[6], _03572_, _22731_);
  and _35274_ (_03574_, _03485_, _03144_);
  and _35275_ (_03575_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  or _35276_ (_03577_, _03575_, _03574_);
  and _35277_ (_26859_[0], _03577_, _22731_);
  and _35278_ (_03578_, _03145_, _02728_);
  and _35279_ (_03579_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  or _35280_ (_03580_, _03579_, _03578_);
  and _35281_ (_26859_[1], _03580_, _22731_);
  and _35282_ (_03581_, _03145_, _23880_);
  and _35283_ (_03582_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or _35284_ (_03583_, _03582_, _03581_);
  and _35285_ (_26859_[2], _03583_, _22731_);
  and _35286_ (_03585_, _03145_, _23577_);
  and _35287_ (_03586_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or _35288_ (_03587_, _03586_, _03585_);
  and _35289_ (_26859_[3], _03587_, _22731_);
  and _35290_ (_03588_, _03145_, _02700_);
  and _35291_ (_03589_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or _35292_ (_03590_, _03589_, _03588_);
  and _35293_ (_26859_[4], _03590_, _22731_);
  and _35294_ (_03591_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _35295_ (_03592_, _03145_, _02689_);
  or _35296_ (_03593_, _03592_, _03591_);
  and _35297_ (_26859_[5], _03593_, _22731_);
  and _35298_ (_03594_, _03145_, _02450_);
  and _35299_ (_03595_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _35300_ (_03596_, _03595_, _03594_);
  and _35301_ (_26859_[6], _03596_, _22731_);
  and _35302_ (_03597_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _35303_ (_03599_, _03485_, _03155_);
  or _35304_ (_03600_, _03599_, _03597_);
  and _35305_ (_26860_[0], _03600_, _22731_);
  and _35306_ (_03601_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _35307_ (_03602_, _03554_, _03155_);
  or _35308_ (_03603_, _03602_, _03601_);
  and _35309_ (_26860_[1], _03603_, _22731_);
  and _35310_ (_03604_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _35311_ (_03606_, _03497_, _03155_);
  or _35312_ (_03607_, _03606_, _03604_);
  and _35313_ (_26860_[2], _03607_, _22731_);
  and _35314_ (_03608_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _35315_ (_03610_, _03502_, _03155_);
  or _35316_ (_03611_, _03610_, _03608_);
  and _35317_ (_26860_[3], _03611_, _22731_);
  and _35318_ (_03612_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _35319_ (_03613_, _03506_, _03155_);
  or _35320_ (_03614_, _03613_, _03612_);
  and _35321_ (_26860_[4], _03614_, _22731_);
  nor _35322_ (_03615_, _03157_, _24043_);
  and _35323_ (_03616_, _03157_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _35324_ (_03617_, _03616_, _22979_);
  or _35325_ (_03618_, _03617_, _03615_);
  or _35326_ (_03619_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _35327_ (_03620_, _03619_, _22731_);
  and _35328_ (_26860_[5], _03620_, _03618_);
  and _35329_ (_03621_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _35330_ (_03622_, _03517_, _03155_);
  or _35331_ (_03623_, _03622_, _03621_);
  and _35332_ (_26860_[6], _03623_, _22731_);
  nand _35333_ (_03624_, _03157_, _03147_);
  nor _35334_ (_03625_, _03168_, _03624_);
  or _35335_ (_03626_, _03625_, _22979_);
  and _35336_ (_03628_, _03626_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _35337_ (_03629_, _03485_, _03168_);
  and _35338_ (_03630_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _35339_ (_03632_, _03630_, _03624_);
  or _35340_ (_03633_, _03632_, _03629_);
  or _35341_ (_03634_, _03633_, _03628_);
  and _35342_ (_26861_[0], _03634_, _22731_);
  and _35343_ (_03635_, _03626_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _35344_ (_03636_, _03171_, _23542_);
  and _35345_ (_03637_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _35346_ (_03638_, _03637_, _03624_);
  or _35347_ (_03639_, _03638_, _03636_);
  or _35348_ (_03640_, _03639_, _03635_);
  and _35349_ (_26861_[1], _03640_, _22731_);
  and _35350_ (_03641_, _03170_, _23880_);
  or _35351_ (_03642_, _03137_, _03129_);
  or _35352_ (_03643_, _03642_, _03625_);
  and _35353_ (_03644_, _03624_, _22978_);
  or _35354_ (_03645_, _03644_, _03643_);
  and _35355_ (_03646_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _35356_ (_03647_, _03646_, _03641_);
  and _35357_ (_26861_[2], _03647_, _22731_);
  and _35358_ (_03649_, _03170_, _23577_);
  and _35359_ (_03650_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or _35360_ (_03651_, _03650_, _03649_);
  and _35361_ (_26861_[3], _03651_, _22731_);
  nor _35362_ (_03652_, _03171_, _24082_);
  and _35363_ (_03653_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _35364_ (_03654_, _03653_, _03652_);
  and _35365_ (_26861_[4], _03654_, _22731_);
  and _35366_ (_03655_, _03171_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _35367_ (_03656_, _03171_, _24043_);
  or _35368_ (_03657_, _03656_, _03655_);
  and _35369_ (_26861_[5], _03657_, _22731_);
  nor _35370_ (_03658_, _03171_, _24126_);
  and _35371_ (_03660_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or _35372_ (_03661_, _03660_, _03658_);
  and _35373_ (_26861_[6], _03661_, _22731_);
  and _35374_ (_03662_, _02512_, _24056_);
  not _35375_ (_03663_, _03662_);
  and _35376_ (_03665_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _35377_ (_03666_, _03662_, _23583_);
  or _35378_ (_24958_, _03666_, _03665_);
  and _35379_ (_03667_, _02497_, _24319_);
  and _35380_ (_03668_, _03667_, _24089_);
  not _35381_ (_03669_, _03667_);
  and _35382_ (_03670_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or _35383_ (_25031_, _03670_, _03668_);
  and _35384_ (_03672_, _02970_, _24051_);
  and _35385_ (_03674_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or _35386_ (_25037_, _03674_, _03672_);
  and _35387_ (_03676_, _02502_, _24051_);
  and _35388_ (_03677_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or _35389_ (_25076_, _03677_, _03676_);
  and _35390_ (_03678_, _02890_, _24219_);
  and _35391_ (_03679_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or _35392_ (_25079_, _03679_, _03678_);
  and _35393_ (_03680_, _02502_, _24134_);
  and _35394_ (_03681_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _35395_ (_25082_, _03681_, _03680_);
  and _35396_ (_03682_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and _35397_ (_03683_, _03662_, _23887_);
  or _35398_ (_25087_, _03683_, _03682_);
  and _35399_ (_03684_, _02970_, _23996_);
  and _35400_ (_03685_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or _35401_ (_27229_, _03685_, _03684_);
  and _35402_ (_03686_, _02970_, _24134_);
  and _35403_ (_03687_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or _35404_ (_25170_, _03687_, _03686_);
  not _35405_ (_03688_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _35406_ (_03689_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and _35407_ (_03690_, _03689_, _03688_);
  and _35408_ (_03691_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _22731_);
  and _35409_ (_27314_, _03691_, _03690_);
  nor _35410_ (_03692_, _03690_, rst);
  nand _35411_ (_03693_, _03689_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _35412_ (_03694_, _03689_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _35413_ (_03696_, _03694_, _03693_);
  and _35414_ (_27315_[3], _03696_, _03692_);
  not _35415_ (_03698_, _00051_);
  nor _35416_ (_03699_, _03698_, _00090_);
  not _35417_ (_03700_, _00027_);
  and _35418_ (_03702_, _03700_, _00143_);
  and _35419_ (_03703_, _03702_, _26816_);
  and _35420_ (_03705_, _03703_, _03699_);
  not _35421_ (_03706_, _00325_);
  nand _35422_ (_03707_, _00569_, _03706_);
  nor _35423_ (_03708_, _24533_, _23195_);
  nor _35424_ (_03709_, _03708_, _24534_);
  and _35425_ (_03710_, _00329_, _00326_);
  not _35426_ (_03711_, _03710_);
  nor _35427_ (_03712_, _03711_, _03709_);
  and _35428_ (_03713_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _35429_ (_03714_, _03713_, _00319_);
  nor _35430_ (_03715_, _03714_, _03712_);
  nand _35431_ (_03717_, _03715_, _03707_);
  and _35432_ (_03719_, _01121_, _00319_);
  not _35433_ (_03720_, _03719_);
  nand _35434_ (_03721_, _03720_, _03717_);
  nand _35435_ (_03722_, _00473_, _03706_);
  nor _35436_ (_03723_, _24562_, _23210_);
  nor _35437_ (_03724_, _03723_, _02580_);
  nor _35438_ (_03725_, _03724_, _03711_);
  and _35439_ (_03727_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _35440_ (_03728_, _03727_, _03725_);
  and _35441_ (_03729_, _03728_, _00320_);
  and _35442_ (_03730_, _03729_, _03722_);
  and _35443_ (_03731_, _01061_, _00319_);
  nor _35444_ (_03732_, _03731_, _03730_);
  nand _35445_ (_03733_, _03732_, _03721_);
  or _35446_ (_03734_, _03732_, _03721_);
  nand _35447_ (_03735_, _03734_, _03733_);
  nand _35448_ (_03736_, _26570_, _03706_);
  nor _35449_ (_03737_, _24577_, _23291_);
  nor _35450_ (_03738_, _03737_, _02599_);
  nor _35451_ (_03739_, _03738_, _03711_);
  and _35452_ (_03740_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _35453_ (_03742_, _03740_, _00319_);
  nor _35454_ (_03743_, _03742_, _03739_);
  nand _35455_ (_03744_, _03743_, _03736_);
  or _35456_ (_03745_, _00939_, _00320_);
  and _35457_ (_03746_, _03745_, _03744_);
  nand _35458_ (_03747_, _00393_, _03706_);
  nor _35459_ (_03748_, _24177_, _23260_);
  nor _35460_ (_03750_, _03748_, _02590_);
  nor _35461_ (_03751_, _03750_, _03711_);
  and _35462_ (_03752_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _35463_ (_03754_, _03752_, _00319_);
  nor _35464_ (_03755_, _03754_, _03751_);
  nand _35465_ (_03756_, _03755_, _03747_);
  and _35466_ (_03757_, _01009_, _00319_);
  not _35467_ (_03758_, _03757_);
  nand _35468_ (_03759_, _03758_, _03756_);
  nand _35469_ (_03760_, _03759_, _03746_);
  or _35470_ (_03762_, _03759_, _03746_);
  nand _35471_ (_03763_, _03762_, _03760_);
  nand _35472_ (_03764_, _03763_, _03735_);
  or _35473_ (_03765_, _03763_, _03735_);
  nand _35474_ (_03767_, _03765_, _03764_);
  nand _35475_ (_03769_, _00654_, _03706_);
  nor _35476_ (_03770_, _24636_, _23145_);
  nor _35477_ (_03771_, _03770_, _24637_);
  nor _35478_ (_03772_, _03771_, _03711_);
  and _35479_ (_03773_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _35480_ (_03774_, _03773_, _00319_);
  nor _35481_ (_03775_, _03774_, _03772_);
  nand _35482_ (_03776_, _03775_, _03769_);
  and _35483_ (_03777_, _01192_, _00319_);
  not _35484_ (_03778_, _03777_);
  and _35485_ (_03779_, _03778_, _03776_);
  nand _35486_ (_03781_, _00747_, _03706_);
  nand _35487_ (_03782_, _24607_, _23504_);
  or _35488_ (_03783_, _24607_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _35489_ (_03784_, _03783_, _03710_);
  and _35490_ (_03785_, _03784_, _03782_);
  and _35491_ (_03786_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _35492_ (_03787_, _03786_, _00319_);
  nor _35493_ (_03788_, _03787_, _03785_);
  nand _35494_ (_03789_, _03788_, _03781_);
  and _35495_ (_03790_, _01281_, _00319_);
  not _35496_ (_03791_, _03790_);
  and _35497_ (_03792_, _03791_, _03789_);
  or _35498_ (_03793_, _03792_, _03779_);
  nand _35499_ (_03794_, _03792_, _03779_);
  nand _35500_ (_03795_, _03794_, _03793_);
  or _35501_ (_03796_, _00813_, _00325_);
  not _35502_ (_03797_, _24594_);
  nor _35503_ (_03798_, _03797_, _23504_);
  nor _35504_ (_03799_, _24594_, _23074_);
  nor _35505_ (_03801_, _03799_, _03798_);
  nor _35506_ (_03802_, _03801_, _03711_);
  and _35507_ (_03803_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _35508_ (_03805_, _03803_, _00319_);
  nor _35509_ (_03806_, _03805_, _03802_);
  and _35510_ (_03807_, _03806_, _03796_);
  and _35511_ (_03808_, _01353_, _00319_);
  or _35512_ (_03809_, _03808_, _03807_);
  and _35513_ (_03810_, _00883_, _03706_);
  nor _35514_ (_03811_, _25481_, _23034_);
  or _35515_ (_03813_, _03811_, _25482_);
  and _35516_ (_03814_, _03813_, _03710_);
  and _35517_ (_03815_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _35518_ (_03816_, _03815_, _00319_);
  or _35519_ (_03818_, _03816_, _03814_);
  or _35520_ (_03819_, _03818_, _03810_);
  nor _35521_ (_03821_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _35522_ (_03822_, _23003_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _35523_ (_03823_, _03822_, _03821_);
  nor _35524_ (_03824_, _03823_, _01319_);
  and _35525_ (_03825_, _03823_, _01319_);
  or _35526_ (_03826_, _03825_, _03824_);
  and _35527_ (_03828_, _03826_, _23390_);
  or _35528_ (_03829_, _26539_, _26501_);
  and _35529_ (_03830_, _03829_, _26540_);
  and _35530_ (_03831_, _03830_, _23531_);
  and _35531_ (_03832_, _01259_, _23120_);
  and _35532_ (_03833_, _03832_, _23086_);
  nor _35533_ (_03834_, _03833_, _01329_);
  or _35534_ (_03835_, _03834_, _01341_);
  or _35535_ (_03837_, _03835_, _23049_);
  nand _35536_ (_03838_, _03835_, _23049_);
  and _35537_ (_03839_, _03838_, _23514_);
  and _35538_ (_03840_, _03839_, _03837_);
  and _35539_ (_03841_, _23364_, _23050_);
  or _35540_ (_03842_, _03841_, _23472_);
  and _35541_ (_03843_, _03842_, _23506_);
  and _35542_ (_03844_, _23488_, _23563_);
  and _35543_ (_03845_, _23484_, _23050_);
  and _35544_ (_03846_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or _35545_ (_03847_, _03846_, _03845_);
  or _35546_ (_03849_, _03847_, _03844_);
  or _35547_ (_03850_, _03849_, _03843_);
  or _35548_ (_03851_, _03850_, _03840_);
  or _35549_ (_03852_, _03851_, _03831_);
  or _35550_ (_03853_, _03852_, _03828_);
  or _35551_ (_03855_, _03853_, _00320_);
  and _35552_ (_03857_, _03855_, _03819_);
  or _35553_ (_03858_, _03857_, _03809_);
  nand _35554_ (_03859_, _03857_, _03809_);
  and _35555_ (_03860_, _03859_, _03858_);
  nand _35556_ (_03861_, _03860_, _03795_);
  or _35557_ (_03862_, _03860_, _03795_);
  nand _35558_ (_03863_, _03862_, _03861_);
  nand _35559_ (_03865_, _03863_, _03767_);
  or _35560_ (_03866_, _03863_, _03767_);
  nand _35561_ (_03868_, _03866_, _03865_);
  nand _35562_ (_03869_, _03868_, _00228_);
  and _35563_ (_03870_, _00191_, _00171_);
  or _35564_ (_03871_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _35565_ (_03872_, _03871_, _03870_);
  and _35566_ (_03873_, _03872_, _03869_);
  not _35567_ (_03874_, _00228_);
  not _35568_ (_03875_, _00191_);
  and _35569_ (_03876_, _03875_, _00171_);
  and _35570_ (_03877_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor _35571_ (_03878_, _00191_, _00171_);
  and _35572_ (_03879_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _35573_ (_03880_, _03879_, _03877_);
  and _35574_ (_03881_, _03880_, _03874_);
  not _35575_ (_03882_, _00171_);
  and _35576_ (_03883_, _00191_, _03882_);
  nor _35577_ (_03884_, _00228_, _00546_);
  and _35578_ (_03885_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _35579_ (_03886_, _03885_, _03884_);
  and _35580_ (_03887_, _03886_, _03883_);
  and _35581_ (_03888_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _35582_ (_03889_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _35583_ (_03890_, _03889_, _03888_);
  and _35584_ (_03891_, _03890_, _00228_);
  or _35585_ (_03892_, _03891_, _03887_);
  or _35586_ (_03893_, _03892_, _03881_);
  or _35587_ (_03894_, _03893_, _03873_);
  and _35588_ (_03895_, _03894_, _03705_);
  and _35589_ (_03896_, _00051_, _00090_);
  and _35590_ (_03897_, _00027_, _00143_);
  and _35591_ (_03898_, _03897_, _26816_);
  and _35592_ (_03899_, _23818_, _23824_);
  or _35593_ (_03901_, _23815_, _26723_);
  nor _35594_ (_03902_, _03901_, _03899_);
  not _35595_ (_03903_, _26732_);
  not _35596_ (_03904_, _23826_);
  not _35597_ (_03905_, _26699_);
  and _35598_ (_03906_, _23838_, _23810_);
  nor _35599_ (_03908_, _03906_, _03905_);
  and _35600_ (_03909_, _03908_, _03904_);
  and _35601_ (_03910_, _03909_, _03903_);
  and _35602_ (_03911_, _03910_, _03902_);
  and _35603_ (_03912_, _26720_, _23834_);
  and _35604_ (_03913_, _03912_, _03911_);
  or _35605_ (_03914_, _23806_, _23801_);
  and _35606_ (_03915_, _03914_, _23824_);
  not _35607_ (_03916_, _03915_);
  nor _35608_ (_03917_, _26757_, _23840_);
  not _35609_ (_03919_, _03917_);
  nor _35610_ (_03920_, _03919_, _26735_);
  and _35611_ (_03922_, _03920_, _03916_);
  and _35612_ (_03923_, _03922_, _26745_);
  and _35613_ (_03925_, _03923_, _03913_);
  nor _35614_ (_03926_, _03925_, _24279_);
  nor _35615_ (_03927_, _03926_, p0_in[0]);
  and _35616_ (_03928_, _03926_, _25360_);
  nor _35617_ (_03929_, _03928_, _03927_);
  or _35618_ (_03930_, _03929_, _03874_);
  nor _35619_ (_03931_, _03926_, p0_in[4]);
  and _35620_ (_03933_, _03926_, _25409_);
  nor _35621_ (_03934_, _03933_, _03931_);
  or _35622_ (_03935_, _03934_, _00228_);
  and _35623_ (_03936_, _03935_, _03870_);
  and _35624_ (_03937_, _03936_, _03930_);
  nor _35625_ (_03938_, _03926_, p0_in[3]);
  not _35626_ (_03939_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _35627_ (_03940_, _03926_, _03939_);
  nor _35628_ (_03941_, _03940_, _03938_);
  or _35629_ (_03942_, _03941_, _03874_);
  nor _35630_ (_03943_, _03926_, p0_in[7]);
  not _35631_ (_03944_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _35632_ (_03945_, _03926_, _03944_);
  nor _35633_ (_03946_, _03945_, _03943_);
  or _35634_ (_03947_, _03946_, _00228_);
  and _35635_ (_03949_, _03947_, _03878_);
  and _35636_ (_03950_, _03949_, _03942_);
  or _35637_ (_03951_, _03950_, _03937_);
  nor _35638_ (_03952_, _03926_, p0_in[1]);
  and _35639_ (_03953_, _03926_, _25347_);
  nor _35640_ (_03954_, _03953_, _03952_);
  or _35641_ (_03955_, _03954_, _03874_);
  or _35642_ (_03956_, _03926_, p0_in[5]);
  not _35643_ (_03957_, _03926_);
  or _35644_ (_03958_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _35645_ (_03959_, _03958_, _03956_);
  or _35646_ (_03960_, _03959_, _00228_);
  and _35647_ (_03962_, _03960_, _03876_);
  and _35648_ (_03963_, _03962_, _03955_);
  nor _35649_ (_03964_, _03926_, p0_in[2]);
  and _35650_ (_03965_, _03926_, _25333_);
  nor _35651_ (_03966_, _03965_, _03964_);
  or _35652_ (_03967_, _03966_, _03874_);
  nor _35653_ (_03968_, _03926_, p0_in[6]);
  and _35654_ (_03970_, _03926_, _25392_);
  nor _35655_ (_03972_, _03970_, _03968_);
  or _35656_ (_03973_, _03972_, _00228_);
  and _35657_ (_03975_, _03973_, _03883_);
  and _35658_ (_03976_, _03975_, _03967_);
  or _35659_ (_03977_, _03976_, _03963_);
  or _35660_ (_03978_, _03977_, _03951_);
  and _35661_ (_03979_, _03978_, _03898_);
  nor _35662_ (_03980_, _03926_, p1_in[0]);
  and _35663_ (_03981_, _03926_, _25277_);
  nor _35664_ (_03982_, _03981_, _03980_);
  or _35665_ (_03983_, _03982_, _03874_);
  nor _35666_ (_03984_, _03926_, p1_in[4]);
  not _35667_ (_03985_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _35668_ (_03987_, _03926_, _03985_);
  nor _35669_ (_03988_, _03987_, _03984_);
  or _35670_ (_03990_, _03988_, _00228_);
  and _35671_ (_03991_, _03990_, _03870_);
  and _35672_ (_03993_, _03991_, _03983_);
  nor _35673_ (_03995_, _03926_, p1_in[3]);
  and _35674_ (_03996_, _03926_, _25234_);
  nor _35675_ (_03997_, _03996_, _03995_);
  or _35676_ (_03998_, _03997_, _03874_);
  nor _35677_ (_04000_, _03926_, p1_in[7]);
  not _35678_ (_04001_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _35679_ (_04003_, _03926_, _04001_);
  nor _35680_ (_04004_, _04003_, _04000_);
  or _35681_ (_04006_, _04004_, _00228_);
  and _35682_ (_04008_, _04006_, _03878_);
  and _35683_ (_04009_, _04008_, _03998_);
  or _35684_ (_04011_, _04009_, _03993_);
  nor _35685_ (_04012_, _03926_, p1_in[1]);
  and _35686_ (_04014_, _03926_, _25263_);
  nor _35687_ (_04016_, _04014_, _04012_);
  or _35688_ (_04017_, _04016_, _03874_);
  or _35689_ (_04018_, _03926_, p1_in[5]);
  or _35690_ (_04019_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _35691_ (_04020_, _04019_, _04018_);
  or _35692_ (_04021_, _04020_, _00228_);
  and _35693_ (_04022_, _04021_, _03876_);
  and _35694_ (_04023_, _04022_, _04017_);
  nor _35695_ (_04024_, _03926_, p1_in[2]);
  and _35696_ (_04025_, _03926_, _25250_);
  nor _35697_ (_04027_, _04025_, _04024_);
  or _35698_ (_04028_, _04027_, _03874_);
  nor _35699_ (_04029_, _03926_, p1_in[6]);
  and _35700_ (_04030_, _03926_, _25295_);
  nor _35701_ (_04031_, _04030_, _04029_);
  or _35702_ (_04032_, _04031_, _00228_);
  and _35703_ (_04033_, _04032_, _03883_);
  and _35704_ (_04034_, _04033_, _04028_);
  or _35705_ (_04035_, _04034_, _04023_);
  or _35706_ (_04036_, _04035_, _04011_);
  and _35707_ (_04038_, _04036_, _03703_);
  not _35708_ (_04039_, _26816_);
  and _35709_ (_04041_, _03702_, _04039_);
  and _35710_ (_04042_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor _35711_ (_04043_, _00228_, _02660_);
  or _35712_ (_04045_, _04043_, _04042_);
  and _35713_ (_04047_, _04045_, _03878_);
  nor _35714_ (_04048_, _00228_, _02674_);
  and _35715_ (_04049_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _35716_ (_04051_, _04049_, _04048_);
  and _35717_ (_04052_, _04051_, _03883_);
  or _35718_ (_04053_, _04052_, _04047_);
  and _35719_ (_04054_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  not _35720_ (_04056_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _35721_ (_04057_, _00228_, _04056_);
  or _35722_ (_04058_, _04057_, _04054_);
  and _35723_ (_04059_, _04058_, _03870_);
  and _35724_ (_04060_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor _35725_ (_04061_, _00228_, _02604_);
  or _35726_ (_04062_, _04061_, _04060_);
  and _35727_ (_04063_, _04062_, _03876_);
  or _35728_ (_04064_, _04063_, _04059_);
  or _35729_ (_04065_, _04064_, _04053_);
  and _35730_ (_04066_, _04065_, _04041_);
  or _35731_ (_04067_, _04066_, _04038_);
  or _35732_ (_04069_, _04067_, _03979_);
  and _35733_ (_04070_, _04069_, _03896_);
  and _35734_ (_04071_, _03897_, _04039_);
  and _35735_ (_04073_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _35736_ (_04074_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _35737_ (_04076_, _04074_, _04073_);
  and _35738_ (_04078_, _04076_, _03878_);
  or _35739_ (_04079_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or _35740_ (_04080_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _35741_ (_04081_, _04080_, _03870_);
  and _35742_ (_04082_, _04081_, _04079_);
  or _35743_ (_04083_, _04082_, _04078_);
  nor _35744_ (_04084_, _00228_, _02243_);
  and _35745_ (_04085_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _35746_ (_04086_, _04085_, _04084_);
  and _35747_ (_04088_, _04086_, _03883_);
  or _35748_ (_04090_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  not _35749_ (_04091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand _35750_ (_04093_, _00228_, _04091_);
  and _35751_ (_04094_, _04093_, _03876_);
  and _35752_ (_04095_, _04094_, _04090_);
  or _35753_ (_04096_, _04095_, _04088_);
  or _35754_ (_04098_, _04096_, _04083_);
  and _35755_ (_04099_, _04098_, _03896_);
  and _35756_ (_04100_, _03698_, _00090_);
  and _35757_ (_04102_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _35758_ (_04103_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _35759_ (_04104_, _04103_, _04102_);
  and _35760_ (_04105_, _04104_, _03878_);
  or _35761_ (_04106_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _35762_ (_04108_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _35763_ (_04110_, _04108_, _03870_);
  and _35764_ (_04111_, _04110_, _04106_);
  or _35765_ (_04113_, _04111_, _04105_);
  and _35766_ (_04114_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _35767_ (_04115_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _35768_ (_04117_, _04115_, _04114_);
  and _35769_ (_04118_, _04117_, _03883_);
  or _35770_ (_04119_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _35771_ (_04120_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _35772_ (_04121_, _04120_, _03876_);
  and _35773_ (_04122_, _04121_, _04119_);
  or _35774_ (_04123_, _04122_, _04118_);
  or _35775_ (_04124_, _04123_, _04113_);
  and _35776_ (_04125_, _04124_, _04100_);
  or _35777_ (_04127_, _04125_, _04099_);
  and _35778_ (_04128_, _04127_, _04071_);
  nor _35779_ (_04129_, _03926_, p3_in[0]);
  and _35780_ (_04130_, _03926_, _25074_);
  nor _35781_ (_04131_, _04130_, _04129_);
  or _35782_ (_04132_, _04131_, _03874_);
  nor _35783_ (_04133_, _03926_, p3_in[4]);
  not _35784_ (_04134_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _35785_ (_04135_, _03926_, _04134_);
  nor _35786_ (_04136_, _04135_, _04133_);
  or _35787_ (_04138_, _04136_, _00228_);
  and _35788_ (_04139_, _04138_, _03870_);
  and _35789_ (_04140_, _04139_, _04132_);
  nor _35790_ (_04141_, _03926_, p3_in[3]);
  and _35791_ (_04142_, _03926_, _25033_);
  nor _35792_ (_04143_, _04142_, _04141_);
  or _35793_ (_04144_, _04143_, _03874_);
  nor _35794_ (_04145_, _03926_, p3_in[7]);
  not _35795_ (_04146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _35796_ (_04147_, _03926_, _04146_);
  nor _35797_ (_04148_, _04147_, _04145_);
  or _35798_ (_04149_, _04148_, _00228_);
  and _35799_ (_04150_, _04149_, _03878_);
  and _35800_ (_04151_, _04150_, _04144_);
  or _35801_ (_04152_, _04151_, _04140_);
  nor _35802_ (_04153_, _03926_, p3_in[1]);
  and _35803_ (_04154_, _03926_, _25062_);
  nor _35804_ (_04155_, _04154_, _04153_);
  or _35805_ (_04156_, _04155_, _03874_);
  or _35806_ (_04157_, _03926_, p3_in[5]);
  or _35807_ (_04158_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _35808_ (_04160_, _04158_, _04157_);
  or _35809_ (_04161_, _04160_, _00228_);
  and _35810_ (_04163_, _04161_, _03876_);
  and _35811_ (_04164_, _04163_, _04156_);
  nor _35812_ (_04166_, _03926_, p3_in[2]);
  and _35813_ (_04167_, _03926_, _25049_);
  nor _35814_ (_04169_, _04167_, _04166_);
  or _35815_ (_04170_, _04169_, _03874_);
  nor _35816_ (_04172_, _03926_, p3_in[6]);
  and _35817_ (_04173_, _03926_, _25098_);
  nor _35818_ (_04175_, _04173_, _04172_);
  or _35819_ (_04176_, _04175_, _00228_);
  and _35820_ (_04178_, _04176_, _03883_);
  and _35821_ (_04179_, _04178_, _04170_);
  or _35822_ (_04180_, _04179_, _04164_);
  or _35823_ (_04181_, _04180_, _04152_);
  and _35824_ (_04182_, _04181_, _03703_);
  nor _35825_ (_04183_, _03926_, p2_in[0]);
  and _35826_ (_04184_, _03926_, _25200_);
  nor _35827_ (_04186_, _04184_, _04183_);
  or _35828_ (_04188_, _04186_, _03874_);
  nor _35829_ (_04190_, _03926_, p2_in[4]);
  and _35830_ (_04192_, _03926_, _25160_);
  nor _35831_ (_04193_, _04192_, _04190_);
  or _35832_ (_04195_, _04193_, _00228_);
  and _35833_ (_04196_, _04195_, _03870_);
  and _35834_ (_04197_, _04196_, _04188_);
  nor _35835_ (_04199_, _03926_, p2_in[3]);
  and _35836_ (_04201_, _03926_, _25175_);
  nor _35837_ (_04202_, _04201_, _04199_);
  or _35838_ (_04203_, _04202_, _03874_);
  nor _35839_ (_04204_, _03926_, p2_in[7]);
  not _35840_ (_04206_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _35841_ (_04207_, _03926_, _04206_);
  nor _35842_ (_04209_, _04207_, _04204_);
  or _35843_ (_04210_, _04209_, _00228_);
  and _35844_ (_04211_, _04210_, _03878_);
  and _35845_ (_04212_, _04211_, _04203_);
  or _35846_ (_04213_, _04212_, _04197_);
  nor _35847_ (_04214_, _03926_, p2_in[1]);
  and _35848_ (_04215_, _03926_, _25135_);
  nor _35849_ (_04216_, _04215_, _04214_);
  or _35850_ (_04217_, _04216_, _03874_);
  or _35851_ (_04219_, _03926_, p2_in[5]);
  or _35852_ (_04220_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _35853_ (_04221_, _04220_, _04219_);
  or _35854_ (_04222_, _04221_, _00228_);
  and _35855_ (_04223_, _04222_, _03876_);
  and _35856_ (_04224_, _04223_, _04217_);
  nor _35857_ (_04225_, _03926_, p2_in[2]);
  and _35858_ (_04226_, _03926_, _25188_);
  nor _35859_ (_04227_, _04226_, _04225_);
  or _35860_ (_04228_, _04227_, _03874_);
  nor _35861_ (_04229_, _03926_, p2_in[6]);
  not _35862_ (_04230_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _35863_ (_04231_, _03926_, _04230_);
  nor _35864_ (_04232_, _04231_, _04229_);
  or _35865_ (_04233_, _04232_, _00228_);
  and _35866_ (_04234_, _04233_, _03883_);
  and _35867_ (_04235_, _04234_, _04228_);
  or _35868_ (_04236_, _04235_, _04224_);
  or _35869_ (_04237_, _04236_, _04213_);
  and _35870_ (_04238_, _04237_, _03898_);
  or _35871_ (_04239_, _04238_, _04182_);
  and _35872_ (_04240_, _04239_, _04100_);
  nor _35873_ (_04241_, _00051_, _00090_);
  and _35874_ (_04242_, _04241_, _03898_);
  and _35875_ (_04243_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _35876_ (_04244_, _00228_, _23109_);
  or _35877_ (_04245_, _04244_, _04243_);
  and _35878_ (_04246_, _04245_, _03876_);
  nand _35879_ (_04247_, _00228_, _23210_);
  or _35880_ (_04248_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _35881_ (_04249_, _04248_, _03883_);
  and _35882_ (_04250_, _04249_, _04247_);
  nor _35883_ (_04251_, _00228_, _23034_);
  and _35884_ (_04252_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _35885_ (_04253_, _04252_, _04251_);
  and _35886_ (_04255_, _04253_, _03878_);
  or _35887_ (_04256_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _35888_ (_04257_, _00228_, _23291_);
  and _35889_ (_04258_, _04257_, _03870_);
  and _35890_ (_04259_, _04258_, _04256_);
  or _35891_ (_04260_, _04259_, _04255_);
  or _35892_ (_04261_, _04260_, _04250_);
  or _35893_ (_04263_, _04261_, _04246_);
  and _35894_ (_04264_, _04263_, _04242_);
  nand _35895_ (_04265_, _00143_, _00090_);
  or _35896_ (_04266_, _04265_, _26816_);
  not _35897_ (_04267_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _35898_ (_04268_, _03703_, _04267_);
  and _35899_ (_04270_, _04268_, _04266_);
  and _35900_ (_04272_, _04071_, _03699_);
  not _35901_ (_04274_, _03699_);
  and _35902_ (_04275_, _03898_, _04274_);
  nor _35903_ (_04276_, _04275_, _04272_);
  and _35904_ (_04277_, _04276_, _04270_);
  and _35905_ (_04278_, _04100_, _04041_);
  or _35906_ (_04280_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand _35907_ (_04281_, _00228_, _24789_);
  and _35908_ (_04283_, _04281_, _03878_);
  and _35909_ (_04285_, _04283_, _04280_);
  and _35910_ (_04286_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _35911_ (_04287_, _00228_, _24786_);
  or _35912_ (_04288_, _04287_, _04286_);
  and _35913_ (_04289_, _04288_, _03876_);
  or _35914_ (_04290_, _04289_, _04285_);
  and _35915_ (_04291_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor _35916_ (_04292_, _00228_, _24784_);
  or _35917_ (_04293_, _04292_, _04291_);
  and _35918_ (_04295_, _04293_, _03870_);
  nand _35919_ (_04297_, _00228_, _24800_);
  or _35920_ (_04298_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _35921_ (_04300_, _04298_, _03883_);
  and _35922_ (_04301_, _04300_, _04297_);
  or _35923_ (_04302_, _04301_, _04295_);
  or _35924_ (_04303_, _04302_, _04290_);
  and _35925_ (_04304_, _04303_, _04278_);
  and _35926_ (_04305_, _04241_, _03703_);
  and _35927_ (_04306_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not _35928_ (_04308_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor _35929_ (_04309_, _00228_, _04308_);
  or _35930_ (_04311_, _04309_, _04306_);
  and _35931_ (_04312_, _04311_, _03878_);
  and _35932_ (_04314_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not _35933_ (_04315_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor _35934_ (_04317_, _00228_, _04315_);
  or _35935_ (_04319_, _04317_, _04314_);
  and _35936_ (_04320_, _04319_, _03876_);
  or _35937_ (_04322_, _04320_, _04312_);
  and _35938_ (_04323_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _35939_ (_04325_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor _35940_ (_04326_, _00228_, _04325_);
  or _35941_ (_04327_, _04326_, _04323_);
  and _35942_ (_04328_, _04327_, _03870_);
  not _35943_ (_04329_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor _35944_ (_04330_, _00228_, _04329_);
  and _35945_ (_04331_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _35946_ (_04332_, _04331_, _04330_);
  and _35947_ (_04333_, _04332_, _03883_);
  or _35948_ (_04334_, _04333_, _04328_);
  or _35949_ (_04335_, _04334_, _04322_);
  and _35950_ (_04336_, _04335_, _04305_);
  or _35951_ (_04337_, _04336_, _04304_);
  or _35952_ (_04338_, _04337_, _04277_);
  or _35953_ (_04339_, _04338_, _04264_);
  and _35954_ (_04340_, _00235_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _35955_ (_04341_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _35956_ (_04342_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _35957_ (_04343_, _00228_, _04342_);
  or _35958_ (_04344_, _04343_, _04341_);
  and _35959_ (_04345_, _04344_, _03876_);
  or _35960_ (_04347_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _35961_ (_04348_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _35962_ (_04349_, _04348_, _03883_);
  and _35963_ (_04350_, _04349_, _04347_);
  and _35964_ (_04352_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _35965_ (_04353_, _00228_, _25483_);
  or _35966_ (_04355_, _04353_, _04352_);
  and _35967_ (_04356_, _04355_, _03878_);
  or _35968_ (_04357_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _35969_ (_04358_, _00228_, _25527_);
  and _35970_ (_04360_, _04358_, _03870_);
  and _35971_ (_04361_, _04360_, _04357_);
  or _35972_ (_04362_, _04361_, _04356_);
  or _35973_ (_04363_, _04362_, _04350_);
  or _35974_ (_04364_, _04363_, _04345_);
  and _35975_ (_04366_, _04364_, _04272_);
  or _35976_ (_04367_, _04366_, _04340_);
  or _35977_ (_04368_, _04367_, _04339_);
  or _35978_ (_04370_, _04368_, _04240_);
  or _35979_ (_04372_, _04370_, _04128_);
  or _35980_ (_04373_, _04372_, _04070_);
  or _35981_ (_04374_, _04373_, _03895_);
  and _35982_ (_04375_, _04242_, _00322_);
  nor _35983_ (_04376_, _04375_, _00151_);
  nand _35984_ (_04377_, _04340_, _23504_);
  and _35985_ (_04378_, _04377_, _04376_);
  and _35986_ (_04379_, _04378_, _04374_);
  nor _35987_ (_04380_, _00228_, _24043_);
  and _35988_ (_04382_, _00228_, _02728_);
  or _35989_ (_04383_, _04382_, _04380_);
  and _35990_ (_04384_, _04383_, _03876_);
  or _35991_ (_04385_, _00228_, _02450_);
  or _35992_ (_04387_, _03874_, _23880_);
  and _35993_ (_04388_, _04387_, _03883_);
  and _35994_ (_04389_, _04388_, _04385_);
  nor _35995_ (_04390_, _00228_, _23989_);
  and _35996_ (_04392_, _00228_, _23577_);
  or _35997_ (_04394_, _04392_, _04390_);
  and _35998_ (_04395_, _04394_, _03878_);
  nand _35999_ (_04396_, _00228_, _24210_);
  or _36000_ (_04397_, _00228_, _02700_);
  and _36001_ (_04399_, _04397_, _03870_);
  and _36002_ (_04400_, _04399_, _04396_);
  or _36003_ (_04401_, _04400_, _04395_);
  or _36004_ (_04402_, _04401_, _04389_);
  nor _36005_ (_04403_, _04402_, _04384_);
  nor _36006_ (_04404_, _04403_, _04376_);
  or _36007_ (_04405_, _04404_, _04379_);
  and _36008_ (_27316_, _04405_, _22731_);
  and _36009_ (_04406_, _24539_, _22844_);
  and _36010_ (_04407_, _03878_, _03874_);
  not _36011_ (_04409_, _04407_);
  and _36012_ (_04410_, _04409_, _04406_);
  and _36013_ (_04412_, _04410_, _00149_);
  not _36014_ (_04413_, _00143_);
  nor _36015_ (_04414_, _04413_, _00090_);
  and _36016_ (_04416_, _00228_, _26816_);
  and _36017_ (_04418_, _04416_, _03870_);
  nor _36018_ (_04419_, _00051_, _03700_);
  and _36019_ (_04420_, _04419_, _04418_);
  and _36020_ (_04421_, _04420_, _04414_);
  and _36021_ (_04423_, _04421_, _00322_);
  or _36022_ (_04425_, _04423_, _00237_);
  or _36023_ (_04426_, _04425_, _04412_);
  and _36024_ (_04427_, _04421_, _00319_);
  and _36025_ (_04428_, _00051_, _03700_);
  and _36026_ (_04429_, _04428_, _04418_);
  and _36027_ (_04430_, _04429_, _04414_);
  and _36028_ (_04431_, _04430_, _00312_);
  and _36029_ (_04433_, _00318_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _36030_ (_04434_, _03897_, _03896_);
  and _36031_ (_04435_, _04434_, _03878_);
  and _36032_ (_04436_, _04435_, _04416_);
  and _36033_ (_04437_, _04436_, _04433_);
  or _36034_ (_04438_, _04437_, _04431_);
  nor _36035_ (_04439_, _04438_, _04427_);
  nor _36036_ (_04440_, _04439_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _36037_ (_04441_, _04440_, _04426_);
  and _36038_ (_04442_, _04434_, _03883_);
  and _36039_ (_04443_, _04442_, _04416_);
  and _36040_ (_04444_, _04443_, _04433_);
  nor _36041_ (_04446_, _04444_, rst);
  and _36042_ (_27317_, _04446_, _04441_);
  not _36043_ (_04447_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _36044_ (_04448_, _03897_, _03699_);
  nor _36045_ (_04449_, _00228_, _26816_);
  and _36046_ (_04450_, _04449_, _03870_);
  and _36047_ (_04451_, _04450_, _04448_);
  and _36048_ (_04452_, _00228_, _04039_);
  and _36049_ (_04454_, _04452_, _03870_);
  and _36050_ (_04456_, _04454_, _04448_);
  nor _36051_ (_04458_, _04456_, _04451_);
  and _36052_ (_04459_, _04449_, _03876_);
  and _36053_ (_04461_, _04459_, _04448_);
  and _36054_ (_04462_, _04452_, _03883_);
  and _36055_ (_04463_, _04462_, _04448_);
  nor _36056_ (_04464_, _04463_, _04461_);
  and _36057_ (_04465_, _04464_, _04458_);
  and _36058_ (_04466_, _04454_, _04434_);
  and _36059_ (_04467_, _04452_, _03878_);
  and _36060_ (_04468_, _04467_, _04448_);
  nor _36061_ (_04469_, _04468_, _04466_);
  and _36062_ (_04470_, _04407_, _26816_);
  and _36063_ (_04472_, _04100_, _03702_);
  and _36064_ (_04474_, _04472_, _04470_);
  and _36065_ (_04475_, _04100_, _03897_);
  and _36066_ (_04476_, _04475_, _04454_);
  nor _36067_ (_04477_, _04476_, _04474_);
  and _36068_ (_04478_, _04477_, _04469_);
  and _36069_ (_04479_, _04478_, _04465_);
  and _36070_ (_04480_, _04467_, _04434_);
  and _36071_ (_04481_, _04452_, _03876_);
  and _36072_ (_04482_, _04481_, _04434_);
  nor _36073_ (_04483_, _04482_, _04480_);
  and _36074_ (_04484_, _04459_, _04434_);
  and _36075_ (_04485_, _04462_, _04434_);
  nor _36076_ (_04486_, _04485_, _04484_);
  and _36077_ (_04488_, _04486_, _04483_);
  and _36078_ (_04489_, _04470_, _04434_);
  and _36079_ (_04491_, _04450_, _04434_);
  nor _36080_ (_04493_, _04491_, _04489_);
  and _36081_ (_04494_, _03896_, _03702_);
  and _36082_ (_04495_, _04494_, _04454_);
  and _36083_ (_04496_, _04481_, _04494_);
  nor _36084_ (_04497_, _04496_, _04495_);
  and _36085_ (_04498_, _04497_, _04493_);
  and _36086_ (_04499_, _04498_, _04488_);
  and _36087_ (_04500_, _04499_, _04479_);
  not _36088_ (_04501_, _04418_);
  or _36089_ (_04502_, _04501_, _04265_);
  and _36090_ (_04503_, _04416_, _03878_);
  and _36091_ (_04505_, _04503_, _04434_);
  nor _36092_ (_04507_, _04443_, _04505_);
  and _36093_ (_04508_, _04241_, _03702_);
  and _36094_ (_04510_, _04508_, _04418_);
  and _36095_ (_04512_, _04416_, _03876_);
  and _36096_ (_04513_, _04512_, _04434_);
  nor _36097_ (_04514_, _04513_, _04510_);
  and _36098_ (_04516_, _04514_, _04507_);
  and _36099_ (_04517_, _04516_, _04502_);
  nor _36100_ (_04518_, _04430_, _04421_);
  and _36101_ (_04519_, _04518_, _04517_);
  and _36102_ (_04520_, _04519_, _04500_);
  nor _36103_ (_04521_, _04520_, _04441_);
  nor _36104_ (_04522_, _04521_, _04447_);
  not _36105_ (_04523_, _04444_);
  nand _36106_ (_04524_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _36107_ (_04526_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _36108_ (_04527_, _04526_, _04524_);
  nand _36109_ (_04528_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand _36110_ (_04529_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _36111_ (_04530_, _04529_, _04528_);
  and _36112_ (_04531_, _04530_, _04527_);
  nand _36113_ (_04532_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _36114_ (_04533_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _36115_ (_04534_, _04533_, _04532_);
  nand _36116_ (_04535_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nand _36117_ (_04536_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _36118_ (_04537_, _04536_, _04535_);
  and _36119_ (_04538_, _04537_, _04534_);
  and _36120_ (_04539_, _04538_, _04531_);
  nand _36121_ (_04540_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand _36122_ (_04541_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _36123_ (_04542_, _04541_, _04540_);
  nand _36124_ (_04543_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _36125_ (_04544_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _36126_ (_04545_, _04544_, _04543_);
  and _36127_ (_04547_, _04545_, _04542_);
  nand _36128_ (_04548_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand _36129_ (_04549_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _36130_ (_04550_, _04549_, _04548_);
  nand _36131_ (_04551_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _36132_ (_04552_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _36133_ (_04553_, _04552_, _04551_);
  and _36134_ (_04554_, _04553_, _04550_);
  and _36135_ (_04555_, _04554_, _04547_);
  and _36136_ (_04556_, _04555_, _04539_);
  nand _36137_ (_04557_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand _36138_ (_04558_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _36139_ (_04559_, _04558_, _04557_);
  nand _36140_ (_04560_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _36141_ (_04561_, _04513_, _00105_);
  and _36142_ (_04563_, _04561_, _04560_);
  and _36143_ (_04564_, _04563_, _04559_);
  and _36144_ (_04565_, _04475_, _04418_);
  nand _36145_ (_04566_, _04565_, _04209_);
  and _36146_ (_04567_, _04472_, _04418_);
  nand _36147_ (_04568_, _04567_, _04148_);
  and _36148_ (_04569_, _04568_, _04566_);
  and _36149_ (_04570_, _04434_, _04418_);
  nand _36150_ (_04572_, _04570_, _03946_);
  and _36151_ (_04573_, _04494_, _04418_);
  nand _36152_ (_04574_, _04573_, _04004_);
  and _36153_ (_04575_, _04574_, _04572_);
  and _36154_ (_04577_, _04575_, _04569_);
  and _36155_ (_04578_, _04577_, _04564_);
  nand _36156_ (_04579_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand _36157_ (_04580_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _36158_ (_04581_, _04580_, _04579_);
  and _36159_ (_04582_, _04581_, _04578_);
  and _36160_ (_04583_, _04582_, _04556_);
  or _36161_ (_04584_, _04583_, _04441_);
  nand _36162_ (_04585_, _04584_, _04523_);
  or _36163_ (_04586_, _04585_, _04522_);
  or _36164_ (_04587_, _04523_, _00883_);
  and _36165_ (_04589_, _04587_, _22731_);
  and _36166_ (_27318_[7], _04589_, _04586_);
  and _36167_ (_04590_, _03667_, _23583_);
  and _36168_ (_04592_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _36169_ (_25237_, _04592_, _04590_);
  and _36170_ (_04593_, _03667_, _23887_);
  and _36171_ (_04594_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _36172_ (_25239_, _04594_, _04593_);
  and _36173_ (_04595_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _36174_ (_04596_, _03662_, _23548_);
  or _36175_ (_25245_, _04596_, _04595_);
  and _36176_ (_04597_, _03667_, _23996_);
  and _36177_ (_04598_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _36178_ (_25265_, _04598_, _04597_);
  and _36179_ (_04599_, _03667_, _24134_);
  and _36180_ (_04601_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or _36181_ (_27228_, _04601_, _04599_);
  and _36182_ (_04602_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and _36183_ (_04603_, _03662_, _24134_);
  or _36184_ (_25273_, _04603_, _04602_);
  and _36185_ (_04604_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _36186_ (_04605_, _03662_, _24051_);
  or _36187_ (_25282_, _04605_, _04604_);
  and _36188_ (_04606_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _36189_ (_04607_, _03662_, _24089_);
  or _36190_ (_27095_, _04607_, _04606_);
  and _36191_ (_04608_, _02497_, _22974_);
  and _36192_ (_04609_, _04608_, _23996_);
  not _36193_ (_04610_, _04608_);
  and _36194_ (_04611_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _36195_ (_25304_, _04611_, _04609_);
  and _36196_ (_04612_, _04608_, _24134_);
  and _36197_ (_04613_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _36198_ (_25317_, _04613_, _04612_);
  and _36199_ (_04614_, _02512_, _24223_);
  not _36200_ (_04615_, _04614_);
  and _36201_ (_04616_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and _36202_ (_04617_, _04614_, _23887_);
  or _36203_ (_25324_, _04617_, _04616_);
  and _36204_ (_04619_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  and _36205_ (_04620_, _04614_, _24089_);
  or _36206_ (_25326_, _04620_, _04619_);
  and _36207_ (_04622_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and _36208_ (_04623_, _04614_, _23583_);
  or _36209_ (_25337_, _04623_, _04622_);
  and _36210_ (_04625_, _03667_, _24219_);
  and _36211_ (_04626_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _36212_ (_25348_, _04626_, _04625_);
  and _36213_ (_04627_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  and _36214_ (_04628_, _04614_, _24134_);
  or _36215_ (_25373_, _04628_, _04627_);
  and _36216_ (_04629_, _24219_, _24008_);
  and _36217_ (_04630_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or _36218_ (_25379_, _04630_, _04629_);
  and _36219_ (_04631_, _04608_, _23548_);
  and _36220_ (_04632_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _36221_ (_25389_, _04632_, _04631_);
  and _36222_ (_04633_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  and _36223_ (_04634_, _04614_, _23996_);
  or _36224_ (_27094_, _04634_, _04633_);
  and _36225_ (_04635_, _04608_, _24219_);
  and _36226_ (_04636_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _36227_ (_25399_, _04636_, _04635_);
  and _36228_ (_04637_, _04608_, _24089_);
  and _36229_ (_04638_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _36230_ (_25427_, _04638_, _04637_);
  and _36231_ (_04639_, _04608_, _23583_);
  and _36232_ (_04640_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _36233_ (_27213_, _04640_, _04639_);
  and _36234_ (_04641_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and _36235_ (_04642_, _04614_, _24219_);
  or _36236_ (_25437_, _04642_, _04641_);
  and _36237_ (_04643_, _04608_, _23887_);
  and _36238_ (_04644_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _36239_ (_25439_, _04644_, _04643_);
  and _36240_ (_04645_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and _36241_ (_04646_, _02836_, _23548_);
  or _36242_ (_25452_, _04646_, _04645_);
  and _36243_ (_04647_, _02497_, _24095_);
  and _36244_ (_04648_, _04647_, _24134_);
  not _36245_ (_04649_, _04647_);
  and _36246_ (_04650_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _36247_ (_25464_, _04650_, _04648_);
  and _36248_ (_04651_, _04647_, _24051_);
  and _36249_ (_04652_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _36250_ (_25468_, _04652_, _04651_);
  and _36251_ (_04653_, _02512_, _24095_);
  not _36252_ (_04654_, _04653_);
  and _36253_ (_04656_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _36254_ (_04657_, _04653_, _24219_);
  or _36255_ (_25471_, _04657_, _04656_);
  and _36256_ (_04658_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  and _36257_ (_04659_, _03011_, _23996_);
  or _36258_ (_25476_, _04659_, _04658_);
  and _36259_ (_04660_, _04647_, _23996_);
  and _36260_ (_04661_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _36261_ (_25498_, _04661_, _04660_);
  and _36262_ (_04662_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and _36263_ (_04663_, _04653_, _24089_);
  or _36264_ (_27092_, _04663_, _04662_);
  and _36265_ (_04665_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _36266_ (_04667_, _04653_, _23583_);
  or _36267_ (_25525_, _04667_, _04665_);
  and _36268_ (_04668_, _04647_, _23548_);
  and _36269_ (_04669_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _36270_ (_25530_, _04669_, _04668_);
  and _36271_ (_04670_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and _36272_ (_04671_, _04653_, _23887_);
  or _36273_ (_27091_, _04671_, _04670_);
  and _36274_ (_04672_, _04647_, _24219_);
  and _36275_ (_04673_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _36276_ (_25537_, _04673_, _04672_);
  and _36277_ (_04674_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  and _36278_ (_04675_, _03011_, _23583_);
  or _36279_ (_25555_, _04675_, _04674_);
  and _36280_ (_04676_, _04647_, _23583_);
  and _36281_ (_04677_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _36282_ (_25559_, _04677_, _04676_);
  and _36283_ (_04678_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and _36284_ (_04680_, _03011_, _23887_);
  or _36285_ (_25562_, _04680_, _04678_);
  and _36286_ (_04681_, _04647_, _23887_);
  and _36287_ (_04682_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _36288_ (_25570_, _04682_, _04681_);
  not _36289_ (_04683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _36290_ (_04684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _36291_ (_04685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor _36292_ (_04686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _36293_ (_04687_, _04686_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _36294_ (_04688_, _04687_, _04685_);
  and _36295_ (_04689_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02674_);
  or _36296_ (_04690_, _04689_, _04688_);
  nor _36297_ (_04691_, _04690_, _04684_);
  nand _36298_ (_04692_, _04691_, _04683_);
  nor _36299_ (_04693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor _36300_ (_04694_, _04693_, _04691_);
  nand _36301_ (_04695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _36302_ (_04696_, _04695_, _04694_);
  and _36303_ (_04697_, _04696_, _22731_);
  and _36304_ (_25638_, _04697_, _04692_);
  and _36305_ (_04698_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  and _36306_ (_04699_, _03011_, _24134_);
  or _36307_ (_25641_, _04699_, _04698_);
  not _36308_ (_04700_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and _36309_ (_04701_, _02652_, _04700_);
  and _36310_ (_04702_, _04701_, _02755_);
  and _36311_ (_04703_, _04702_, _02752_);
  nand _36312_ (_04704_, _04703_, _02648_);
  not _36313_ (_04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _36314_ (_04706_, _02757_, _04705_);
  and _36315_ (_04707_, _04706_, _04704_);
  or _36316_ (_04708_, _04707_, _02658_);
  and _36317_ (_25646_, _04708_, _22731_);
  and _36318_ (_04709_, _02497_, _24372_);
  and _36319_ (_04710_, _04709_, _24089_);
  not _36320_ (_04711_, _04709_);
  and _36321_ (_04712_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _36322_ (_25653_, _04712_, _04710_);
  and _36323_ (_25655_, _04694_, _22731_);
  and _36324_ (_04714_, _04709_, _23583_);
  and _36325_ (_04715_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _36326_ (_25667_, _04715_, _04714_);
  and _36327_ (_04716_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and _36328_ (_04718_, _03011_, _24051_);
  or _36329_ (_25671_, _04718_, _04716_);
  and _36330_ (_04719_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  and _36331_ (_04721_, _03011_, _24089_);
  or _36332_ (_25676_, _04721_, _04719_);
  and _36333_ (_04722_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or _36334_ (_04723_, _04722_, _02658_);
  nor _36335_ (_04724_, _02675_, rst);
  and _36336_ (_25678_, _04724_, _04723_);
  nand _36337_ (_04725_, _02910_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or _36338_ (_04726_, _02910_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _36339_ (_04727_, _04726_, _22731_);
  nand _36340_ (_04729_, _04727_, _04725_);
  nor _36341_ (_25680_, _04729_, _02658_);
  not _36342_ (_04730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _36343_ (_04732_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _36344_ (_04733_, _04687_, _04342_);
  or _36345_ (_04735_, _04733_, _04689_);
  nor _36346_ (_04736_, _04735_, _04732_);
  nand _36347_ (_04737_, _04736_, _04730_);
  nor _36348_ (_04738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _36349_ (_04739_, _04738_, _04736_);
  nand _36350_ (_04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _36351_ (_04742_, _04741_, _04739_);
  and _36352_ (_04743_, _04742_, _22731_);
  and _36353_ (_25688_, _04743_, _04737_);
  and _36354_ (_25690_, _04739_, _22731_);
  and _36355_ (_04744_, _04709_, _23996_);
  and _36356_ (_04745_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _36357_ (_27189_, _04745_, _04744_);
  and _36358_ (_04747_, _04709_, _24134_);
  and _36359_ (_04748_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _36360_ (_25702_, _04748_, _04747_);
  not _36361_ (_04749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor _36362_ (_04750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _04056_);
  not _36363_ (_04751_, _04750_);
  nor _36364_ (_04752_, _02568_, _02810_);
  and _36365_ (_04753_, _04752_, _04751_);
  and _36366_ (_04754_, _04753_, _02820_);
  nor _36367_ (_04755_, _04754_, _04749_);
  and _36368_ (_04756_, _04754_, rxd_i);
  or _36369_ (_04757_, _04756_, rst);
  or _36370_ (_25706_, _04757_, _04755_);
  or _36371_ (_04758_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _36372_ (_04759_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _36373_ (_04760_, _04759_, _02568_);
  or _36374_ (_04761_, _04760_, _02778_);
  nand _36375_ (_04762_, _04761_, _04758_);
  nand _36376_ (_25708_, _04762_, _02080_);
  and _36377_ (_04763_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _36378_ (_04764_, _04653_, _23996_);
  or _36379_ (_25717_, _04764_, _04763_);
  and _36380_ (_04766_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _36381_ (_04767_, _04653_, _24134_);
  or _36382_ (_25725_, _04767_, _04766_);
  and _36383_ (_04768_, _02497_, _24146_);
  and _36384_ (_04769_, _04768_, _24134_);
  not _36385_ (_04770_, _04768_);
  and _36386_ (_04772_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _36387_ (_25731_, _04772_, _04769_);
  and _36388_ (_04773_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _36389_ (_04774_, _04653_, _24051_);
  or _36390_ (_25733_, _04774_, _04773_);
  and _36391_ (_04775_, _04768_, _23996_);
  and _36392_ (_04777_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _36393_ (_25742_, _04777_, _04775_);
  and _36394_ (_04778_, _02502_, _23996_);
  and _36395_ (_04779_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _36396_ (_25747_, _04779_, _04778_);
  and _36397_ (_04781_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _36398_ (_04782_, _23687_);
  nor _36399_ (_04783_, _26748_, _04782_);
  and _36400_ (_04785_, _24257_, _23797_);
  or _36401_ (_04786_, _04785_, _01985_);
  nor _36402_ (_04787_, _23782_, _23749_);
  and _36403_ (_04789_, _04787_, _23838_);
  or _36404_ (_04790_, _04789_, _23897_);
  or _36405_ (_04791_, _04790_, _04786_);
  or _36406_ (_04792_, _04791_, _04783_);
  and _36407_ (_04793_, _23784_, _23687_);
  or _36408_ (_04794_, _01979_, _04793_);
  and _36409_ (_04795_, _23911_, _23687_);
  or _36410_ (_04796_, _03905_, _23841_);
  or _36411_ (_04797_, _04796_, _04795_);
  nor _36412_ (_04798_, _04797_, _04794_);
  nand _36413_ (_04799_, _04798_, _26733_);
  and _36414_ (_04800_, _23780_, _23772_);
  and _36415_ (_04801_, _26730_, _23687_);
  or _36416_ (_04802_, _04801_, _04800_);
  or _36417_ (_04803_, _26757_, _24259_);
  and _36418_ (_04804_, _04803_, _23791_);
  or _36419_ (_04806_, _04804_, _04802_);
  or _36420_ (_04807_, _04806_, _04799_);
  or _36421_ (_04808_, _04807_, _04792_);
  and _36422_ (_04809_, _04808_, _22737_);
  or _36423_ (_04810_, _04809_, _04781_);
  and _36424_ (_26847_[0], _04810_, _22731_);
  and _36425_ (_04812_, _24408_, _23941_);
  and _36426_ (_04813_, _04812_, _23996_);
  not _36427_ (_04815_, _04812_);
  and _36428_ (_04816_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _36429_ (_25762_, _04816_, _04813_);
  and _36430_ (_04818_, _04812_, _24051_);
  and _36431_ (_04819_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _36432_ (_25774_, _04819_, _04818_);
  and _36433_ (_04820_, _04812_, _23583_);
  and _36434_ (_04821_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _36435_ (_27138_, _04821_, _04820_);
  and _36436_ (_04823_, _24134_, _22983_);
  and _36437_ (_04824_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or _36438_ (_25847_, _04824_, _04823_);
  and _36439_ (_04825_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _36440_ (_04826_, _03319_, _23548_);
  or _36441_ (_25853_, _04826_, _04825_);
  and _36442_ (_04827_, _04709_, _24219_);
  and _36443_ (_04828_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _36444_ (_25857_, _04828_, _04827_);
  and _36445_ (_04829_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _36446_ (_04830_, _03319_, _24219_);
  or _36447_ (_25871_, _04830_, _04829_);
  and _36448_ (_04831_, _24518_, _23583_);
  and _36449_ (_04832_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or _36450_ (_25875_, _04832_, _04831_);
  and _36451_ (_04833_, _02432_, _24219_);
  and _36452_ (_04835_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  or _36453_ (_25883_, _04835_, _04833_);
  and _36454_ (_04837_, _04768_, _24219_);
  and _36455_ (_04838_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _36456_ (_25887_, _04838_, _04837_);
  and _36457_ (_04840_, _04768_, _23887_);
  and _36458_ (_04841_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _36459_ (_25889_, _04841_, _04840_);
  and _36460_ (_04843_, _04768_, _23548_);
  and _36461_ (_04844_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _36462_ (_25904_, _04844_, _04843_);
  and _36463_ (_04846_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _36464_ (_04847_, _03319_, _23887_);
  or _36465_ (_25906_, _04847_, _04846_);
  and _36466_ (_04848_, _03360_, _24219_);
  and _36467_ (_04849_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or _36468_ (_25927_, _04849_, _04848_);
  and _36469_ (_04851_, _04768_, _23583_);
  and _36470_ (_04852_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _36471_ (_27080_, _04852_, _04851_);
  and _36472_ (_04853_, _02039_, _24140_);
  not _36473_ (_04854_, _04853_);
  and _36474_ (_04855_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and _36475_ (_04856_, _04853_, _23583_);
  or _36476_ (_25939_, _04856_, _04855_);
  and _36477_ (_04858_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  and _36478_ (_04859_, _04853_, _23887_);
  or _36479_ (_25946_, _04859_, _04858_);
  and _36480_ (_04860_, _04768_, _24089_);
  and _36481_ (_04861_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or _36482_ (_25949_, _04861_, _04860_);
  and _36483_ (_04862_, _03360_, _23583_);
  and _36484_ (_04864_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _36485_ (_25953_, _04864_, _04862_);
  and _36486_ (_04865_, _03308_, _24056_);
  and _36487_ (_04866_, _04865_, _24134_);
  not _36488_ (_04867_, _04865_);
  and _36489_ (_04868_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or _36490_ (_25957_, _04868_, _04866_);
  and _36491_ (_04869_, _24518_, _24089_);
  and _36492_ (_04871_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or _36493_ (_25960_, _04871_, _04869_);
  and _36494_ (_04872_, _02432_, _24089_);
  and _36495_ (_04874_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  or _36496_ (_25966_, _04874_, _04872_);
  and _36497_ (_04875_, _02432_, _23887_);
  and _36498_ (_04876_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or _36499_ (_25972_, _04876_, _04875_);
  and _36500_ (_04877_, _03360_, _24051_);
  and _36501_ (_04878_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or _36502_ (_25993_, _04878_, _04877_);
  and _36503_ (_04879_, _02039_, _24319_);
  not _36504_ (_04880_, _04879_);
  and _36505_ (_04881_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _36506_ (_04882_, _04879_, _23548_);
  or _36507_ (_25996_, _04882_, _04881_);
  and _36508_ (_04884_, _03313_, _23887_);
  and _36509_ (_04885_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  or _36510_ (_26004_, _04885_, _04884_);
  and _36511_ (_04886_, _03313_, _24134_);
  and _36512_ (_04887_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  or _36513_ (_26009_, _04887_, _04886_);
  and _36514_ (_04888_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and _36515_ (_04890_, _04879_, _23887_);
  or _36516_ (_26012_, _04890_, _04888_);
  and _36517_ (_04891_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _36518_ (_04892_, _04879_, _24089_);
  or _36519_ (_26015_, _04892_, _04891_);
  and _36520_ (_04893_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _36521_ (_04894_, _04879_, _24051_);
  or _36522_ (_26019_, _04894_, _04893_);
  and _36523_ (_04895_, _03313_, _24051_);
  and _36524_ (_04896_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or _36525_ (_26026_, _04896_, _04895_);
  and _36526_ (_04897_, _02039_, _24146_);
  not _36527_ (_04898_, _04897_);
  and _36528_ (_04899_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _36529_ (_04900_, _04897_, _24089_);
  or _36530_ (_26029_, _04900_, _04899_);
  and _36531_ (_04901_, _03033_, _23548_);
  and _36532_ (_04902_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _36533_ (_26030_, _04902_, _04901_);
  and _36534_ (_04903_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and _36535_ (_04904_, _04897_, _24134_);
  or _36536_ (_26033_, _04904_, _04903_);
  and _36537_ (_04905_, _02039_, _24372_);
  not _36538_ (_04907_, _04905_);
  and _36539_ (_04908_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _36540_ (_04909_, _04905_, _23548_);
  or _36541_ (_27010_, _04909_, _04908_);
  and _36542_ (_04910_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _36543_ (_04912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _36544_ (_04913_, _22740_, _04912_);
  or _36545_ (_04915_, _04913_, _04910_);
  and _36546_ (_26862_[15], _04915_, _22731_);
  and _36547_ (_04916_, _03033_, _23583_);
  and _36548_ (_04918_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or _36549_ (_26046_, _04918_, _04916_);
  and _36550_ (_04920_, _24301_, _24236_);
  and _36551_ (_04921_, _04920_, _24051_);
  not _36552_ (_04923_, _04920_);
  and _36553_ (_04924_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _36554_ (_26052_, _04924_, _04921_);
  and _36555_ (_04925_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and _36556_ (_04926_, _04905_, _23583_);
  or _36557_ (_26056_, _04926_, _04925_);
  and _36558_ (_04928_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _36559_ (_04930_, _04905_, _24051_);
  or _36560_ (_26062_, _04930_, _04928_);
  and _36561_ (_04932_, _25672_, _23548_);
  and _36562_ (_04933_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _36563_ (_26065_, _04933_, _04932_);
  and _36564_ (_04935_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _36565_ (_04936_, _04905_, _23996_);
  or _36566_ (_26069_, _04936_, _04935_);
  and _36567_ (_04937_, _02039_, _24095_);
  not _36568_ (_04938_, _04937_);
  and _36569_ (_04939_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and _36570_ (_04940_, _04937_, _24219_);
  or _36571_ (_27012_, _04940_, _04939_);
  and _36572_ (_04941_, _03033_, _24219_);
  and _36573_ (_04942_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _36574_ (_26075_, _04942_, _04941_);
  and _36575_ (_04943_, _03001_, _24134_);
  and _36576_ (_04944_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _36577_ (_26078_, _04944_, _04943_);
  and _36578_ (_04946_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  and _36579_ (_04947_, _04937_, _23887_);
  or _36580_ (_26086_, _04947_, _04946_);
  and _36581_ (_04948_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and _36582_ (_04949_, _04937_, _24089_);
  or _36583_ (_26096_, _04949_, _04948_);
  and _36584_ (_04950_, _25413_, _22974_);
  and _36585_ (_04951_, _04950_, _24089_);
  not _36586_ (_04952_, _04950_);
  and _36587_ (_04953_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or _36588_ (_26105_, _04953_, _04951_);
  or _36589_ (_04955_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _36590_ (_04956_, _04955_, _22731_);
  nand _36591_ (_04957_, _02071_, _24082_);
  and _36592_ (_26109_, _04957_, _04956_);
  nor _36593_ (_27315_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _36594_ (_04959_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor _36595_ (_04961_, _03689_, rst);
  and _36596_ (_27315_[1], _04961_, _04959_);
  nor _36597_ (_04964_, _03689_, _03688_);
  or _36598_ (_04965_, _04964_, _03690_);
  and _36599_ (_04967_, _03693_, _22731_);
  and _36600_ (_27315_[2], _04967_, _04965_);
  and _36601_ (_04969_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and _36602_ (_04970_, _04937_, _24134_);
  or _36603_ (_26117_, _04970_, _04969_);
  nand _36604_ (_04971_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _36605_ (_04973_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _36606_ (_04974_, _04973_, _04971_);
  nand _36607_ (_04975_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _36608_ (_04976_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _36609_ (_04977_, _04976_, _04975_);
  and _36610_ (_04978_, _04977_, _04974_);
  nand _36611_ (_04979_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _36612_ (_04980_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _36613_ (_04981_, _04980_, _04979_);
  nand _36614_ (_04982_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand _36615_ (_04983_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _36616_ (_04984_, _04983_, _04982_);
  and _36617_ (_04985_, _04984_, _04981_);
  and _36618_ (_04986_, _04985_, _04978_);
  nand _36619_ (_04987_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand _36620_ (_04988_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _36621_ (_04989_, _04988_, _04987_);
  nand _36622_ (_04990_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _36623_ (_04991_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _36624_ (_04992_, _04991_, _04990_);
  and _36625_ (_04993_, _04992_, _04989_);
  nand _36626_ (_04994_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand _36627_ (_04995_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _36628_ (_04996_, _04995_, _04994_);
  nand _36629_ (_04997_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _36630_ (_04998_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _36631_ (_04999_, _04998_, _04997_);
  and _36632_ (_05000_, _04999_, _04996_);
  and _36633_ (_05001_, _05000_, _04993_);
  and _36634_ (_05002_, _05001_, _04986_);
  nand _36635_ (_05003_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand _36636_ (_05004_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _36637_ (_05006_, _05004_, _05003_);
  nand _36638_ (_05007_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _36639_ (_05008_, _00187_);
  nand _36640_ (_05009_, _04513_, _05008_);
  and _36641_ (_05010_, _05009_, _05007_);
  and _36642_ (_05011_, _05010_, _05006_);
  nand _36643_ (_05012_, _04565_, _04186_);
  nand _36644_ (_05013_, _04567_, _04131_);
  and _36645_ (_05014_, _05013_, _05012_);
  nand _36646_ (_05015_, _04570_, _03929_);
  nand _36647_ (_05016_, _04573_, _03982_);
  and _36648_ (_05017_, _05016_, _05015_);
  and _36649_ (_05018_, _05017_, _05014_);
  and _36650_ (_05020_, _05018_, _05011_);
  not _36651_ (_05021_, _04430_);
  or _36652_ (_05022_, _05021_, _03868_);
  nand _36653_ (_05023_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _36654_ (_05025_, _05023_, _05022_);
  and _36655_ (_05026_, _05025_, _05020_);
  and _36656_ (_05028_, _05026_, _05002_);
  nor _36657_ (_05030_, _05028_, _04441_);
  not _36658_ (_05031_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nor _36659_ (_05032_, _04521_, _05031_);
  or _36660_ (_05033_, _05032_, _04444_);
  or _36661_ (_05034_, _05033_, _05030_);
  or _36662_ (_05035_, _04523_, _26570_);
  and _36663_ (_05036_, _05035_, _22731_);
  and _36664_ (_27318_[0], _05036_, _05034_);
  not _36665_ (_05037_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nor _36666_ (_05038_, _04521_, _05037_);
  nand _36667_ (_05039_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _36668_ (_05040_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _36669_ (_05041_, _05040_, _05039_);
  nand _36670_ (_05042_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _36671_ (_05043_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _36672_ (_05044_, _05043_, _05042_);
  and _36673_ (_05045_, _05044_, _05041_);
  nand _36674_ (_05046_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _36675_ (_05047_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _36676_ (_05048_, _05047_, _05046_);
  nand _36677_ (_05049_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _36678_ (_05050_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _36679_ (_05051_, _05050_, _05049_);
  and _36680_ (_05053_, _05051_, _05048_);
  and _36681_ (_05054_, _05053_, _05045_);
  nand _36682_ (_05055_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand _36683_ (_05056_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _36684_ (_05057_, _05056_, _05055_);
  nand _36685_ (_05058_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nand _36686_ (_05059_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _36687_ (_05060_, _05059_, _05058_);
  and _36688_ (_05061_, _05060_, _05057_);
  nand _36689_ (_05062_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nand _36690_ (_05063_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _36691_ (_05065_, _05063_, _05062_);
  nand _36692_ (_05066_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _36693_ (_05067_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _36694_ (_05068_, _05067_, _05066_);
  and _36695_ (_05069_, _05068_, _05065_);
  and _36696_ (_05070_, _05069_, _05061_);
  and _36697_ (_05071_, _05070_, _05054_);
  nand _36698_ (_05072_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand _36699_ (_05073_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _36700_ (_05074_, _05073_, _05072_);
  nand _36701_ (_05075_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _36702_ (_05076_, _04513_, _00167_);
  and _36703_ (_05077_, _05076_, _05075_);
  and _36704_ (_05078_, _05077_, _05074_);
  nand _36705_ (_05079_, _04565_, _04216_);
  nand _36706_ (_05080_, _04567_, _04155_);
  and _36707_ (_05081_, _05080_, _05079_);
  nand _36708_ (_05082_, _04570_, _03954_);
  nand _36709_ (_05083_, _04573_, _04016_);
  and _36710_ (_05084_, _05083_, _05082_);
  and _36711_ (_05085_, _05084_, _05081_);
  and _36712_ (_05086_, _05085_, _05078_);
  nand _36713_ (_05087_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand _36714_ (_05088_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _36715_ (_05090_, _05088_, _05087_);
  and _36716_ (_05092_, _05090_, _05086_);
  and _36717_ (_05094_, _05092_, _05071_);
  nor _36718_ (_05095_, _05094_, _04441_);
  or _36719_ (_05096_, _05095_, _04444_);
  or _36720_ (_05097_, _05096_, _05038_);
  or _36721_ (_05098_, _04523_, _00393_);
  and _36722_ (_05099_, _05098_, _22731_);
  and _36723_ (_27318_[1], _05099_, _05097_);
  not _36724_ (_05100_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nor _36725_ (_05101_, _04521_, _05100_);
  nand _36726_ (_05102_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand _36727_ (_05103_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _36728_ (_05104_, _05103_, _05102_);
  nand _36729_ (_05105_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  nand _36730_ (_05106_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _36731_ (_05107_, _05106_, _05105_);
  and _36732_ (_05108_, _05107_, _05104_);
  nand _36733_ (_05109_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand _36734_ (_05110_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _36735_ (_05111_, _05110_, _05109_);
  nand _36736_ (_05112_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _36737_ (_05114_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _36738_ (_05115_, _05114_, _05112_);
  and _36739_ (_05117_, _05115_, _05111_);
  and _36740_ (_05118_, _05117_, _05108_);
  nand _36741_ (_05119_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _36742_ (_05120_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _36743_ (_05121_, _05120_, _05119_);
  nand _36744_ (_05122_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand _36745_ (_05123_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _36746_ (_05124_, _05123_, _05122_);
  and _36747_ (_05125_, _05124_, _05121_);
  nand _36748_ (_05126_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand _36749_ (_05127_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _36750_ (_05128_, _05127_, _05126_);
  nand _36751_ (_05129_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand _36752_ (_05130_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _36753_ (_05131_, _05130_, _05129_);
  and _36754_ (_05132_, _05131_, _05128_);
  and _36755_ (_05133_, _05132_, _05125_);
  and _36756_ (_05134_, _05133_, _05118_);
  nand _36757_ (_05136_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand _36758_ (_05137_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _36759_ (_05138_, _05137_, _05136_);
  nand _36760_ (_05139_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _36761_ (_05140_, _04513_, _00205_);
  and _36762_ (_05141_, _05140_, _05139_);
  and _36763_ (_05142_, _05141_, _05138_);
  nand _36764_ (_05144_, _04565_, _04227_);
  nand _36765_ (_05145_, _04567_, _04169_);
  and _36766_ (_05146_, _05145_, _05144_);
  nand _36767_ (_05147_, _04573_, _04027_);
  nand _36768_ (_05148_, _04570_, _03966_);
  and _36769_ (_05149_, _05148_, _05147_);
  and _36770_ (_05150_, _05149_, _05146_);
  and _36771_ (_05151_, _05150_, _05142_);
  nand _36772_ (_05152_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand _36773_ (_05153_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _36774_ (_05155_, _05153_, _05152_);
  and _36775_ (_05156_, _05155_, _05151_);
  and _36776_ (_05157_, _05156_, _05134_);
  or _36777_ (_05158_, _05157_, _04441_);
  nand _36778_ (_05159_, _05158_, _04523_);
  or _36779_ (_05160_, _05159_, _05101_);
  or _36780_ (_05161_, _04523_, _00473_);
  and _36781_ (_05162_, _05161_, _22731_);
  and _36782_ (_27318_[2], _05162_, _05160_);
  not _36783_ (_05164_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nor _36784_ (_05165_, _04521_, _05164_);
  nand _36785_ (_05167_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  nand _36786_ (_05169_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _36787_ (_05170_, _05169_, _05167_);
  nand _36788_ (_05171_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _36789_ (_05173_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _36790_ (_05174_, _05173_, _05171_);
  and _36791_ (_05176_, _05174_, _05170_);
  nand _36792_ (_05177_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand _36793_ (_05178_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _36794_ (_05179_, _05178_, _05177_);
  nand _36795_ (_05180_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _36796_ (_05181_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _36797_ (_05182_, _05181_, _05180_);
  and _36798_ (_05183_, _05182_, _05179_);
  and _36799_ (_05184_, _05183_, _05176_);
  nand _36800_ (_05185_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand _36801_ (_05186_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _36802_ (_05188_, _05186_, _05185_);
  nand _36803_ (_05190_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nand _36804_ (_05191_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _36805_ (_05192_, _05191_, _05190_);
  and _36806_ (_05193_, _05192_, _05188_);
  nand _36807_ (_05194_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand _36808_ (_05195_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _36809_ (_05196_, _05195_, _05194_);
  nand _36810_ (_05197_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand _36811_ (_05198_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _36812_ (_05199_, _05198_, _05197_);
  and _36813_ (_05200_, _05199_, _05196_);
  and _36814_ (_05201_, _05200_, _05193_);
  and _36815_ (_05202_, _05201_, _05184_);
  nand _36816_ (_05203_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nand _36817_ (_05204_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _36818_ (_05205_, _05204_, _05203_);
  nand _36819_ (_05207_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _36820_ (_05208_, _04513_, _26805_);
  and _36821_ (_05209_, _05208_, _05207_);
  and _36822_ (_05210_, _05209_, _05205_);
  nand _36823_ (_05211_, _04565_, _04202_);
  nand _36824_ (_05212_, _04567_, _04143_);
  and _36825_ (_05213_, _05212_, _05211_);
  nand _36826_ (_05214_, _04573_, _03997_);
  nand _36827_ (_05215_, _04570_, _03941_);
  and _36828_ (_05216_, _05215_, _05214_);
  and _36829_ (_05218_, _05216_, _05213_);
  and _36830_ (_05219_, _05218_, _05210_);
  nand _36831_ (_05221_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand _36832_ (_05223_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _36833_ (_05224_, _05223_, _05221_);
  and _36834_ (_05225_, _05224_, _05219_);
  and _36835_ (_05226_, _05225_, _05202_);
  or _36836_ (_05227_, _05226_, _04441_);
  nand _36837_ (_05228_, _05227_, _04523_);
  or _36838_ (_05229_, _05228_, _05165_);
  or _36839_ (_05230_, _04523_, _00569_);
  and _36840_ (_05231_, _05230_, _22731_);
  and _36841_ (_27318_[3], _05231_, _05229_);
  not _36842_ (_05232_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor _36843_ (_05233_, _04521_, _05232_);
  nand _36844_ (_05234_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  nand _36845_ (_05235_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _36846_ (_05236_, _05235_, _05234_);
  nand _36847_ (_05237_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand _36848_ (_05239_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _36849_ (_05240_, _05239_, _05237_);
  and _36850_ (_05242_, _05240_, _05236_);
  nand _36851_ (_05243_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _36852_ (_05244_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _36853_ (_05246_, _05244_, _05243_);
  nand _36854_ (_05247_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _36855_ (_05248_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _36856_ (_05249_, _05248_, _05247_);
  and _36857_ (_05250_, _05249_, _05246_);
  and _36858_ (_05251_, _05250_, _05242_);
  nand _36859_ (_05253_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _36860_ (_05254_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _36861_ (_05255_, _05254_, _05253_);
  nand _36862_ (_05256_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _36863_ (_05257_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _36864_ (_05258_, _05257_, _05256_);
  and _36865_ (_05259_, _05258_, _05255_);
  nand _36866_ (_05260_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand _36867_ (_05261_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _36868_ (_05262_, _05261_, _05260_);
  nand _36869_ (_05263_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _36870_ (_05264_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _36871_ (_05265_, _05264_, _05263_);
  and _36872_ (_05266_, _05265_, _05262_);
  and _36873_ (_05267_, _05266_, _05259_);
  and _36874_ (_05268_, _05267_, _05251_);
  nand _36875_ (_05269_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand _36876_ (_05270_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _36877_ (_05271_, _05270_, _05269_);
  nand _36878_ (_05273_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not _36879_ (_05274_, _00014_);
  nand _36880_ (_05275_, _04513_, _05274_);
  and _36881_ (_05276_, _05275_, _05273_);
  and _36882_ (_05277_, _05276_, _05271_);
  nand _36883_ (_05278_, _04565_, _04193_);
  nand _36884_ (_05279_, _04567_, _04136_);
  and _36885_ (_05280_, _05279_, _05278_);
  nand _36886_ (_05281_, _04573_, _03988_);
  nand _36887_ (_05282_, _04570_, _03934_);
  and _36888_ (_05284_, _05282_, _05281_);
  and _36889_ (_05285_, _05284_, _05280_);
  and _36890_ (_05286_, _05285_, _05277_);
  nand _36891_ (_05287_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand _36892_ (_05288_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _36893_ (_05289_, _05288_, _05287_);
  and _36894_ (_05291_, _05289_, _05286_);
  and _36895_ (_05292_, _05291_, _05268_);
  or _36896_ (_05293_, _05292_, _04441_);
  nand _36897_ (_05294_, _05293_, _04523_);
  or _36898_ (_05295_, _05294_, _05233_);
  or _36899_ (_05296_, _04523_, _00654_);
  and _36900_ (_05297_, _05296_, _22731_);
  and _36901_ (_27318_[4], _05297_, _05295_);
  not _36902_ (_05298_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _36903_ (_05299_, _04426_, _05298_);
  and _36904_ (_05300_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _36905_ (_05301_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _36906_ (_05302_, _05301_, _05300_);
  and _36907_ (_05304_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _36908_ (_05305_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _36909_ (_05306_, _05305_, _05304_);
  or _36910_ (_05307_, _05306_, _05302_);
  and _36911_ (_05308_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _36912_ (_05309_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _36913_ (_05310_, _05309_, _05308_);
  and _36914_ (_05311_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _36915_ (_05312_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _36916_ (_05313_, _05312_, _05311_);
  or _36917_ (_05314_, _05313_, _05310_);
  or _36918_ (_05315_, _05314_, _05307_);
  and _36919_ (_05316_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _36920_ (_05317_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _36921_ (_05318_, _05317_, _05316_);
  and _36922_ (_05319_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _36923_ (_05321_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _36924_ (_05322_, _05321_, _05319_);
  or _36925_ (_05323_, _05322_, _05318_);
  and _36926_ (_05324_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _36927_ (_05326_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _36928_ (_05327_, _05326_, _05324_);
  and _36929_ (_05328_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _36930_ (_05329_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _36931_ (_05331_, _05329_, _05328_);
  or _36932_ (_05332_, _05331_, _05327_);
  or _36933_ (_05333_, _05332_, _05323_);
  or _36934_ (_05334_, _05333_, _05315_);
  and _36935_ (_05335_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _36936_ (_05337_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _36937_ (_05338_, _05337_, _05335_);
  and _36938_ (_05339_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not _36939_ (_05340_, _00046_);
  and _36940_ (_05341_, _04513_, _05340_);
  or _36941_ (_05342_, _05341_, _05339_);
  or _36942_ (_05343_, _05342_, _05338_);
  and _36943_ (_05344_, _04565_, _04221_);
  and _36944_ (_05345_, _04567_, _04160_);
  or _36945_ (_05347_, _05345_, _05344_);
  and _36946_ (_05348_, _04570_, _03959_);
  and _36947_ (_05349_, _04573_, _04020_);
  or _36948_ (_05350_, _05349_, _05348_);
  or _36949_ (_05351_, _05350_, _05347_);
  or _36950_ (_05352_, _05351_, _05343_);
  and _36951_ (_05353_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _36952_ (_05355_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _36953_ (_05356_, _05355_, _05353_);
  or _36954_ (_05358_, _05356_, _05352_);
  nor _36955_ (_05359_, _05358_, _05334_);
  nor _36956_ (_05360_, _05359_, _04440_);
  nor _36957_ (_05361_, _04521_, _05298_);
  or _36958_ (_05362_, _05361_, _05360_);
  and _36959_ (_05363_, _05362_, _05299_);
  or _36960_ (_05364_, _05363_, _04444_);
  or _36961_ (_05365_, _04523_, _00747_);
  and _36962_ (_05366_, _05365_, _22731_);
  and _36963_ (_27318_[5], _05366_, _05364_);
  not _36964_ (_05367_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor _36965_ (_05368_, _04521_, _05367_);
  nand _36966_ (_05370_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand _36967_ (_05371_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _36968_ (_05372_, _05371_, _05370_);
  nand _36969_ (_05373_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand _36970_ (_05374_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _36971_ (_05375_, _05374_, _05373_);
  and _36972_ (_05376_, _05375_, _05372_);
  nand _36973_ (_05377_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _36974_ (_05378_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _36975_ (_05380_, _05378_, _05377_);
  nand _36976_ (_05381_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand _36977_ (_05382_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _36978_ (_05384_, _05382_, _05381_);
  and _36979_ (_05385_, _05384_, _05380_);
  and _36980_ (_05386_, _05385_, _05376_);
  nand _36981_ (_05387_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand _36982_ (_05388_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _36983_ (_05389_, _05388_, _05387_);
  nand _36984_ (_05391_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  nand _36985_ (_05392_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _36986_ (_05393_, _05392_, _05391_);
  and _36987_ (_05394_, _05393_, _05389_);
  nand _36988_ (_05395_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _36989_ (_05396_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _36990_ (_05397_, _05396_, _05395_);
  nand _36991_ (_05398_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _36992_ (_05399_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _36993_ (_05400_, _05399_, _05398_);
  and _36994_ (_05401_, _05400_, _05397_);
  and _36995_ (_05402_, _05401_, _05394_);
  and _36996_ (_05403_, _05402_, _05386_);
  nand _36997_ (_05404_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand _36998_ (_05405_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _36999_ (_05406_, _05405_, _05404_);
  nand _37000_ (_05407_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not _37001_ (_05408_, _00084_);
  nand _37002_ (_05409_, _04513_, _05408_);
  and _37003_ (_05410_, _05409_, _05407_);
  and _37004_ (_05411_, _05410_, _05406_);
  nand _37005_ (_05412_, _04565_, _04232_);
  nand _37006_ (_05413_, _04567_, _04175_);
  and _37007_ (_05414_, _05413_, _05412_);
  nand _37008_ (_05415_, _04570_, _03972_);
  nand _37009_ (_05416_, _04573_, _04031_);
  and _37010_ (_05417_, _05416_, _05415_);
  and _37011_ (_05418_, _05417_, _05414_);
  and _37012_ (_05419_, _05418_, _05411_);
  nand _37013_ (_05420_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _37014_ (_05421_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _37015_ (_05422_, _05421_, _05420_);
  and _37016_ (_05424_, _05422_, _05419_);
  and _37017_ (_05425_, _05424_, _05403_);
  or _37018_ (_05426_, _05425_, _04441_);
  nand _37019_ (_05427_, _05426_, _04523_);
  or _37020_ (_05428_, _05427_, _05368_);
  nand _37021_ (_05429_, _04444_, _00813_);
  and _37022_ (_05430_, _05429_, _22731_);
  and _37023_ (_27318_[6], _05430_, _05428_);
  and _37024_ (_05431_, _24474_, _24408_);
  and _37025_ (_05432_, _05431_, _23583_);
  not _37026_ (_05434_, _05431_);
  and _37027_ (_05435_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or _37028_ (_26604_, _05435_, _05432_);
  and _37029_ (_05436_, _05431_, _23548_);
  and _37030_ (_05437_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or _37031_ (_26621_, _05437_, _05436_);
  and _37032_ (_05438_, _24476_, _24349_);
  and _37033_ (_05439_, _05438_, _24219_);
  not _37034_ (_05440_, _05438_);
  and _37035_ (_05441_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _37036_ (_27185_, _05441_, _05439_);
  and _37037_ (_05442_, _24476_, _24159_);
  and _37038_ (_05443_, _05442_, _23548_);
  not _37039_ (_05444_, _05442_);
  and _37040_ (_05446_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _37041_ (_26661_, _05446_, _05443_);
  and _37042_ (_05448_, _02502_, _23583_);
  and _37043_ (_05449_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or _37044_ (_26685_, _05449_, _05448_);
  and _37045_ (_05451_, _02502_, _24089_);
  and _37046_ (_05453_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _37047_ (_26725_, _05453_, _05451_);
  and _37048_ (_05454_, _02502_, _23887_);
  and _37049_ (_05455_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or _37050_ (_26728_, _05455_, _05454_);
  and _37051_ (_05456_, _24408_, _24056_);
  and _37052_ (_05457_, _05456_, _24134_);
  not _37053_ (_05458_, _05456_);
  and _37054_ (_05459_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _37055_ (_26746_, _05459_, _05457_);
  and _37056_ (_05460_, _24140_, _24006_);
  and _37057_ (_05461_, _05460_, _24219_);
  not _37058_ (_05462_, _05460_);
  and _37059_ (_05464_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or _37060_ (_26771_, _05464_, _05461_);
  and _37061_ (_05465_, _24297_, _23945_);
  and _37062_ (_05467_, _05465_, _23887_);
  not _37063_ (_05468_, _05465_);
  and _37064_ (_05469_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or _37065_ (_26774_, _05469_, _05467_);
  and _37066_ (_05471_, _05456_, _24089_);
  and _37067_ (_05472_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _37068_ (_27126_, _05472_, _05471_);
  and _37069_ (_05473_, _05456_, _23887_);
  and _37070_ (_05475_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _37071_ (_26785_, _05475_, _05473_);
  and _37072_ (_05478_, _24496_, _24349_);
  and _37073_ (_05479_, _05478_, _24051_);
  not _37074_ (_05480_, _05478_);
  and _37075_ (_05481_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or _37076_ (_26817_, _05481_, _05479_);
  and _37077_ (_05482_, _05456_, _24219_);
  and _37078_ (_05484_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _37079_ (_00007_, _05484_, _05482_);
  and _37080_ (_05485_, _24899_, _24408_);
  and _37081_ (_05486_, _05485_, _24051_);
  not _37082_ (_05487_, _05485_);
  and _37083_ (_05488_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _37084_ (_00019_, _05488_, _05486_);
  and _37085_ (_05489_, _05478_, _24134_);
  and _37086_ (_05490_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or _37087_ (_00022_, _05490_, _05489_);
  and _37088_ (_05491_, _24408_, _24223_);
  and _37089_ (_05492_, _05491_, _23996_);
  not _37090_ (_05493_, _05491_);
  and _37091_ (_05494_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or _37092_ (_00032_, _05494_, _05492_);
  and _37093_ (_05495_, _05460_, _23548_);
  and _37094_ (_05496_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _37095_ (_00044_, _05496_, _05495_);
  and _37096_ (_05497_, _02045_, _23548_);
  and _37097_ (_05498_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _37098_ (_00074_, _05498_, _05497_);
  and _37099_ (_05499_, _05460_, _23887_);
  and _37100_ (_05500_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _37101_ (_00079_, _05500_, _05499_);
  and _37102_ (_05501_, _05478_, _23996_);
  and _37103_ (_05502_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or _37104_ (_00082_, _05502_, _05501_);
  and _37105_ (_05504_, _05491_, _24089_);
  and _37106_ (_05505_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or _37107_ (_00087_, _05505_, _05504_);
  and _37108_ (_05506_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and _37109_ (_05507_, _04937_, _23996_);
  or _37110_ (_00103_, _05507_, _05506_);
  and _37111_ (_05508_, _05465_, _24219_);
  and _37112_ (_05509_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or _37113_ (_00172_, _05509_, _05508_);
  or _37114_ (_05510_, _03083_, _00143_);
  or _37115_ (_05511_, _05510_, _26816_);
  not _37116_ (_05512_, _03083_);
  or _37117_ (_05513_, _05512_, _00191_);
  nand _37118_ (_05514_, _05513_, _05511_);
  and _37119_ (_05515_, _05514_, _22888_);
  nor _37120_ (_05516_, _05514_, _22888_);
  nor _37121_ (_05517_, _05516_, _05515_);
  and _37122_ (_05518_, _05510_, _03700_);
  nor _37123_ (_05519_, _05518_, _24096_);
  and _37124_ (_05520_, _05510_, _00051_);
  nor _37125_ (_05521_, _05520_, _24001_);
  nor _37126_ (_05522_, _05521_, _05519_);
  nor _37127_ (_05523_, _22968_, _22871_);
  not _37128_ (_05524_, _05523_);
  not _37129_ (_05525_, _05510_);
  nor _37130_ (_05526_, _05525_, _00090_);
  nor _37131_ (_05527_, _05526_, _05524_);
  and _37132_ (_05528_, _05526_, _05524_);
  nor _37133_ (_05529_, _05528_, _05527_);
  and _37134_ (_05530_, _05529_, _05522_);
  and _37135_ (_05531_, _05530_, _05517_);
  not _37136_ (_05532_, _22953_);
  nor _37137_ (_05533_, _05510_, _00051_);
  nor _37138_ (_05534_, _05512_, _00228_);
  nor _37139_ (_05535_, _05534_, _05533_);
  nor _37140_ (_05536_, _05535_, _05532_);
  and _37141_ (_05537_, _05535_, _05532_);
  nor _37142_ (_05538_, _05537_, _05536_);
  not _37143_ (_05539_, _05538_);
  and _37144_ (_05540_, _05510_, _26816_);
  and _37145_ (_05541_, _05525_, _00090_);
  nor _37146_ (_05542_, _05541_, _05540_);
  and _37147_ (_05543_, _05542_, _22972_);
  nor _37148_ (_05544_, _05542_, _22972_);
  or _37149_ (_05545_, _05544_, _05543_);
  nor _37150_ (_05546_, _05545_, _05539_);
  or _37151_ (_05547_, _05510_, _00027_);
  or _37152_ (_05548_, _05512_, _00171_);
  nand _37153_ (_05549_, _05548_, _05547_);
  and _37154_ (_05550_, _05549_, _22921_);
  nor _37155_ (_05551_, _05549_, _22921_);
  nor _37156_ (_05552_, _05551_, _05550_);
  and _37157_ (_05553_, _05520_, _24001_);
  not _37158_ (_05554_, _05553_);
  and _37159_ (_05555_, _05518_, _24096_);
  not _37160_ (_05556_, _05555_);
  nor _37161_ (_05558_, _00146_, _22849_);
  and _37162_ (_05559_, _05558_, _05556_);
  and _37163_ (_05560_, _05559_, _05554_);
  and _37164_ (_05561_, _05560_, _05552_);
  and _37165_ (_05562_, _05561_, _05546_);
  and _37166_ (_05563_, _05562_, _05531_);
  and _37167_ (_26890_, _05563_, _22731_);
  and _37168_ (_26891_[7], _23995_, _22731_);
  nor _37169_ (_26893_[2], _00228_, rst);
  and _37170_ (_05565_, _04865_, _24051_);
  and _37171_ (_05566_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or _37172_ (_00184_, _05566_, _05565_);
  and _37173_ (_05567_, _02039_, _22974_);
  not _37174_ (_05568_, _05567_);
  and _37175_ (_05569_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  and _37176_ (_05570_, _05567_, _23548_);
  or _37177_ (_00203_, _05570_, _05569_);
  and _37178_ (_05571_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and _37179_ (_05572_, _05567_, _23583_);
  or _37180_ (_00209_, _05572_, _05571_);
  and _37181_ (_05573_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  and _37182_ (_05574_, _05567_, _24051_);
  or _37183_ (_00212_, _05574_, _05573_);
  and _37184_ (_05576_, _03281_, _23996_);
  and _37185_ (_05577_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or _37186_ (_00215_, _05577_, _05576_);
  and _37187_ (_05578_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and _37188_ (_05579_, _05567_, _24134_);
  or _37189_ (_00262_, _05579_, _05578_);
  and _37190_ (_05580_, _02039_, _24223_);
  not _37191_ (_05582_, _05580_);
  and _37192_ (_05583_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _37193_ (_05584_, _05580_, _23548_);
  or _37194_ (_00270_, _05584_, _05583_);
  and _37195_ (_05585_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _37196_ (_05587_, _05580_, _23583_);
  or _37197_ (_00276_, _05587_, _05585_);
  and _37198_ (_05589_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _37199_ (_05591_, _05580_, _24051_);
  or _37200_ (_00280_, _05591_, _05589_);
  and _37201_ (_05592_, _04920_, _23996_);
  and _37202_ (_05593_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _37203_ (_00289_, _05593_, _05592_);
  and _37204_ (_05594_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _37205_ (_05595_, _05580_, _24134_);
  or _37206_ (_00291_, _05595_, _05594_);
  and _37207_ (_05596_, _02039_, _24056_);
  not _37208_ (_05597_, _05596_);
  and _37209_ (_05598_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and _37210_ (_05599_, _05596_, _24219_);
  or _37211_ (_00299_, _05599_, _05598_);
  and _37212_ (_05600_, _03275_, _23887_);
  and _37213_ (_05601_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or _37214_ (_00302_, _05601_, _05600_);
  and _37215_ (_05603_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and _37216_ (_05604_, _05596_, _23887_);
  or _37217_ (_00305_, _05604_, _05603_);
  and _37218_ (_05605_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and _37219_ (_05606_, _05596_, _24089_);
  or _37220_ (_00310_, _05606_, _05605_);
  and _37221_ (_26891_[0], _24218_, _22731_);
  and _37222_ (_26891_[1], _23547_, _22731_);
  and _37223_ (_26891_[2], _23886_, _22731_);
  and _37224_ (_26891_[3], _23582_, _22731_);
  and _37225_ (_26891_[4], _24088_, _22731_);
  and _37226_ (_26891_[5], _24050_, _22731_);
  and _37227_ (_26891_[6], _24133_, _22731_);
  nor _37228_ (_26893_[0], _00191_, rst);
  nor _37229_ (_26893_[1], _00171_, rst);
  and _37230_ (_05609_, _05491_, _23548_);
  and _37231_ (_05610_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or _37232_ (_00515_, _05610_, _05609_);
  nor _37233_ (_05611_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _37234_ (_05612_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01836_);
  nor _37235_ (_05613_, _05612_, _05611_);
  not _37236_ (_05614_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _37237_ (_05615_, _00613_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _37238_ (_05616_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01836_);
  nor _37239_ (_05617_, _05616_, _05615_);
  nor _37240_ (_05618_, _05617_, _05614_);
  and _37241_ (_05619_, _05617_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _37242_ (_05620_, _05619_, _05618_);
  not _37243_ (_05621_, _05620_);
  nor _37244_ (_05622_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _37245_ (_05623_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01836_);
  nor _37246_ (_05624_, _05623_, _05622_);
  not _37247_ (_05625_, _05624_);
  nor _37248_ (_05626_, _00517_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _37249_ (_05627_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01836_);
  nor _37250_ (_05628_, _05627_, _05626_);
  and _37251_ (_05629_, _05628_, _05625_);
  nand _37252_ (_05630_, _05629_, _05621_);
  and _37253_ (_05631_, _05630_, _05613_);
  nor _37254_ (_05632_, _05628_, _05625_);
  not _37255_ (_05633_, _05632_);
  not _37256_ (_05634_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _37257_ (_05635_, _05617_, _05634_);
  and _37258_ (_05636_, _05617_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _37259_ (_05637_, _05636_, _05635_);
  nor _37260_ (_05638_, _05637_, _05633_);
  and _37261_ (_05639_, _05628_, _05624_);
  not _37262_ (_05640_, _05639_);
  not _37263_ (_05641_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _37264_ (_05642_, _05617_, _05641_);
  and _37265_ (_05643_, _05617_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _37266_ (_05645_, _05643_, _05642_);
  nor _37267_ (_05646_, _05645_, _05640_);
  nor _37268_ (_05647_, _05646_, _05638_);
  nor _37269_ (_05649_, _05628_, _05624_);
  not _37270_ (_05651_, _05649_);
  and _37271_ (_05652_, _05617_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not _37272_ (_05653_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _37273_ (_05654_, _05617_, _05653_);
  nor _37274_ (_05655_, _05654_, _05652_);
  or _37275_ (_05656_, _05655_, _05651_);
  and _37276_ (_05657_, _05656_, _05647_);
  and _37277_ (_05658_, _05657_, _05631_);
  not _37278_ (_05659_, _05628_);
  not _37279_ (_05660_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _37280_ (_05661_, _05617_, _05660_);
  and _37281_ (_05662_, _05617_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _37282_ (_05663_, _05662_, _05661_);
  nor _37283_ (_05664_, _05663_, _05659_);
  not _37284_ (_05665_, _05664_);
  nor _37285_ (_05667_, _05628_, _05617_);
  and _37286_ (_05668_, _05667_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _37287_ (_05669_, _05659_, _05617_);
  and _37288_ (_05670_, _05669_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _37289_ (_05671_, _05670_, _05668_);
  and _37290_ (_05672_, _05671_, _05665_);
  nor _37291_ (_05673_, _05672_, _05624_);
  and _37292_ (_05674_, _05667_, _05624_);
  and _37293_ (_05675_, _05674_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _37294_ (_05677_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _37295_ (_05678_, _05617_, _05677_);
  nor _37296_ (_05679_, _05617_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _37297_ (_05680_, _05679_, _05678_);
  nor _37298_ (_05681_, _05680_, _05640_);
  and _37299_ (_05682_, _05617_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _37300_ (_05683_, _05682_, _05632_);
  or _37301_ (_05684_, _05683_, _05613_);
  or _37302_ (_05685_, _05684_, _05681_);
  or _37303_ (_05686_, _05685_, _05675_);
  nor _37304_ (_05687_, _05686_, _05673_);
  nor _37305_ (_05688_, _05687_, _05658_);
  not _37306_ (_05689_, _05688_);
  and _37307_ (_05690_, _05689_, word_in[7]);
  not _37308_ (_05691_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _37309_ (_05692_, _05613_, _05691_);
  or _37310_ (_05693_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _37311_ (_05694_, _05693_, _05692_);
  and _37312_ (_05696_, _05694_, _05639_);
  not _37313_ (_05697_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _37314_ (_05698_, _05613_, _05697_);
  or _37315_ (_05699_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _37316_ (_05700_, _05699_, _05698_);
  and _37317_ (_05701_, _05700_, _05632_);
  or _37318_ (_05702_, _05701_, _05696_);
  not _37319_ (_05704_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _37320_ (_05705_, _05613_, _05704_);
  or _37321_ (_05706_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _37322_ (_05707_, _05706_, _05705_);
  and _37323_ (_05708_, _05707_, _05629_);
  not _37324_ (_05709_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _37325_ (_05710_, _05613_, _05709_);
  or _37326_ (_05711_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _37327_ (_05712_, _05711_, _05710_);
  and _37328_ (_05713_, _05712_, _05649_);
  or _37329_ (_05715_, _05713_, _05708_);
  or _37330_ (_05716_, _05715_, _05702_);
  and _37331_ (_05717_, _05716_, _05617_);
  not _37332_ (_05719_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _37333_ (_05720_, _05613_, _05719_);
  or _37334_ (_05721_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _37335_ (_05722_, _05721_, _05720_);
  and _37336_ (_05723_, _05722_, _05674_);
  not _37337_ (_05724_, _05617_);
  and _37338_ (_05725_, _05639_, _05724_);
  not _37339_ (_05726_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _37340_ (_05727_, _05613_, _05726_);
  or _37341_ (_05728_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _37342_ (_05730_, _05728_, _05727_);
  and _37343_ (_05731_, _05730_, _05725_);
  not _37344_ (_05732_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _37345_ (_05733_, _05613_, _05732_);
  or _37346_ (_05734_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _37347_ (_05735_, _05734_, _05733_);
  and _37348_ (_05736_, _05735_, _05629_);
  not _37349_ (_05737_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _37350_ (_05738_, _05613_, _05737_);
  or _37351_ (_05739_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _37352_ (_05741_, _05739_, _05738_);
  and _37353_ (_05742_, _05741_, _05649_);
  or _37354_ (_05743_, _05742_, _05736_);
  and _37355_ (_05744_, _05743_, _05724_);
  or _37356_ (_05745_, _05744_, _05731_);
  or _37357_ (_05746_, _05745_, _05723_);
  or _37358_ (_05747_, _05746_, _05717_);
  and _37359_ (_05748_, _05747_, _05688_);
  or _37360_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _05748_, _05690_);
  and _37361_ (_05749_, _03275_, _24134_);
  and _37362_ (_05750_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _37363_ (_00527_, _05750_, _05749_);
  and _37364_ (_05751_, _05625_, _05613_);
  not _37365_ (_05752_, _05751_);
  and _37366_ (_05753_, _05624_, _05613_);
  and _37367_ (_05754_, _05753_, _05628_);
  nor _37368_ (_05755_, _05753_, _05628_);
  nor _37369_ (_05756_, _05755_, _05754_);
  not _37370_ (_05757_, _05756_);
  nor _37371_ (_05758_, _05757_, _05680_);
  nor _37372_ (_05759_, _05754_, _05724_);
  nor _37373_ (_05760_, _05659_, _05617_);
  and _37374_ (_05761_, _05760_, _05753_);
  nor _37375_ (_05762_, _05761_, _05759_);
  nor _37376_ (_05763_, _05762_, _05756_);
  and _37377_ (_05765_, _05763_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _37378_ (_05766_, _05755_, _05617_);
  nor _37379_ (_05767_, _05766_, _05759_);
  and _37380_ (_05768_, _05767_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _37381_ (_05769_, _05768_, _05765_);
  nor _37382_ (_05770_, _05769_, _05758_);
  nor _37383_ (_05771_, _05770_, _05752_);
  not _37384_ (_05772_, _05753_);
  nor _37385_ (_05773_, _05757_, _05663_);
  and _37386_ (_05774_, _05767_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _37387_ (_05775_, _05774_, _05773_);
  or _37388_ (_05776_, _05775_, _05772_);
  nand _37389_ (_05777_, _05761_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _37390_ (_05779_, _05777_, _05776_);
  not _37391_ (_05780_, _05779_);
  nor _37392_ (_05782_, _05780_, _05771_);
  nor _37393_ (_05784_, _05624_, _05613_);
  or _37394_ (_05785_, _05753_, _05784_);
  not _37395_ (_05787_, _05785_);
  nor _37396_ (_05789_, _05757_, _05620_);
  and _37397_ (_05790_, _05763_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _37398_ (_05792_, _05767_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _37399_ (_05793_, _05792_, _05790_);
  nor _37400_ (_05795_, _05793_, _05789_);
  or _37401_ (_05796_, _05795_, _05787_);
  and _37402_ (_05797_, _05756_, _05724_);
  and _37403_ (_05798_, _05797_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _37404_ (_05799_, _05763_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _37405_ (_05800_, _05756_, _05617_);
  and _37406_ (_05801_, _05800_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _37407_ (_05802_, _05767_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _37408_ (_05803_, _05802_, _05801_);
  or _37409_ (_05804_, _05803_, _05799_);
  nor _37410_ (_05806_, _05804_, _05798_);
  or _37411_ (_05807_, _05806_, _05785_);
  and _37412_ (_05808_, _05807_, _05796_);
  or _37413_ (_05809_, _05808_, _05613_);
  and _37414_ (_05810_, _05809_, _05782_);
  not _37415_ (_05811_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _37416_ (_05813_, _05613_, _05811_);
  or _37417_ (_05814_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _37418_ (_05815_, _05814_, _05813_);
  and _37419_ (_05817_, _05815_, _05787_);
  not _37420_ (_05818_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _37421_ (_05819_, _05613_, _05818_);
  or _37422_ (_05821_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _37423_ (_05822_, _05821_, _05819_);
  and _37424_ (_05823_, _05822_, _05785_);
  or _37425_ (_05824_, _05823_, _05817_);
  and _37426_ (_05826_, _05824_, _05800_);
  not _37427_ (_05827_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _37428_ (_05828_, _05613_, _05827_);
  or _37429_ (_05829_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _37430_ (_05830_, _05829_, _05828_);
  and _37431_ (_05831_, _05830_, _05787_);
  not _37432_ (_05832_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _37433_ (_05834_, _05613_, _05832_);
  or _37434_ (_05835_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _37435_ (_05836_, _05835_, _05834_);
  and _37436_ (_05837_, _05836_, _05785_);
  or _37437_ (_05838_, _05837_, _05831_);
  and _37438_ (_05839_, _05838_, _05763_);
  or _37439_ (_05841_, _05839_, _05826_);
  not _37440_ (_05842_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _37441_ (_05844_, _05613_, _05842_);
  or _37442_ (_05845_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _37443_ (_05846_, _05845_, _05844_);
  and _37444_ (_05847_, _05846_, _05785_);
  not _37445_ (_05848_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _37446_ (_05849_, _05613_, _05848_);
  or _37447_ (_05850_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _37448_ (_05851_, _05850_, _05849_);
  and _37449_ (_05852_, _05851_, _05787_);
  or _37450_ (_05853_, _05852_, _05847_);
  and _37451_ (_05854_, _05853_, _05767_);
  not _37452_ (_05855_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _37453_ (_05856_, _05613_, _05855_);
  or _37454_ (_05857_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _37455_ (_05858_, _05857_, _05856_);
  and _37456_ (_05860_, _05858_, _05785_);
  not _37457_ (_05862_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _37458_ (_05863_, _05613_, _05862_);
  or _37459_ (_05864_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _37460_ (_05865_, _05864_, _05863_);
  and _37461_ (_05867_, _05865_, _05787_);
  or _37462_ (_05868_, _05867_, _05860_);
  and _37463_ (_05869_, _05868_, _05797_);
  or _37464_ (_05870_, _05869_, _05854_);
  nor _37465_ (_05871_, _05870_, _05841_);
  nor _37466_ (_05872_, _05871_, _05810_);
  and _37467_ (_05873_, _05810_, word_in[15]);
  or _37468_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _05873_, _05872_);
  and _37469_ (_05874_, _05639_, _05617_);
  and _37470_ (_05875_, _05649_, _05724_);
  or _37471_ (_05876_, _05875_, _05874_);
  and _37472_ (_05877_, _05876_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _37473_ (_05878_, _05877_);
  nor _37474_ (_05879_, _05639_, _05649_);
  not _37475_ (_05880_, _05879_);
  nor _37476_ (_05881_, _05880_, _05620_);
  or _37477_ (_05883_, _05639_, _05617_);
  or _37478_ (_05884_, _05649_, _05724_);
  and _37479_ (_05885_, _05884_, _05883_);
  and _37480_ (_05886_, _05885_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _37481_ (_05887_, _05886_, _05881_);
  and _37482_ (_05888_, _05887_, _05878_);
  nor _37483_ (_05889_, _05888_, _05772_);
  nor _37484_ (_05890_, _05880_, _05645_);
  and _37485_ (_05891_, _05876_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _37486_ (_05893_, _05885_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _37487_ (_05894_, _05893_, _05891_);
  nor _37488_ (_05895_, _05894_, _05890_);
  nor _37489_ (_05896_, _05895_, _05752_);
  nor _37490_ (_05897_, _05896_, _05889_);
  not _37491_ (_05898_, _05784_);
  nor _37492_ (_05899_, _05880_, _05680_);
  and _37493_ (_05900_, _05876_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _37494_ (_05901_, _05885_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _37495_ (_05902_, _05901_, _05900_);
  nor _37496_ (_05903_, _05902_, _05899_);
  nor _37497_ (_05904_, _05903_, _05898_);
  not _37498_ (_05905_, _05613_);
  and _37499_ (_05906_, _05624_, _05905_);
  not _37500_ (_05907_, _05906_);
  nor _37501_ (_05908_, _05880_, _05663_);
  and _37502_ (_05910_, _05876_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _37503_ (_05911_, _05885_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _37504_ (_05912_, _05911_, _05910_);
  nor _37505_ (_05914_, _05912_, _05908_);
  nor _37506_ (_05915_, _05914_, _05907_);
  nor _37507_ (_05916_, _05915_, _05904_);
  and _37508_ (_05918_, _05916_, _05897_);
  and _37509_ (_05919_, _05918_, word_in[23]);
  and _37510_ (_05920_, _05640_, _05617_);
  or _37511_ (_05921_, _05920_, _05725_);
  and _37512_ (_05922_, _05730_, _05629_);
  and _37513_ (_05923_, _05722_, _05649_);
  or _37514_ (_05924_, _05923_, _05922_);
  and _37515_ (_05925_, _05735_, _05632_);
  and _37516_ (_05926_, _05741_, _05639_);
  or _37517_ (_05927_, _05926_, _05925_);
  or _37518_ (_05929_, _05927_, _05924_);
  or _37519_ (_05930_, _05929_, _05921_);
  and _37520_ (_05931_, _05707_, _05632_);
  and _37521_ (_05933_, _05700_, _05649_);
  or _37522_ (_05934_, _05933_, _05931_);
  and _37523_ (_05936_, _05694_, _05629_);
  and _37524_ (_05937_, _05712_, _05639_);
  or _37525_ (_05938_, _05937_, _05936_);
  nor _37526_ (_05939_, _05938_, _05934_);
  nand _37527_ (_05941_, _05939_, _05921_);
  nand _37528_ (_05942_, _05941_, _05930_);
  nor _37529_ (_05943_, _05942_, _05918_);
  or _37530_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _05943_, _05919_);
  and _37531_ (_05944_, _03269_, _24089_);
  and _37532_ (_05946_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or _37533_ (_00541_, _05946_, _05944_);
  and _37534_ (_05947_, _05898_, _05628_);
  nor _37535_ (_05948_, _05898_, _05628_);
  nor _37536_ (_05949_, _05948_, _05947_);
  not _37537_ (_05950_, _05949_);
  or _37538_ (_05952_, _05950_, _05663_);
  and _37539_ (_05953_, _05947_, _05617_);
  nor _37540_ (_05955_, _05947_, _05617_);
  nor _37541_ (_05956_, _05955_, _05953_);
  and _37542_ (_05957_, _05956_, _05950_);
  nand _37543_ (_05958_, _05957_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _37544_ (_05959_, _05958_, _05952_);
  or _37545_ (_05961_, _05959_, _05752_);
  and _37546_ (_05962_, _05628_, _05617_);
  and _37547_ (_05963_, _05751_, _05962_);
  and _37548_ (_05964_, _05963_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _37549_ (_05965_, _05754_, _05617_);
  and _37550_ (_05966_, _05965_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _37551_ (_05967_, _05680_, _05950_);
  and _37552_ (_05968_, _05957_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _37553_ (_05969_, _05968_, _05967_);
  and _37554_ (_05970_, _05969_, _05753_);
  or _37555_ (_05971_, _05970_, _05966_);
  nor _37556_ (_05972_, _05971_, _05964_);
  and _37557_ (_05973_, _05972_, _05961_);
  or _37558_ (_05975_, _05950_, _05620_);
  nand _37559_ (_05976_, _05957_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _37560_ (_05977_, _05976_, _05975_);
  or _37561_ (_05979_, _05977_, _05907_);
  and _37562_ (_05980_, _05948_, _05635_);
  and _37563_ (_05982_, _05874_, _05905_);
  and _37564_ (_05983_, _05982_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _37565_ (_05984_, _05950_, _05645_);
  and _37566_ (_05985_, _05957_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _37567_ (_05986_, _05985_, _05984_);
  and _37568_ (_05987_, _05986_, _05784_);
  or _37569_ (_05988_, _05987_, _05983_);
  nor _37570_ (_05989_, _05988_, _05980_);
  and _37571_ (_05990_, _05989_, _05979_);
  and _37572_ (_05991_, _05990_, _05973_);
  and _37573_ (_05992_, _05836_, _05787_);
  and _37574_ (_05993_, _05830_, _05785_);
  or _37575_ (_05994_, _05993_, _05992_);
  and _37576_ (_05995_, _05994_, _05957_);
  nor _37577_ (_05996_, _05956_, _05949_);
  and _37578_ (_05997_, _05846_, _05787_);
  and _37579_ (_05999_, _05851_, _05785_);
  or _37580_ (_06000_, _05999_, _05997_);
  and _37581_ (_06001_, _06000_, _05996_);
  not _37582_ (_06002_, _05948_);
  and _37583_ (_06003_, _05955_, _06002_);
  and _37584_ (_06004_, _05858_, _05787_);
  and _37585_ (_06005_, _05865_, _05785_);
  or _37586_ (_06006_, _06005_, _06004_);
  and _37587_ (_06007_, _06006_, _06003_);
  and _37588_ (_06008_, _05949_, _05617_);
  and _37589_ (_06009_, _05822_, _05787_);
  and _37590_ (_06010_, _05815_, _05785_);
  or _37591_ (_06011_, _06010_, _06009_);
  and _37592_ (_06012_, _06011_, _06008_);
  or _37593_ (_06013_, _06012_, _06007_);
  or _37594_ (_06014_, _06013_, _06001_);
  nor _37595_ (_06015_, _06014_, _05995_);
  nor _37596_ (_06016_, _06015_, _05991_);
  and _37597_ (_06017_, _05991_, word_in[31]);
  or _37598_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _06017_, _06016_);
  or _37599_ (_06018_, _05962_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _37600_ (_26822_[15], _06018_, _22731_);
  and _37601_ (_06019_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and _37602_ (_06020_, _05596_, _24051_);
  or _37603_ (_00596_, _06020_, _06019_);
  and _37604_ (_06022_, _05918_, _22731_);
  and _37605_ (_06023_, _06022_, _05879_);
  and _37606_ (_06024_, _06023_, _05921_);
  and _37607_ (_06026_, _06024_, _05751_);
  not _37608_ (_06027_, _06026_);
  and _37609_ (_06028_, _05810_, _22731_);
  and _37610_ (_06029_, _06028_, _05906_);
  and _37611_ (_06030_, _06029_, _05800_);
  and _37612_ (_06031_, _05658_, _22731_);
  and _37613_ (_06032_, _06031_, _05624_);
  nor _37614_ (_06033_, _05688_, rst);
  and _37615_ (_06034_, _06033_, _05962_);
  and _37616_ (_06035_, _06034_, _06032_);
  and _37617_ (_06036_, _06035_, word_in[7]);
  nor _37618_ (_06037_, _06035_, _05691_);
  nor _37619_ (_06038_, _06037_, _06036_);
  nor _37620_ (_06039_, _06038_, _06030_);
  and _37621_ (_06040_, _06030_, word_in[15]);
  or _37622_ (_06041_, _06040_, _06039_);
  and _37623_ (_06042_, _06041_, _06027_);
  and _37624_ (_06043_, _05991_, _22731_);
  and _37625_ (_06044_, _06043_, _05784_);
  and _37626_ (_06046_, _06044_, _05962_);
  and _37627_ (_06047_, _06022_, word_in[23]);
  and _37628_ (_06048_, _06047_, _06026_);
  or _37629_ (_06049_, _06048_, _06046_);
  or _37630_ (_06050_, _06049_, _06042_);
  not _37631_ (_06051_, _06046_);
  and _37632_ (_06052_, _06043_, word_in[31]);
  or _37633_ (_06053_, _06052_, _06051_);
  and _37634_ (_26829_[7], _06053_, _06050_);
  or _37635_ (_06055_, _05996_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _37636_ (_26839_, _06055_, _22731_);
  and _37637_ (_06057_, _04920_, _24134_);
  and _37638_ (_06058_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _37639_ (_00657_, _06058_, _06057_);
  or _37640_ (_06060_, _05965_, _05875_);
  or _37641_ (_06061_, _05982_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _37642_ (_06062_, _06061_, _06060_);
  and _37643_ (_26822_[1], _06062_, _22731_);
  and _37644_ (_06063_, _03001_, _23887_);
  and _37645_ (_06064_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _37646_ (_00674_, _06064_, _06063_);
  or _37647_ (_06066_, _05617_, _05613_);
  nor _37648_ (_06067_, _06066_, _05633_);
  or _37649_ (_06069_, _06067_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _37650_ (_06070_, _06060_, _06069_);
  and _37651_ (_26822_[2], _06070_, _22731_);
  or _37652_ (_06072_, _05667_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _37653_ (_26822_[3], _06072_, _22731_);
  and _37654_ (_06073_, _05753_, _05667_);
  and _37655_ (_06074_, _05751_, _06003_);
  and _37656_ (_06075_, _05948_, _05724_);
  and _37657_ (_06077_, _06075_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _37658_ (_06078_, _06077_, _06074_);
  not _37659_ (_06079_, _05667_);
  and _37660_ (_06080_, _05760_, _05784_);
  or _37661_ (_06081_, _06080_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _37662_ (_06082_, _06081_, _06079_);
  or _37663_ (_06083_, _06082_, _06078_);
  or _37664_ (_06084_, _06083_, _06073_);
  or _37665_ (_06085_, _06084_, _06067_);
  and _37666_ (_26822_[4], _06085_, _22731_);
  or _37667_ (_06087_, _06080_, _06073_);
  or _37668_ (_06089_, _06087_, _05883_);
  and _37669_ (_06090_, _06089_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _37670_ (_06091_, _05760_, _05751_);
  and _37671_ (_06092_, _06067_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _37672_ (_06093_, _06092_, _06091_);
  nor _37673_ (_06094_, _06093_, _06090_);
  nor _37674_ (_06096_, _06094_, _05955_);
  and _37675_ (_06097_, _05649_, _05618_);
  or _37676_ (_06098_, _06097_, _06067_);
  or _37677_ (_06099_, _06098_, _06080_);
  or _37678_ (_06100_, _06099_, _06073_);
  or _37679_ (_06101_, _06100_, _06096_);
  and _37680_ (_26822_[5], _06101_, _22731_);
  and _37681_ (_06102_, _05947_, _05724_);
  or _37682_ (_06103_, _05759_, _06102_);
  or _37683_ (_06104_, _05759_, _05725_);
  nor _37684_ (_06105_, _06066_, _05640_);
  not _37685_ (_06106_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _37686_ (_06108_, _05667_, _06106_);
  and _37687_ (_06109_, _06108_, _06066_);
  or _37688_ (_06110_, _06109_, _06105_);
  and _37689_ (_06111_, _06110_, _06104_);
  and _37690_ (_06112_, _06087_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _37691_ (_06113_, _06112_, _06091_);
  or _37692_ (_06114_, _06113_, _06111_);
  and _37693_ (_06115_, _06114_, _06103_);
  or _37694_ (_06116_, _06112_, _06110_);
  and _37695_ (_06117_, _06116_, _05965_);
  and _37696_ (_06118_, _06067_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _37697_ (_06119_, _05875_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _37698_ (_06121_, _06119_, _06073_);
  or _37699_ (_06122_, _06121_, _06118_);
  or _37700_ (_06124_, _06122_, _06080_);
  or _37701_ (_06125_, _06124_, _06117_);
  or _37702_ (_06126_, _06125_, _06115_);
  and _37703_ (_26822_[6], _06126_, _22731_);
  and _37704_ (_06127_, _24320_, _24219_);
  and _37705_ (_06128_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _37706_ (_00972_, _06128_, _06127_);
  and _37707_ (_06129_, _24496_, _24223_);
  and _37708_ (_06130_, _06129_, _23996_);
  not _37709_ (_06131_, _06129_);
  and _37710_ (_06132_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or _37711_ (_00985_, _06132_, _06130_);
  and _37712_ (_06133_, _25658_, _24219_);
  and _37713_ (_06134_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _37714_ (_00994_, _06134_, _06133_);
  or _37715_ (_06135_, _05754_, _05617_);
  or _37716_ (_06136_, _06105_, _05617_);
  and _37717_ (_06137_, _06136_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _37718_ (_06138_, _05642_, _05640_);
  or _37719_ (_06139_, _06138_, _05761_);
  or _37720_ (_06140_, _06139_, _06137_);
  and _37721_ (_06141_, _06140_, _06135_);
  and _37722_ (_06142_, _05667_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _37723_ (_06143_, _06142_, _06080_);
  or _37724_ (_06144_, _06143_, _06091_);
  or _37725_ (_06145_, _06144_, _06105_);
  or _37726_ (_06146_, _06145_, _06141_);
  and _37727_ (_26822_[7], _06146_, _22731_);
  or _37728_ (_06148_, _05957_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _37729_ (_26822_[8], _06148_, _22731_);
  and _37730_ (_06150_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and _37731_ (_06152_, _02513_, _24219_);
  or _37732_ (_01070_, _06152_, _06150_);
  nand _37733_ (_06153_, _02294_, _24082_);
  or _37734_ (_06154_, _02616_, _02281_);
  and _37735_ (_06155_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _37736_ (_06156_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _37737_ (_06157_, _06156_, _02285_);
  not _37738_ (_06158_, _02281_);
  nor _37739_ (_06159_, _02258_, _02249_);
  nor _37740_ (_06160_, _06159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _37741_ (_06162_, _02259_, _02248_);
  nor _37742_ (_06163_, _06162_, _06160_);
  and _37743_ (_06164_, _06163_, _06158_);
  nor _37744_ (_06165_, _06164_, _06157_);
  nor _37745_ (_06166_, _06165_, _02616_);
  or _37746_ (_06167_, _06166_, _06155_);
  or _37747_ (_06168_, _06167_, _02294_);
  and _37748_ (_06170_, _06168_, _22731_);
  and _37749_ (_01093_, _06170_, _06153_);
  and _37750_ (_06171_, _05759_, _06002_);
  and _37751_ (_06172_, _05725_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _37752_ (_06173_, _05751_, _06008_);
  or _37753_ (_06174_, _06173_, _05652_);
  or _37754_ (_06175_, _06174_, _06172_);
  and _37755_ (_06176_, _06175_, _06171_);
  and _37756_ (_06177_, _05948_, _05617_);
  or _37757_ (_06178_, _06172_, _06177_);
  or _37758_ (_06180_, _06178_, _06176_);
  and _37759_ (_06181_, _06180_, _05759_);
  and _37760_ (_06182_, _06175_, _05965_);
  or _37761_ (_06183_, _06091_, _06003_);
  and _37762_ (_06184_, _06183_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _37763_ (_06185_, _06075_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _37764_ (_06186_, _06185_, _05725_);
  or _37765_ (_06187_, _06186_, _06184_);
  or _37766_ (_06188_, _06187_, _06182_);
  or _37767_ (_06189_, _06188_, _06181_);
  and _37768_ (_26822_[9], _06189_, _22731_);
  and _37769_ (_06190_, _05906_, _06008_);
  not _37770_ (_06191_, _05755_);
  and _37771_ (_06192_, _06191_, _05682_);
  or _37772_ (_06193_, _06192_, _06190_);
  and _37773_ (_06194_, _05879_, _05724_);
  and _37774_ (_06195_, _06194_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _37775_ (_06196_, _06105_, _05875_);
  and _37776_ (_06197_, _06196_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _37777_ (_06198_, _06197_, _05761_);
  or _37778_ (_06199_, _06198_, _06195_);
  or _37779_ (_06200_, _06199_, _06177_);
  or _37780_ (_06201_, _06200_, _06173_);
  or _37781_ (_06202_, _06201_, _06193_);
  and _37782_ (_26822_[10], _06202_, _22731_);
  and _37783_ (_06203_, _02512_, _24140_);
  not _37784_ (_06204_, _06203_);
  and _37785_ (_06205_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _37786_ (_06206_, _06203_, _23996_);
  or _37787_ (_01196_, _06206_, _06205_);
  and _37788_ (_06208_, _24474_, _24301_);
  and _37789_ (_06209_, _06208_, _23887_);
  not _37790_ (_06210_, _06208_);
  and _37791_ (_06211_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _37792_ (_01224_, _06211_, _06209_);
  and _37793_ (_06212_, _25658_, _23583_);
  and _37794_ (_06213_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or _37795_ (_01235_, _06213_, _06212_);
  and _37796_ (_06215_, _25658_, _23887_);
  and _37797_ (_06216_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or _37798_ (_01254_, _06216_, _06215_);
  and _37799_ (_06217_, _05787_, _05667_);
  or _37800_ (_06218_, _06217_, _05766_);
  or _37801_ (_06219_, _06218_, _05962_);
  and _37802_ (_06220_, _06219_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _37803_ (_06221_, _05753_, _06008_);
  and _37804_ (_06222_, _06075_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _37805_ (_06223_, _06222_, _06177_);
  or _37806_ (_06224_, _06223_, _06173_);
  or _37807_ (_06226_, _06224_, _06190_);
  or _37808_ (_06227_, _06226_, _06221_);
  or _37809_ (_06228_, _06227_, _06220_);
  and _37810_ (_26822_[11], _06228_, _22731_);
  and _37811_ (_06230_, _25637_, _24051_);
  and _37812_ (_06231_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _37813_ (_01301_, _06231_, _06230_);
  and _37814_ (_06233_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  and _37815_ (_06234_, _02513_, _23548_);
  or _37816_ (_01307_, _06234_, _06233_);
  and _37817_ (_06236_, _02527_, _25481_);
  nand _37818_ (_06237_, _06236_, _23504_);
  or _37819_ (_06238_, _06236_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _37820_ (_06240_, _06238_, _02534_);
  and _37821_ (_06241_, _06240_, _06237_);
  nor _37822_ (_06242_, _02534_, _23989_);
  or _37823_ (_06244_, _06242_, _06241_);
  and _37824_ (_01332_, _06244_, _22731_);
  or _37825_ (_06245_, _02925_, _02865_);
  and _37826_ (_06246_, _06245_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _37827_ (_06247_, _06246_, _02898_);
  and _37828_ (_01334_, _06247_, _22731_);
  nor _37829_ (_01336_, _04686_, rst);
  and _37830_ (_06249_, _24008_, _23583_);
  and _37831_ (_06250_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or _37832_ (_27083_, _06250_, _06249_);
  or _37833_ (_06251_, _05957_, _05724_);
  and _37834_ (_06252_, _06251_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _37835_ (_06253_, _05953_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _37836_ (_06254_, _06253_, _06008_);
  or _37837_ (_06255_, _06254_, _06252_);
  and _37838_ (_26822_[12], _06255_, _22731_);
  and _37839_ (_06256_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _37840_ (_06257_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _37841_ (_01355_, _06257_, _06256_);
  or _37842_ (_06258_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _37843_ (_06259_, _06258_, _22731_);
  and _37844_ (_06260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or _37845_ (_06261_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _37846_ (_06262_, _06261_, rxd_i);
  or _37847_ (_06263_, _06262_, _06260_);
  and _37848_ (_06264_, _06263_, _02785_);
  and _37849_ (_06265_, _02812_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _37850_ (_06267_, _06265_, _06264_);
  and _37851_ (_06269_, _02799_, rxd_i);
  or _37852_ (_06270_, _06269_, _02810_);
  or _37853_ (_06271_, _06270_, _06267_);
  and _37854_ (_01368_, _06271_, _06259_);
  and _37855_ (_06272_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  and _37856_ (_06273_, _02513_, _23887_);
  or _37857_ (_01379_, _06273_, _06272_);
  and _37858_ (_06274_, _04865_, _24219_);
  and _37859_ (_06276_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _37860_ (_01388_, _06276_, _06274_);
  and _37861_ (_06278_, _06129_, _23887_);
  and _37862_ (_06279_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or _37863_ (_01392_, _06279_, _06278_);
  and _37864_ (_06281_, _02970_, _23548_);
  and _37865_ (_06283_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or _37866_ (_01404_, _06283_, _06281_);
  and _37867_ (_06284_, _06129_, _23548_);
  and _37868_ (_06286_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or _37869_ (_01407_, _06286_, _06284_);
  and _37870_ (_06287_, _02877_, _02780_);
  and _37871_ (_06289_, _02867_, _06287_);
  nand _37872_ (_06290_, _06289_, _02900_);
  or _37873_ (_06291_, _06289_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _37874_ (_06292_, _06291_, _22731_);
  and _37875_ (_01409_, _06292_, _06290_);
  and _37876_ (_06293_, _05632_, _05617_);
  or _37877_ (_06294_, _05963_, _06293_);
  and _37878_ (_06295_, _05962_, _05784_);
  and _37879_ (_06296_, _05874_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _37880_ (_06298_, _05884_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or _37881_ (_06299_, _06298_, _06296_);
  or _37882_ (_06300_, _06299_, _06295_);
  or _37883_ (_06301_, _06300_, _06294_);
  and _37884_ (_26822_[13], _06301_, _22731_);
  nor _37885_ (_06302_, _02792_, _02786_);
  and _37886_ (_06303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _02900_);
  and _37887_ (_06305_, _06303_, _02792_);
  or _37888_ (_06306_, _06305_, _06302_);
  and _37889_ (_06307_, _06306_, _02569_);
  not _37890_ (_06308_, _02798_);
  nand _37891_ (_06310_, _02824_, _06308_);
  or _37892_ (_06311_, _06310_, _06307_);
  and _37893_ (_01421_, _06311_, _02080_);
  or _37894_ (_06312_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _37895_ (_06313_, _06312_, _22731_);
  nand _37896_ (_06315_, _02071_, _23989_);
  and _37897_ (_01423_, _06315_, _06313_);
  not _37898_ (_06316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _37899_ (_06317_, _02652_, _06316_);
  or _37900_ (_06318_, _06317_, _04703_);
  and _37901_ (_06319_, _06318_, _02649_);
  nand _37902_ (_06320_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _37903_ (_06321_, _06320_, _02648_);
  nor _37904_ (_06322_, _06321_, _06319_);
  nor _37905_ (_06323_, _06322_, _02647_);
  or _37906_ (_06324_, _06323_, _02757_);
  nand _37907_ (_06325_, _06324_, _22731_);
  nor _37908_ (_01426_, _06325_, _02658_);
  or _37909_ (_06326_, _05800_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _37910_ (_26822_[14], _06326_, _22731_);
  and _37911_ (_06328_, _06129_, _24051_);
  and _37912_ (_06329_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or _37913_ (_01495_, _06329_, _06328_);
  and _37914_ (_06330_, _24008_, _23887_);
  and _37915_ (_06331_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _37916_ (_01500_, _06331_, _06330_);
  and _37917_ (_06332_, _02970_, _24219_);
  and _37918_ (_06334_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or _37919_ (_01504_, _06334_, _06332_);
  and _37920_ (_06335_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  and _37921_ (_06337_, _05596_, _23996_);
  or _37922_ (_01600_, _06337_, _06335_);
  and _37923_ (_06339_, _02039_, _24474_);
  not _37924_ (_06341_, _06339_);
  and _37925_ (_06342_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _37926_ (_06343_, _06339_, _24219_);
  or _37927_ (_01604_, _06343_, _06342_);
  and _37928_ (_06344_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _37929_ (_06345_, _06339_, _23887_);
  or _37930_ (_01606_, _06345_, _06344_);
  and _37931_ (_06347_, _03245_, _24089_);
  and _37932_ (_06348_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  or _37933_ (_27170_, _06348_, _06347_);
  and _37934_ (_06351_, _02767_, _23583_);
  and _37935_ (_06352_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or _37936_ (_01662_, _06352_, _06351_);
  and _37937_ (_06353_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _37938_ (_06354_, _06339_, _23583_);
  or _37939_ (_27015_, _06354_, _06353_);
  and _37940_ (_06356_, _25413_, _24159_);
  and _37941_ (_06357_, _06356_, _24089_);
  not _37942_ (_06358_, _06356_);
  and _37943_ (_06359_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _37944_ (_01688_, _06359_, _06357_);
  and _37945_ (_06360_, _06356_, _23887_);
  and _37946_ (_06361_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _37947_ (_01698_, _06361_, _06360_);
  and _37948_ (_06362_, _06356_, _23996_);
  and _37949_ (_06363_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _37950_ (_01729_, _06363_, _06362_);
  and _37951_ (_06364_, _06043_, word_in[24]);
  and _37952_ (_06365_, _06364_, _05963_);
  and _37953_ (_06366_, _06022_, _05982_);
  and _37954_ (_06367_, _06028_, _05965_);
  not _37955_ (_06368_, _06367_);
  and _37956_ (_06369_, _06033_, _05624_);
  nor _37957_ (_06370_, _06369_, _06031_);
  and _37958_ (_06371_, _06033_, _05667_);
  and _37959_ (_06372_, _06371_, _06370_);
  and _37960_ (_06374_, _06372_, word_in[0]);
  not _37961_ (_06375_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _37962_ (_06376_, _06372_, _06375_);
  or _37963_ (_06377_, _06376_, _06374_);
  and _37964_ (_06378_, _06377_, _06368_);
  and _37965_ (_06379_, _06367_, word_in[8]);
  or _37966_ (_06381_, _06379_, _06378_);
  or _37967_ (_06383_, _06381_, _06366_);
  and _37968_ (_06384_, _06043_, _05963_);
  not _37969_ (_06385_, _06384_);
  not _37970_ (_06386_, _06366_);
  or _37971_ (_06387_, _06386_, word_in[16]);
  and _37972_ (_06388_, _06387_, _06385_);
  and _37973_ (_06389_, _06388_, _06383_);
  or _37974_ (_26823_[0], _06389_, _06365_);
  and _37975_ (_06391_, _06022_, word_in[17]);
  and _37976_ (_06392_, _06391_, _05982_);
  not _37977_ (_06393_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _37978_ (_06394_, _06372_, _06393_);
  and _37979_ (_06395_, _06372_, word_in[1]);
  or _37980_ (_06397_, _06395_, _06394_);
  and _37981_ (_06398_, _06397_, _06368_);
  and _37982_ (_06399_, _06367_, word_in[9]);
  or _37983_ (_06400_, _06399_, _06398_);
  and _37984_ (_06402_, _06400_, _06386_);
  or _37985_ (_06404_, _06402_, _06392_);
  and _37986_ (_06405_, _06404_, _06385_);
  and _37987_ (_06406_, _06384_, word_in[25]);
  or _37988_ (_26823_[1], _06406_, _06405_);
  and _37989_ (_06407_, _06043_, word_in[26]);
  and _37990_ (_06409_, _06407_, _05963_);
  not _37991_ (_06410_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _37992_ (_06411_, _06372_, _06410_);
  and _37993_ (_06412_, _06033_, word_in[2]);
  and _37994_ (_06413_, _06412_, _06372_);
  or _37995_ (_06415_, _06413_, _06411_);
  or _37996_ (_06417_, _06415_, _06367_);
  or _37997_ (_06418_, _06368_, word_in[10]);
  and _37998_ (_06419_, _06418_, _06417_);
  or _37999_ (_06421_, _06419_, _06366_);
  or _38000_ (_06422_, _06386_, word_in[18]);
  and _38001_ (_06423_, _06422_, _06385_);
  and _38002_ (_06424_, _06423_, _06421_);
  or _38003_ (_26823_[2], _06424_, _06409_);
  not _38004_ (_06425_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _38005_ (_06426_, _06372_, _06425_);
  and _38006_ (_06427_, _06033_, word_in[3]);
  and _38007_ (_06429_, _06427_, _06372_);
  or _38008_ (_06430_, _06429_, _06426_);
  or _38009_ (_06431_, _06430_, _06367_);
  or _38010_ (_06432_, _06368_, word_in[11]);
  and _38011_ (_06433_, _06432_, _06431_);
  or _38012_ (_06435_, _06433_, _06366_);
  or _38013_ (_06437_, _06386_, word_in[19]);
  and _38014_ (_06438_, _06437_, _06385_);
  and _38015_ (_06440_, _06438_, _06435_);
  and _38016_ (_06441_, _06043_, word_in[27]);
  and _38017_ (_06443_, _06441_, _05963_);
  or _38018_ (_26823_[3], _06443_, _06440_);
  and _38019_ (_06446_, _06043_, word_in[28]);
  and _38020_ (_06447_, _06446_, _05963_);
  not _38021_ (_06448_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _38022_ (_06449_, _06372_, _06448_);
  and _38023_ (_06450_, _06033_, word_in[4]);
  and _38024_ (_06451_, _06450_, _06372_);
  or _38025_ (_06452_, _06451_, _06449_);
  or _38026_ (_06453_, _06452_, _06367_);
  or _38027_ (_06454_, _06368_, word_in[12]);
  and _38028_ (_06455_, _06454_, _06453_);
  or _38029_ (_06456_, _06455_, _06366_);
  or _38030_ (_06458_, _06386_, word_in[20]);
  and _38031_ (_06460_, _06458_, _06385_);
  and _38032_ (_06461_, _06460_, _06456_);
  or _38033_ (_26823_[4], _06461_, _06447_);
  and _38034_ (_06463_, _06043_, word_in[29]);
  and _38035_ (_06464_, _06463_, _05963_);
  not _38036_ (_06466_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _38037_ (_06468_, _06372_, _06466_);
  and _38038_ (_06469_, _06033_, word_in[5]);
  and _38039_ (_06470_, _06469_, _06372_);
  or _38040_ (_06471_, _06470_, _06468_);
  or _38041_ (_06472_, _06471_, _06367_);
  or _38042_ (_06473_, _06368_, word_in[13]);
  and _38043_ (_06474_, _06473_, _06472_);
  or _38044_ (_06475_, _06474_, _06366_);
  or _38045_ (_06476_, _06386_, word_in[21]);
  and _38046_ (_06478_, _06476_, _06385_);
  and _38047_ (_06479_, _06478_, _06475_);
  or _38048_ (_26823_[5], _06479_, _06464_);
  and _38049_ (_06480_, _06384_, word_in[30]);
  not _38050_ (_06481_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _38051_ (_06482_, _06372_, _06481_);
  and _38052_ (_06483_, _06372_, word_in[6]);
  or _38053_ (_06484_, _06483_, _06482_);
  and _38054_ (_06486_, _06484_, _06368_);
  and _38055_ (_06487_, _06367_, word_in[14]);
  or _38056_ (_06488_, _06487_, _06486_);
  or _38057_ (_06489_, _06488_, _06366_);
  or _38058_ (_06490_, _06386_, word_in[22]);
  and _38059_ (_06491_, _06490_, _06385_);
  and _38060_ (_06492_, _06491_, _06489_);
  or _38061_ (_26823_[6], _06492_, _06480_);
  and _38062_ (_06493_, _24442_, _23583_);
  and _38063_ (_06494_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or _38064_ (_01799_, _06494_, _06493_);
  nor _38065_ (_06495_, _06372_, _05842_);
  and _38066_ (_06496_, _06033_, word_in[7]);
  and _38067_ (_06497_, _06372_, _06496_);
  or _38068_ (_06498_, _06497_, _06495_);
  or _38069_ (_06499_, _06498_, _06367_);
  or _38070_ (_06500_, _06368_, word_in[15]);
  and _38071_ (_06502_, _06500_, _06499_);
  or _38072_ (_06503_, _06502_, _06366_);
  or _38073_ (_06505_, _06386_, word_in[23]);
  and _38074_ (_06507_, _06505_, _06385_);
  and _38075_ (_06508_, _06507_, _06503_);
  and _38076_ (_06509_, _06384_, word_in[31]);
  or _38077_ (_26823_[7], _06509_, _06508_);
  and _38078_ (_06512_, _06022_, _05753_);
  and _38079_ (_06513_, _06512_, _05876_);
  and _38080_ (_06515_, _06028_, _05784_);
  and _38081_ (_06516_, _06515_, _05767_);
  not _38082_ (_06518_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _38083_ (_06520_, _06033_, _06079_);
  and _38084_ (_06521_, _06031_, _05625_);
  not _38085_ (_06522_, _06521_);
  nor _38086_ (_06523_, _06522_, _06520_);
  nor _38087_ (_06524_, _06523_, _06518_);
  and _38088_ (_06525_, _06033_, word_in[0]);
  and _38089_ (_06527_, _06523_, _06525_);
  or _38090_ (_06528_, _06527_, _06524_);
  or _38091_ (_06529_, _06528_, _06516_);
  not _38092_ (_06531_, _06516_);
  or _38093_ (_06532_, _06531_, word_in[8]);
  and _38094_ (_06533_, _06532_, _06529_);
  or _38095_ (_06534_, _06533_, _06513_);
  and _38096_ (_06535_, _06043_, _05982_);
  not _38097_ (_06537_, _06535_);
  and _38098_ (_06538_, _06022_, word_in[16]);
  not _38099_ (_06539_, _06513_);
  or _38100_ (_06540_, _06539_, _06538_);
  and _38101_ (_06542_, _06540_, _06537_);
  and _38102_ (_06543_, _06542_, _06534_);
  and _38103_ (_06544_, _06535_, word_in[24]);
  or _38104_ (_26830_[0], _06544_, _06543_);
  not _38105_ (_06545_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _38106_ (_06546_, _06523_, _06545_);
  and _38107_ (_06548_, _06033_, word_in[1]);
  and _38108_ (_06549_, _06523_, _06548_);
  or _38109_ (_06550_, _06549_, _06546_);
  or _38110_ (_06551_, _06550_, _06516_);
  or _38111_ (_06552_, _06531_, word_in[9]);
  and _38112_ (_06553_, _06552_, _06551_);
  or _38113_ (_06554_, _06553_, _06513_);
  or _38114_ (_06556_, _06539_, _06391_);
  and _38115_ (_06557_, _06556_, _06537_);
  and _38116_ (_06559_, _06557_, _06554_);
  and _38117_ (_06561_, _06535_, word_in[25]);
  or _38118_ (_26830_[1], _06561_, _06559_);
  not _38119_ (_06562_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _38120_ (_06563_, _06523_, _06562_);
  and _38121_ (_06565_, _06523_, _06412_);
  or _38122_ (_06566_, _06565_, _06563_);
  or _38123_ (_06567_, _06566_, _06516_);
  or _38124_ (_06568_, _06531_, word_in[10]);
  and _38125_ (_06570_, _06568_, _06567_);
  or _38126_ (_06571_, _06570_, _06513_);
  and _38127_ (_06572_, _06022_, word_in[18]);
  or _38128_ (_06573_, _06539_, _06572_);
  and _38129_ (_06575_, _06573_, _06537_);
  and _38130_ (_06576_, _06575_, _06571_);
  and _38131_ (_06577_, _06535_, word_in[26]);
  or _38132_ (_26830_[2], _06577_, _06576_);
  not _38133_ (_06578_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _38134_ (_06579_, _06523_, _06578_);
  and _38135_ (_06580_, _06523_, _06427_);
  or _38136_ (_06581_, _06580_, _06579_);
  or _38137_ (_06582_, _06581_, _06516_);
  or _38138_ (_06583_, _06531_, word_in[11]);
  and _38139_ (_06584_, _06583_, _06582_);
  or _38140_ (_06585_, _06584_, _06513_);
  and _38141_ (_06586_, _06022_, word_in[19]);
  or _38142_ (_06587_, _06539_, _06586_);
  and _38143_ (_06588_, _06587_, _06537_);
  and _38144_ (_06589_, _06588_, _06585_);
  and _38145_ (_06590_, _06535_, word_in[27]);
  or _38146_ (_26830_[3], _06590_, _06589_);
  and _38147_ (_06591_, _06022_, word_in[20]);
  and _38148_ (_06592_, _06513_, _06591_);
  and _38149_ (_06593_, _06523_, _06450_);
  not _38150_ (_06594_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _38151_ (_06595_, _06523_, _06594_);
  nor _38152_ (_06596_, _06595_, _06593_);
  nor _38153_ (_06597_, _06596_, _06516_);
  and _38154_ (_06598_, _06516_, word_in[12]);
  or _38155_ (_06599_, _06598_, _06597_);
  and _38156_ (_06600_, _06599_, _06539_);
  or _38157_ (_06602_, _06600_, _06592_);
  and _38158_ (_06603_, _06602_, _06537_);
  and _38159_ (_06605_, _06535_, word_in[28]);
  or _38160_ (_26830_[4], _06605_, _06603_);
  and _38161_ (_06606_, _06022_, word_in[21]);
  and _38162_ (_06607_, _06513_, _06606_);
  and _38163_ (_06608_, _06523_, _06469_);
  not _38164_ (_06609_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _38165_ (_06610_, _06523_, _06609_);
  nor _38166_ (_06611_, _06610_, _06608_);
  nor _38167_ (_06612_, _06611_, _06516_);
  and _38168_ (_06613_, _06516_, word_in[13]);
  or _38169_ (_06615_, _06613_, _06612_);
  and _38170_ (_06616_, _06615_, _06539_);
  or _38171_ (_06617_, _06616_, _06607_);
  and _38172_ (_06618_, _06617_, _06537_);
  and _38173_ (_06619_, _06535_, word_in[29]);
  or _38174_ (_26830_[5], _06619_, _06618_);
  and _38175_ (_06620_, _06022_, word_in[22]);
  and _38176_ (_06621_, _06513_, _06620_);
  and _38177_ (_06623_, _06033_, word_in[6]);
  and _38178_ (_06624_, _06523_, _06623_);
  not _38179_ (_06625_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _38180_ (_06626_, _06523_, _06625_);
  nor _38181_ (_06628_, _06626_, _06624_);
  nor _38182_ (_06629_, _06628_, _06516_);
  and _38183_ (_06630_, _06516_, word_in[14]);
  or _38184_ (_06631_, _06630_, _06629_);
  and _38185_ (_06632_, _06631_, _06539_);
  or _38186_ (_06633_, _06632_, _06621_);
  and _38187_ (_06634_, _06633_, _06537_);
  and _38188_ (_06635_, _06535_, word_in[30]);
  or _38189_ (_26830_[6], _06635_, _06634_);
  and _38190_ (_06636_, _06513_, _06047_);
  and _38191_ (_06637_, _06523_, _06496_);
  nor _38192_ (_06638_, _06523_, _05737_);
  nor _38193_ (_06639_, _06638_, _06637_);
  nor _38194_ (_06640_, _06639_, _06516_);
  and _38195_ (_06641_, _06516_, word_in[15]);
  or _38196_ (_06642_, _06641_, _06640_);
  and _38197_ (_06643_, _06642_, _06539_);
  or _38198_ (_06644_, _06643_, _06636_);
  and _38199_ (_06645_, _06644_, _06537_);
  and _38200_ (_06646_, _06535_, word_in[31]);
  or _38201_ (_26830_[7], _06646_, _06645_);
  and _38202_ (_06647_, _06043_, _05753_);
  and _38203_ (_06648_, _06647_, _05996_);
  and _38204_ (_06649_, _06022_, _05784_);
  and _38205_ (_06650_, _06649_, _05876_);
  not _38206_ (_06651_, _06650_);
  or _38207_ (_06652_, _06651_, _06538_);
  and _38208_ (_06653_, _06028_, _05751_);
  and _38209_ (_06654_, _06653_, _05767_);
  not _38210_ (_06655_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not _38211_ (_06656_, _06031_);
  and _38212_ (_06657_, _06369_, _06656_);
  and _38213_ (_06658_, _06657_, _05667_);
  nor _38214_ (_06659_, _06658_, _06655_);
  and _38215_ (_06660_, _06658_, _06525_);
  or _38216_ (_06661_, _06660_, _06659_);
  or _38217_ (_06662_, _06661_, _06654_);
  not _38218_ (_06663_, _06654_);
  or _38219_ (_06664_, _06663_, word_in[8]);
  and _38220_ (_06665_, _06664_, _06662_);
  or _38221_ (_06666_, _06665_, _06650_);
  and _38222_ (_06668_, _06666_, _06652_);
  or _38223_ (_06669_, _06668_, _06648_);
  not _38224_ (_06670_, _06648_);
  or _38225_ (_06671_, _06670_, word_in[24]);
  and _38226_ (_26831_[0], _06671_, _06669_);
  and _38227_ (_06672_, _06650_, _06391_);
  and _38228_ (_06673_, _06658_, _06548_);
  not _38229_ (_06674_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _38230_ (_06675_, _06658_, _06674_);
  nor _38231_ (_06676_, _06675_, _06673_);
  nor _38232_ (_06677_, _06676_, _06654_);
  and _38233_ (_06678_, _06654_, word_in[9]);
  or _38234_ (_06679_, _06678_, _06677_);
  and _38235_ (_06680_, _06679_, _06651_);
  or _38236_ (_06682_, _06680_, _06672_);
  and _38237_ (_06683_, _06682_, _06670_);
  and _38238_ (_06684_, _06648_, word_in[25]);
  or _38239_ (_26831_[1], _06684_, _06683_);
  and _38240_ (_06685_, _06658_, _06412_);
  not _38241_ (_06686_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _38242_ (_06687_, _06658_, _06686_);
  nor _38243_ (_06688_, _06687_, _06685_);
  nor _38244_ (_06689_, _06688_, _06654_);
  and _38245_ (_06690_, _06654_, word_in[10]);
  or _38246_ (_06691_, _06690_, _06689_);
  and _38247_ (_06692_, _06691_, _06651_);
  and _38248_ (_06693_, _06650_, _06572_);
  or _38249_ (_06694_, _06693_, _06648_);
  or _38250_ (_06695_, _06694_, _06692_);
  or _38251_ (_06696_, _06670_, word_in[26]);
  and _38252_ (_26831_[2], _06696_, _06695_);
  and _38253_ (_06697_, _06650_, _06586_);
  and _38254_ (_06698_, _06658_, _06427_);
  not _38255_ (_06699_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _38256_ (_06700_, _06658_, _06699_);
  nor _38257_ (_06702_, _06700_, _06698_);
  nor _38258_ (_06703_, _06702_, _06654_);
  and _38259_ (_06704_, _06654_, word_in[11]);
  or _38260_ (_06705_, _06704_, _06703_);
  and _38261_ (_06706_, _06705_, _06651_);
  or _38262_ (_06708_, _06706_, _06697_);
  and _38263_ (_06709_, _06708_, _06670_);
  and _38264_ (_06710_, _06648_, word_in[27]);
  or _38265_ (_26831_[3], _06710_, _06709_);
  not _38266_ (_06711_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _38267_ (_06712_, _06658_, _06711_);
  and _38268_ (_06713_, _06658_, _06450_);
  or _38269_ (_06714_, _06713_, _06712_);
  or _38270_ (_06715_, _06714_, _06654_);
  or _38271_ (_06716_, _06663_, word_in[12]);
  and _38272_ (_06717_, _06716_, _06715_);
  or _38273_ (_06718_, _06717_, _06650_);
  or _38274_ (_06719_, _06651_, _06591_);
  and _38275_ (_06720_, _06719_, _06670_);
  and _38276_ (_06721_, _06720_, _06718_);
  and _38277_ (_06723_, _06648_, word_in[28]);
  or _38278_ (_26831_[4], _06723_, _06721_);
  and _38279_ (_06724_, _06650_, _06606_);
  and _38280_ (_06725_, _06658_, _06469_);
  not _38281_ (_06726_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _38282_ (_06727_, _06658_, _06726_);
  nor _38283_ (_06728_, _06727_, _06725_);
  nor _38284_ (_06729_, _06728_, _06654_);
  and _38285_ (_06730_, _06654_, word_in[13]);
  or _38286_ (_06731_, _06730_, _06729_);
  and _38287_ (_06733_, _06731_, _06651_);
  or _38288_ (_06734_, _06733_, _06724_);
  and _38289_ (_06735_, _06734_, _06670_);
  and _38290_ (_06736_, _06648_, word_in[29]);
  or _38291_ (_26831_[5], _06736_, _06735_);
  and _38292_ (_06737_, _06658_, _06623_);
  not _38293_ (_06738_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _38294_ (_06739_, _06658_, _06738_);
  nor _38295_ (_06740_, _06739_, _06737_);
  nor _38296_ (_06741_, _06740_, _06654_);
  and _38297_ (_06742_, _06654_, word_in[14]);
  or _38298_ (_06743_, _06742_, _06741_);
  and _38299_ (_06745_, _06743_, _06651_);
  and _38300_ (_06746_, _06650_, _06620_);
  or _38301_ (_06747_, _06746_, _06648_);
  or _38302_ (_06748_, _06747_, _06745_);
  or _38303_ (_06749_, _06670_, word_in[30]);
  and _38304_ (_26831_[6], _06749_, _06748_);
  and _38305_ (_06750_, _06658_, _06496_);
  nor _38306_ (_06751_, _06658_, _05848_);
  nor _38307_ (_06753_, _06751_, _06750_);
  nor _38308_ (_06754_, _06753_, _06654_);
  and _38309_ (_06755_, _06654_, word_in[15]);
  or _38310_ (_06756_, _06755_, _06754_);
  and _38311_ (_06757_, _06756_, _06651_);
  and _38312_ (_06758_, _06650_, _06047_);
  or _38313_ (_06759_, _06758_, _06648_);
  or _38314_ (_06761_, _06759_, _06757_);
  or _38315_ (_06762_, _06670_, word_in[31]);
  and _38316_ (_26831_[7], _06762_, _06761_);
  and _38317_ (_06763_, _24899_, _24006_);
  and _38318_ (_06764_, _06763_, _24219_);
  not _38319_ (_06765_, _06763_);
  and _38320_ (_06766_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or _38321_ (_01925_, _06766_, _06764_);
  and _38322_ (_06767_, _06022_, _05751_);
  and _38323_ (_06768_, _06767_, _05876_);
  not _38324_ (_06769_, _06768_);
  and _38325_ (_06770_, _06029_, _05767_);
  not _38326_ (_06771_, _06032_);
  nor _38327_ (_06773_, _06520_, _06771_);
  and _38328_ (_06774_, _06773_, _06525_);
  not _38329_ (_06775_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _38330_ (_06776_, _06773_, _06775_);
  nor _38331_ (_06777_, _06776_, _06774_);
  nor _38332_ (_06778_, _06777_, _06770_);
  and _38333_ (_06779_, _06770_, word_in[8]);
  or _38334_ (_06780_, _06779_, _06778_);
  and _38335_ (_06781_, _06780_, _06769_);
  and _38336_ (_06782_, _06044_, _05996_);
  and _38337_ (_06783_, _06768_, _06538_);
  or _38338_ (_06784_, _06783_, _06782_);
  or _38339_ (_06785_, _06784_, _06781_);
  not _38340_ (_06786_, _06782_);
  or _38341_ (_06788_, _06786_, _06364_);
  and _38342_ (_26832_[0], _06788_, _06785_);
  and _38343_ (_06789_, _06773_, _06548_);
  not _38344_ (_06790_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _38345_ (_06791_, _06773_, _06790_);
  nor _38346_ (_06792_, _06791_, _06789_);
  nor _38347_ (_06794_, _06792_, _06770_);
  and _38348_ (_06795_, _06770_, word_in[9]);
  or _38349_ (_06796_, _06795_, _06794_);
  and _38350_ (_06797_, _06796_, _06769_);
  and _38351_ (_06798_, _06768_, _06391_);
  or _38352_ (_06799_, _06798_, _06782_);
  or _38353_ (_06800_, _06799_, _06797_);
  and _38354_ (_06801_, _06043_, word_in[25]);
  or _38355_ (_06802_, _06786_, _06801_);
  and _38356_ (_26832_[1], _06802_, _06800_);
  and _38357_ (_06803_, _06773_, _06412_);
  not _38358_ (_06804_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _38359_ (_06805_, _06773_, _06804_);
  nor _38360_ (_06807_, _06805_, _06803_);
  nor _38361_ (_06808_, _06807_, _06770_);
  and _38362_ (_06809_, _06770_, word_in[10]);
  or _38363_ (_06810_, _06809_, _06808_);
  and _38364_ (_06811_, _06810_, _06769_);
  and _38365_ (_06812_, _06768_, _06572_);
  or _38366_ (_06813_, _06812_, _06782_);
  or _38367_ (_06815_, _06813_, _06811_);
  or _38368_ (_06816_, _06786_, _06407_);
  and _38369_ (_26832_[2], _06816_, _06815_);
  not _38370_ (_06818_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _38371_ (_06819_, _06773_, _06818_);
  and _38372_ (_06820_, _06773_, _06427_);
  or _38373_ (_06821_, _06820_, _06819_);
  or _38374_ (_06822_, _06821_, _06770_);
  not _38375_ (_06824_, _06770_);
  or _38376_ (_06825_, _06824_, word_in[11]);
  and _38377_ (_06826_, _06825_, _06822_);
  or _38378_ (_06827_, _06826_, _06768_);
  or _38379_ (_06828_, _06769_, _06586_);
  and _38380_ (_06829_, _06828_, _06786_);
  and _38381_ (_06830_, _06829_, _06827_);
  and _38382_ (_06831_, _06782_, _06441_);
  or _38383_ (_26832_[3], _06831_, _06830_);
  not _38384_ (_06832_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _38385_ (_06833_, _06773_, _06832_);
  and _38386_ (_06834_, _06773_, _06450_);
  or _38387_ (_06835_, _06834_, _06833_);
  or _38388_ (_06836_, _06835_, _06770_);
  or _38389_ (_06837_, _06824_, word_in[12]);
  and _38390_ (_06838_, _06837_, _06836_);
  or _38391_ (_06839_, _06838_, _06768_);
  or _38392_ (_06840_, _06769_, _06591_);
  and _38393_ (_06841_, _06840_, _06786_);
  and _38394_ (_06842_, _06841_, _06839_);
  and _38395_ (_06843_, _06782_, _06446_);
  or _38396_ (_26832_[4], _06843_, _06842_);
  and _38397_ (_06844_, _06773_, _06469_);
  not _38398_ (_06845_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _38399_ (_06846_, _06773_, _06845_);
  nor _38400_ (_06847_, _06846_, _06844_);
  nor _38401_ (_06848_, _06847_, _06770_);
  and _38402_ (_06849_, _06770_, word_in[13]);
  or _38403_ (_06850_, _06849_, _06848_);
  and _38404_ (_06851_, _06850_, _06769_);
  and _38405_ (_06852_, _06768_, _06606_);
  or _38406_ (_06853_, _06852_, _06782_);
  or _38407_ (_06854_, _06853_, _06851_);
  or _38408_ (_06855_, _06786_, _06463_);
  and _38409_ (_26832_[5], _06855_, _06854_);
  and _38410_ (_06856_, _06773_, _06623_);
  not _38411_ (_06857_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _38412_ (_06858_, _06773_, _06857_);
  nor _38413_ (_06859_, _06858_, _06856_);
  nor _38414_ (_06860_, _06859_, _06770_);
  and _38415_ (_06861_, _06770_, word_in[14]);
  or _38416_ (_06862_, _06861_, _06860_);
  and _38417_ (_06863_, _06862_, _06769_);
  and _38418_ (_06864_, _06768_, _06620_);
  or _38419_ (_06865_, _06864_, _06782_);
  or _38420_ (_06866_, _06865_, _06863_);
  and _38421_ (_06867_, _06043_, word_in[30]);
  or _38422_ (_06868_, _06786_, _06867_);
  and _38423_ (_26832_[6], _06868_, _06866_);
  and _38424_ (_06870_, _06773_, _06496_);
  nor _38425_ (_06871_, _06773_, _05719_);
  nor _38426_ (_06872_, _06871_, _06870_);
  nor _38427_ (_06873_, _06872_, _06770_);
  and _38428_ (_06874_, _06770_, word_in[15]);
  or _38429_ (_06875_, _06874_, _06873_);
  and _38430_ (_06876_, _06875_, _06769_);
  and _38431_ (_06877_, _06768_, _06047_);
  or _38432_ (_06878_, _06877_, _06782_);
  or _38433_ (_06879_, _06878_, _06876_);
  or _38434_ (_06880_, _06786_, _06052_);
  and _38435_ (_26832_[7], _06880_, _06879_);
  and _38436_ (_06882_, _06043_, _06074_);
  not _38437_ (_06883_, _06882_);
  not _38438_ (_06884_, _05921_);
  and _38439_ (_06885_, _06023_, _06884_);
  and _38440_ (_06887_, _06885_, _05906_);
  and _38441_ (_06888_, _06887_, _06538_);
  not _38442_ (_06889_, _06887_);
  and _38443_ (_06890_, _06028_, _06073_);
  not _38444_ (_06891_, _06890_);
  not _38445_ (_06892_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _38446_ (_06893_, _06033_, _05760_);
  and _38447_ (_06895_, _06893_, _06370_);
  nor _38448_ (_06896_, _06895_, _06892_);
  and _38449_ (_06898_, _06895_, word_in[0]);
  or _38450_ (_06899_, _06898_, _06896_);
  and _38451_ (_06900_, _06899_, _06891_);
  and _38452_ (_06901_, _06890_, word_in[8]);
  or _38453_ (_06902_, _06901_, _06900_);
  and _38454_ (_06903_, _06902_, _06889_);
  or _38455_ (_06904_, _06903_, _06888_);
  and _38456_ (_06905_, _06904_, _06883_);
  and _38457_ (_06906_, _06882_, word_in[24]);
  or _38458_ (_26833_[0], _06906_, _06905_);
  and _38459_ (_06907_, _06887_, _06391_);
  not _38460_ (_06908_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _38461_ (_06909_, _06895_, _06908_);
  and _38462_ (_06910_, _06895_, word_in[1]);
  or _38463_ (_06911_, _06910_, _06909_);
  and _38464_ (_06912_, _06911_, _06891_);
  and _38465_ (_06913_, _06890_, word_in[9]);
  or _38466_ (_06914_, _06913_, _06912_);
  and _38467_ (_06915_, _06914_, _06889_);
  or _38468_ (_06916_, _06915_, _06907_);
  and _38469_ (_06917_, _06916_, _06883_);
  and _38470_ (_06918_, _06882_, word_in[25]);
  or _38471_ (_26833_[1], _06918_, _06917_);
  and _38472_ (_06919_, _06887_, _06572_);
  not _38473_ (_06920_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _38474_ (_06921_, _06895_, _06920_);
  and _38475_ (_06922_, _06895_, word_in[2]);
  or _38476_ (_06924_, _06922_, _06921_);
  and _38477_ (_06925_, _06924_, _06891_);
  and _38478_ (_06926_, _06890_, word_in[10]);
  or _38479_ (_06927_, _06926_, _06925_);
  and _38480_ (_06929_, _06927_, _06889_);
  or _38481_ (_06930_, _06929_, _06919_);
  and _38482_ (_06931_, _06930_, _06883_);
  and _38483_ (_06932_, _06882_, word_in[26]);
  or _38484_ (_26833_[2], _06932_, _06931_);
  and _38485_ (_06933_, _06887_, _06586_);
  not _38486_ (_06934_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _38487_ (_06935_, _06895_, _06934_);
  and _38488_ (_06936_, _06895_, word_in[3]);
  or _38489_ (_06937_, _06936_, _06935_);
  and _38490_ (_06938_, _06937_, _06891_);
  and _38491_ (_06939_, _06890_, word_in[11]);
  or _38492_ (_06940_, _06939_, _06938_);
  and _38493_ (_06941_, _06940_, _06889_);
  or _38494_ (_06942_, _06941_, _06933_);
  and _38495_ (_06943_, _06942_, _06883_);
  and _38496_ (_06944_, _06882_, word_in[27]);
  or _38497_ (_26833_[3], _06944_, _06943_);
  and _38498_ (_06945_, _06887_, _06591_);
  not _38499_ (_06946_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _38500_ (_06947_, _06895_, _06946_);
  and _38501_ (_06949_, _06895_, word_in[4]);
  or _38502_ (_06950_, _06949_, _06947_);
  and _38503_ (_06951_, _06950_, _06891_);
  and _38504_ (_06952_, _06890_, word_in[12]);
  or _38505_ (_06953_, _06952_, _06951_);
  and _38506_ (_06954_, _06953_, _06889_);
  or _38507_ (_06956_, _06954_, _06945_);
  and _38508_ (_06957_, _06956_, _06883_);
  and _38509_ (_06958_, _06882_, word_in[28]);
  or _38510_ (_26833_[4], _06958_, _06957_);
  and _38511_ (_06959_, _06887_, _06606_);
  not _38512_ (_06961_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _38513_ (_06962_, _06895_, _06961_);
  and _38514_ (_06963_, _06895_, word_in[5]);
  or _38515_ (_06965_, _06963_, _06962_);
  and _38516_ (_06966_, _06965_, _06891_);
  and _38517_ (_06968_, _06890_, word_in[13]);
  or _38518_ (_06969_, _06968_, _06966_);
  and _38519_ (_06970_, _06969_, _06889_);
  or _38520_ (_06971_, _06970_, _06959_);
  and _38521_ (_06972_, _06971_, _06883_);
  and _38522_ (_06973_, _06882_, word_in[29]);
  or _38523_ (_26833_[5], _06973_, _06972_);
  and _38524_ (_06975_, _06887_, _06620_);
  not _38525_ (_06976_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _38526_ (_06977_, _06895_, _06976_);
  and _38527_ (_06979_, _06895_, word_in[6]);
  or _38528_ (_06981_, _06979_, _06977_);
  and _38529_ (_06982_, _06981_, _06891_);
  and _38530_ (_06984_, _06890_, word_in[14]);
  or _38531_ (_06985_, _06984_, _06982_);
  and _38532_ (_06986_, _06985_, _06889_);
  or _38533_ (_06987_, _06986_, _06975_);
  and _38534_ (_06989_, _06987_, _06883_);
  and _38535_ (_06991_, _06882_, word_in[30]);
  or _38536_ (_26833_[6], _06991_, _06989_);
  and _38537_ (_06993_, _06887_, _06047_);
  nor _38538_ (_06995_, _06895_, _05855_);
  and _38539_ (_06996_, _06895_, word_in[7]);
  or _38540_ (_06998_, _06996_, _06995_);
  and _38541_ (_07000_, _06998_, _06891_);
  and _38542_ (_07001_, _06890_, word_in[15]);
  or _38543_ (_07002_, _07001_, _07000_);
  and _38544_ (_07004_, _07002_, _06889_);
  or _38545_ (_07005_, _07004_, _06993_);
  and _38546_ (_07006_, _07005_, _06883_);
  and _38547_ (_07007_, _06882_, word_in[31]);
  or _38548_ (_26833_[7], _07007_, _07006_);
  and _38549_ (_07008_, _04920_, _24219_);
  and _38550_ (_07009_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _38551_ (_02030_, _07009_, _07008_);
  and _38552_ (_07011_, _06763_, _23887_);
  and _38553_ (_07012_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _38554_ (_02042_, _07012_, _07011_);
  and _38555_ (_07013_, _24095_, _24006_);
  and _38556_ (_07014_, _07013_, _23548_);
  not _38557_ (_07015_, _07013_);
  and _38558_ (_07016_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _38559_ (_02052_, _07016_, _07014_);
  and _38560_ (_07017_, _06043_, _06067_);
  not _38561_ (_07018_, _07017_);
  and _38562_ (_07019_, _06885_, _05753_);
  and _38563_ (_07020_, _07019_, _06538_);
  not _38564_ (_07021_, _07019_);
  and _38565_ (_07022_, _06515_, _05797_);
  not _38566_ (_07023_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _38567_ (_07025_, _06893_, _06521_);
  nor _38568_ (_07026_, _07025_, _07023_);
  and _38569_ (_07027_, _07025_, word_in[0]);
  nor _38570_ (_07028_, _07027_, _07026_);
  nor _38571_ (_07029_, _07028_, _07022_);
  and _38572_ (_07030_, _07022_, word_in[8]);
  or _38573_ (_07031_, _07030_, _07029_);
  and _38574_ (_07032_, _07031_, _07021_);
  or _38575_ (_07034_, _07032_, _07020_);
  and _38576_ (_07035_, _07034_, _07018_);
  and _38577_ (_07036_, _07017_, word_in[24]);
  or _38578_ (_26834_[0], _07036_, _07035_);
  and _38579_ (_07038_, _24349_, _24301_);
  and _38580_ (_07040_, _07038_, _23996_);
  not _38581_ (_07041_, _07038_);
  and _38582_ (_07042_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _38583_ (_27227_, _07042_, _07040_);
  and _38584_ (_07044_, _07019_, _06391_);
  and _38585_ (_07045_, _07025_, word_in[1]);
  not _38586_ (_07046_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _38587_ (_07048_, _07025_, _07046_);
  nor _38588_ (_07050_, _07048_, _07045_);
  nor _38589_ (_07052_, _07050_, _07022_);
  and _38590_ (_07053_, _07022_, word_in[9]);
  or _38591_ (_07055_, _07053_, _07052_);
  and _38592_ (_07056_, _07055_, _07021_);
  or _38593_ (_07057_, _07056_, _07044_);
  and _38594_ (_07058_, _07057_, _07018_);
  and _38595_ (_07060_, _07017_, word_in[25]);
  or _38596_ (_26834_[1], _07060_, _07058_);
  and _38597_ (_07062_, _07017_, word_in[26]);
  not _38598_ (_07063_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _38599_ (_07064_, _07025_, _07063_);
  and _38600_ (_07065_, _07025_, _06412_);
  or _38601_ (_07066_, _07065_, _07064_);
  or _38602_ (_07067_, _07066_, _07022_);
  not _38603_ (_07068_, _07022_);
  or _38604_ (_07069_, _07068_, word_in[10]);
  and _38605_ (_07070_, _07069_, _07067_);
  or _38606_ (_07071_, _07070_, _07019_);
  or _38607_ (_07073_, _07021_, _06572_);
  and _38608_ (_07074_, _07073_, _07018_);
  and _38609_ (_07076_, _07074_, _07071_);
  or _38610_ (_26834_[2], _07076_, _07062_);
  and _38611_ (_07077_, _07017_, word_in[27]);
  not _38612_ (_07078_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _38613_ (_07079_, _07025_, _07078_);
  and _38614_ (_07080_, _07025_, _06427_);
  or _38615_ (_07082_, _07080_, _07079_);
  or _38616_ (_07084_, _07082_, _07022_);
  or _38617_ (_07085_, _07068_, word_in[11]);
  and _38618_ (_07086_, _07085_, _07084_);
  or _38619_ (_07087_, _07086_, _07019_);
  or _38620_ (_07088_, _07021_, _06586_);
  and _38621_ (_07090_, _07088_, _07018_);
  and _38622_ (_07091_, _07090_, _07087_);
  or _38623_ (_26834_[3], _07091_, _07077_);
  and _38624_ (_07093_, _07019_, _06591_);
  and _38625_ (_07095_, _07025_, word_in[4]);
  not _38626_ (_07096_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _38627_ (_07097_, _07025_, _07096_);
  nor _38628_ (_07098_, _07097_, _07095_);
  nor _38629_ (_07099_, _07098_, _07022_);
  and _38630_ (_07101_, _07022_, word_in[12]);
  or _38631_ (_07102_, _07101_, _07099_);
  and _38632_ (_07104_, _07102_, _07021_);
  or _38633_ (_07105_, _07104_, _07093_);
  and _38634_ (_07106_, _07105_, _07018_);
  and _38635_ (_07108_, _07017_, word_in[28]);
  or _38636_ (_26834_[4], _07108_, _07106_);
  and _38637_ (_07110_, _07017_, word_in[29]);
  and _38638_ (_07111_, _07025_, word_in[5]);
  not _38639_ (_07112_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _38640_ (_07114_, _07025_, _07112_);
  nor _38641_ (_07116_, _07114_, _07111_);
  nor _38642_ (_07118_, _07116_, _07022_);
  and _38643_ (_07119_, _07022_, word_in[13]);
  or _38644_ (_07120_, _07119_, _07118_);
  or _38645_ (_07121_, _07120_, _07019_);
  or _38646_ (_07122_, _07021_, _06606_);
  and _38647_ (_07124_, _07122_, _07018_);
  and _38648_ (_07126_, _07124_, _07121_);
  or _38649_ (_26834_[5], _07126_, _07110_);
  not _38650_ (_07127_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _38651_ (_07128_, _07025_, _07127_);
  and _38652_ (_07129_, _07025_, word_in[6]);
  nor _38653_ (_07131_, _07129_, _07128_);
  nor _38654_ (_07132_, _07131_, _07022_);
  and _38655_ (_07133_, _07022_, word_in[14]);
  or _38656_ (_07134_, _07133_, _07132_);
  and _38657_ (_07136_, _07134_, _07021_);
  and _38658_ (_07137_, _07019_, _06620_);
  or _38659_ (_07138_, _07137_, _07136_);
  and _38660_ (_07139_, _07138_, _07018_);
  and _38661_ (_07140_, _07017_, word_in[30]);
  or _38662_ (_26834_[6], _07140_, _07139_);
  and _38663_ (_07142_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _38664_ (_07143_, _06203_, _23887_);
  or _38665_ (_02081_, _07143_, _07142_);
  and _38666_ (_07144_, _07019_, _06047_);
  nor _38667_ (_07146_, _07025_, _05732_);
  and _38668_ (_07147_, _07025_, word_in[7]);
  nor _38669_ (_07148_, _07147_, _07146_);
  nor _38670_ (_07149_, _07148_, _07022_);
  and _38671_ (_07150_, _07022_, word_in[15]);
  or _38672_ (_07151_, _07150_, _07149_);
  and _38673_ (_07152_, _07151_, _07021_);
  or _38674_ (_07153_, _07152_, _07144_);
  and _38675_ (_07154_, _07153_, _07018_);
  and _38676_ (_07155_, _07017_, word_in[31]);
  or _38677_ (_26834_[7], _07155_, _07154_);
  and _38678_ (_07157_, _06129_, _24089_);
  and _38679_ (_07158_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or _38680_ (_02099_, _07158_, _07157_);
  and _38681_ (_07159_, _07013_, _23583_);
  and _38682_ (_07160_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or _38683_ (_02128_, _07160_, _07159_);
  and _38684_ (_07161_, _06043_, _06073_);
  not _38685_ (_07162_, _07161_);
  and _38686_ (_07163_, _06885_, _05784_);
  and _38687_ (_07165_, _07163_, _06538_);
  not _38688_ (_07166_, _07163_);
  and _38689_ (_07167_, _06653_, _05797_);
  and _38690_ (_07168_, _06657_, _05760_);
  and _38691_ (_07169_, _07168_, word_in[0]);
  not _38692_ (_07170_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _38693_ (_07171_, _07168_, _07170_);
  nor _38694_ (_07172_, _07171_, _07169_);
  nor _38695_ (_07173_, _07172_, _07167_);
  and _38696_ (_07174_, _07167_, word_in[8]);
  or _38697_ (_07175_, _07174_, _07173_);
  and _38698_ (_07176_, _07175_, _07166_);
  or _38699_ (_07178_, _07176_, _07165_);
  and _38700_ (_07179_, _07178_, _07162_);
  and _38701_ (_07181_, _07161_, word_in[24]);
  or _38702_ (_26835_[0], _07181_, _07179_);
  and _38703_ (_07182_, _07163_, _06391_);
  not _38704_ (_07183_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _38705_ (_07184_, _07168_, _07183_);
  and _38706_ (_07186_, _07168_, word_in[1]);
  nor _38707_ (_07187_, _07186_, _07184_);
  nor _38708_ (_07189_, _07187_, _07167_);
  and _38709_ (_07190_, _07167_, word_in[9]);
  or _38710_ (_07191_, _07190_, _07189_);
  and _38711_ (_07192_, _07191_, _07166_);
  or _38712_ (_07193_, _07192_, _07182_);
  and _38713_ (_07195_, _07193_, _07162_);
  and _38714_ (_07196_, _07161_, word_in[25]);
  or _38715_ (_26835_[1], _07196_, _07195_);
  and _38716_ (_07198_, _06763_, _23548_);
  and _38717_ (_07200_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _38718_ (_02151_, _07200_, _07198_);
  and _38719_ (_07202_, _07163_, _06572_);
  not _38720_ (_07203_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _38721_ (_07205_, _07168_, _07203_);
  and _38722_ (_07206_, _07168_, word_in[2]);
  nor _38723_ (_07207_, _07206_, _07205_);
  nor _38724_ (_07208_, _07207_, _07167_);
  and _38725_ (_07209_, _07167_, word_in[10]);
  or _38726_ (_07210_, _07209_, _07208_);
  and _38727_ (_07211_, _07210_, _07166_);
  or _38728_ (_07212_, _07211_, _07202_);
  and _38729_ (_07213_, _07212_, _07162_);
  and _38730_ (_07215_, _07161_, word_in[26]);
  or _38731_ (_26835_[2], _07215_, _07213_);
  and _38732_ (_07217_, _07163_, _06586_);
  not _38733_ (_07218_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _38734_ (_07219_, _07168_, _07218_);
  and _38735_ (_07220_, _07168_, word_in[3]);
  nor _38736_ (_07222_, _07220_, _07219_);
  nor _38737_ (_07224_, _07222_, _07167_);
  and _38738_ (_07225_, _07167_, word_in[11]);
  or _38739_ (_07227_, _07225_, _07224_);
  and _38740_ (_07228_, _07227_, _07166_);
  or _38741_ (_07229_, _07228_, _07217_);
  and _38742_ (_07230_, _07229_, _07162_);
  and _38743_ (_07231_, _07161_, word_in[27]);
  or _38744_ (_26835_[3], _07231_, _07230_);
  and _38745_ (_07233_, _07163_, _06591_);
  not _38746_ (_07234_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _38747_ (_07235_, _07168_, _07234_);
  and _38748_ (_07236_, _07168_, word_in[4]);
  nor _38749_ (_07237_, _07236_, _07235_);
  nor _38750_ (_07238_, _07237_, _07167_);
  and _38751_ (_07239_, _07167_, word_in[12]);
  or _38752_ (_07240_, _07239_, _07238_);
  and _38753_ (_07241_, _07240_, _07166_);
  or _38754_ (_07242_, _07241_, _07233_);
  and _38755_ (_07243_, _07242_, _07162_);
  and _38756_ (_07244_, _07161_, word_in[28]);
  or _38757_ (_26835_[4], _07244_, _07243_);
  and _38758_ (_07246_, _07163_, _06606_);
  not _38759_ (_07247_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _38760_ (_07248_, _07168_, _07247_);
  and _38761_ (_07249_, _07168_, word_in[5]);
  nor _38762_ (_07250_, _07249_, _07248_);
  nor _38763_ (_07252_, _07250_, _07167_);
  and _38764_ (_07253_, _07167_, word_in[13]);
  or _38765_ (_07254_, _07253_, _07252_);
  and _38766_ (_07255_, _07254_, _07166_);
  or _38767_ (_07256_, _07255_, _07246_);
  and _38768_ (_07257_, _07256_, _07162_);
  and _38769_ (_07258_, _07161_, word_in[29]);
  or _38770_ (_26835_[5], _07258_, _07257_);
  and _38771_ (_07259_, _07163_, _06620_);
  not _38772_ (_07260_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _38773_ (_07261_, _07168_, _07260_);
  and _38774_ (_07262_, _07168_, word_in[6]);
  nor _38775_ (_07263_, _07262_, _07261_);
  nor _38776_ (_07264_, _07263_, _07167_);
  and _38777_ (_07265_, _07167_, word_in[14]);
  or _38778_ (_07267_, _07265_, _07264_);
  and _38779_ (_07268_, _07267_, _07166_);
  or _38780_ (_07269_, _07268_, _07259_);
  and _38781_ (_07271_, _07269_, _07162_);
  and _38782_ (_07272_, _07161_, word_in[30]);
  or _38783_ (_26835_[6], _07272_, _07271_);
  and _38784_ (_07273_, _07163_, _06047_);
  nor _38785_ (_07274_, _07168_, _05862_);
  and _38786_ (_07275_, _07168_, word_in[7]);
  nor _38787_ (_07277_, _07275_, _07274_);
  nor _38788_ (_07278_, _07277_, _07167_);
  and _38789_ (_07279_, _07167_, word_in[15]);
  or _38790_ (_07280_, _07279_, _07278_);
  and _38791_ (_07281_, _07280_, _07166_);
  or _38792_ (_07282_, _07281_, _07273_);
  and _38793_ (_07283_, _07282_, _07162_);
  and _38794_ (_07284_, _07161_, word_in[31]);
  or _38795_ (_26835_[7], _07284_, _07283_);
  and _38796_ (_07285_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _38797_ (_07286_, _06203_, _23548_);
  or _38798_ (_02165_, _07286_, _07285_);
  and _38799_ (_07287_, _06043_, _06080_);
  and _38800_ (_07288_, _07287_, word_in[24]);
  and _38801_ (_07289_, _06885_, _05751_);
  and _38802_ (_07290_, _06029_, _05797_);
  and _38803_ (_07291_, _06893_, _06032_);
  and _38804_ (_07292_, _07291_, word_in[0]);
  not _38805_ (_07294_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _38806_ (_07295_, _07291_, _07294_);
  nor _38807_ (_07296_, _07295_, _07292_);
  nor _38808_ (_07298_, _07296_, _07290_);
  and _38809_ (_07299_, _07290_, word_in[8]);
  or _38810_ (_07301_, _07299_, _07298_);
  or _38811_ (_07302_, _07301_, _07289_);
  not _38812_ (_07303_, _07287_);
  not _38813_ (_07304_, _07289_);
  or _38814_ (_07305_, _07304_, _06538_);
  and _38815_ (_07307_, _07305_, _07303_);
  and _38816_ (_07308_, _07307_, _07302_);
  or _38817_ (_26836_[0], _07308_, _07288_);
  not _38818_ (_07310_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _38819_ (_07311_, _07291_, _07310_);
  and _38820_ (_07312_, _07291_, _06548_);
  or _38821_ (_07313_, _07312_, _07311_);
  or _38822_ (_07314_, _07313_, _07290_);
  not _38823_ (_07315_, _07290_);
  or _38824_ (_07316_, _07315_, word_in[9]);
  and _38825_ (_07318_, _07316_, _07314_);
  or _38826_ (_07319_, _07318_, _07289_);
  or _38827_ (_07320_, _07304_, _06391_);
  and _38828_ (_07321_, _07320_, _07303_);
  and _38829_ (_07322_, _07321_, _07319_);
  and _38830_ (_07323_, _07287_, word_in[25]);
  or _38831_ (_26836_[1], _07323_, _07322_);
  and _38832_ (_07325_, _07287_, word_in[26]);
  or _38833_ (_07326_, _07304_, _06572_);
  and _38834_ (_07327_, _07326_, _07303_);
  and _38835_ (_07328_, _07291_, word_in[2]);
  not _38836_ (_07329_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _38837_ (_07330_, _07291_, _07329_);
  nor _38838_ (_07331_, _07330_, _07328_);
  nor _38839_ (_07332_, _07331_, _07290_);
  and _38840_ (_07333_, _07290_, word_in[10]);
  or _38841_ (_07334_, _07333_, _07332_);
  or _38842_ (_07335_, _07334_, _07289_);
  and _38843_ (_07336_, _07335_, _07327_);
  or _38844_ (_26836_[2], _07336_, _07325_);
  and _38845_ (_07337_, _07287_, word_in[27]);
  not _38846_ (_07339_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _38847_ (_07340_, _07291_, _07339_);
  and _38848_ (_07342_, _07291_, _06427_);
  or _38849_ (_07343_, _07342_, _07340_);
  or _38850_ (_07345_, _07343_, _07290_);
  or _38851_ (_07347_, _07315_, word_in[11]);
  and _38852_ (_07348_, _07347_, _07345_);
  or _38853_ (_07350_, _07348_, _07289_);
  or _38854_ (_07351_, _07304_, _06586_);
  and _38855_ (_07352_, _07351_, _07303_);
  and _38856_ (_07354_, _07352_, _07350_);
  or _38857_ (_26836_[3], _07354_, _07337_);
  and _38858_ (_07356_, _07287_, word_in[28]);
  not _38859_ (_07357_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _38860_ (_07358_, _07291_, _07357_);
  and _38861_ (_07359_, _07291_, _06450_);
  or _38862_ (_07361_, _07359_, _07358_);
  or _38863_ (_07362_, _07361_, _07290_);
  or _38864_ (_07363_, _07315_, word_in[12]);
  and _38865_ (_07364_, _07363_, _07362_);
  or _38866_ (_07365_, _07364_, _07289_);
  or _38867_ (_07367_, _07304_, _06591_);
  and _38868_ (_07368_, _07367_, _07303_);
  and _38869_ (_07369_, _07368_, _07365_);
  or _38870_ (_26836_[4], _07369_, _07356_);
  and _38871_ (_07371_, _07287_, word_in[29]);
  or _38872_ (_07372_, _07304_, _06606_);
  and _38873_ (_07373_, _07372_, _07303_);
  and _38874_ (_07374_, _07291_, word_in[5]);
  not _38875_ (_07375_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _38876_ (_07376_, _07291_, _07375_);
  nor _38877_ (_07377_, _07376_, _07374_);
  nor _38878_ (_07378_, _07377_, _07290_);
  and _38879_ (_07379_, _07290_, word_in[13]);
  or _38880_ (_07380_, _07379_, _07378_);
  or _38881_ (_07381_, _07380_, _07289_);
  and _38882_ (_07382_, _07381_, _07373_);
  or _38883_ (_26836_[5], _07382_, _07371_);
  and _38884_ (_07383_, _07287_, word_in[30]);
  not _38885_ (_07384_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _38886_ (_07385_, _07291_, _07384_);
  and _38887_ (_07387_, _07291_, word_in[6]);
  nor _38888_ (_07388_, _07387_, _07385_);
  nor _38889_ (_07389_, _07388_, _07290_);
  and _38890_ (_07390_, _07290_, word_in[14]);
  or _38891_ (_07392_, _07390_, _07389_);
  and _38892_ (_07393_, _07392_, _07304_);
  and _38893_ (_07395_, _07289_, _06620_);
  or _38894_ (_07396_, _07395_, _07393_);
  and _38895_ (_07398_, _07396_, _07303_);
  or _38896_ (_26836_[6], _07398_, _07383_);
  nor _38897_ (_07400_, _07291_, _05726_);
  and _38898_ (_07401_, _07291_, _06496_);
  or _38899_ (_07402_, _07401_, _07400_);
  or _38900_ (_07404_, _07402_, _07290_);
  or _38901_ (_07405_, _07315_, word_in[15]);
  and _38902_ (_07406_, _07405_, _07404_);
  or _38903_ (_07408_, _07406_, _07289_);
  or _38904_ (_07410_, _07304_, _06047_);
  and _38905_ (_07411_, _07410_, _07303_);
  and _38906_ (_07412_, _07411_, _07408_);
  and _38907_ (_07413_, _07287_, word_in[31]);
  or _38908_ (_26836_[7], _07413_, _07412_);
  and _38909_ (_07415_, _07013_, _23887_);
  and _38910_ (_07416_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _38911_ (_02261_, _07416_, _07415_);
  and _38912_ (_07417_, _06043_, _05957_);
  and _38913_ (_07419_, _07417_, _05751_);
  not _38914_ (_07420_, _07419_);
  and _38915_ (_07421_, _06022_, _06105_);
  and _38916_ (_07422_, _07421_, word_in[16]);
  not _38917_ (_07423_, _07421_);
  and _38918_ (_07424_, _06028_, _05761_);
  not _38919_ (_07426_, _07424_);
  not _38920_ (_07428_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _38921_ (_07429_, _06033_, _05669_);
  and _38922_ (_07430_, _07429_, _06370_);
  nor _38923_ (_07431_, _07430_, _07428_);
  and _38924_ (_07432_, _07430_, word_in[0]);
  or _38925_ (_07434_, _07432_, _07431_);
  and _38926_ (_07435_, _07434_, _07426_);
  and _38927_ (_07436_, _07424_, word_in[8]);
  or _38928_ (_07437_, _07436_, _07435_);
  and _38929_ (_07438_, _07437_, _07423_);
  or _38930_ (_07439_, _07438_, _07422_);
  and _38931_ (_07440_, _07439_, _07420_);
  and _38932_ (_07441_, _07419_, word_in[24]);
  or _38933_ (_26837_[0], _07441_, _07440_);
  and _38934_ (_07442_, _07421_, word_in[17]);
  not _38935_ (_07443_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _38936_ (_07445_, _07430_, _07443_);
  and _38937_ (_07446_, _07430_, word_in[1]);
  or _38938_ (_07447_, _07446_, _07445_);
  and _38939_ (_07448_, _07447_, _07426_);
  and _38940_ (_07450_, _07424_, word_in[9]);
  or _38941_ (_07451_, _07450_, _07448_);
  and _38942_ (_07452_, _07451_, _07423_);
  or _38943_ (_07453_, _07452_, _07442_);
  and _38944_ (_07454_, _07453_, _07420_);
  and _38945_ (_07455_, _07419_, word_in[25]);
  or _38946_ (_26837_[1], _07455_, _07454_);
  and _38947_ (_07457_, _07421_, word_in[18]);
  not _38948_ (_07458_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _38949_ (_07459_, _07430_, _07458_);
  and _38950_ (_07460_, _07430_, word_in[2]);
  or _38951_ (_07461_, _07460_, _07459_);
  and _38952_ (_07463_, _07461_, _07426_);
  and _38953_ (_07464_, _07424_, word_in[10]);
  or _38954_ (_07465_, _07464_, _07463_);
  and _38955_ (_07466_, _07465_, _07423_);
  or _38956_ (_07467_, _07466_, _07457_);
  and _38957_ (_07468_, _07467_, _07420_);
  and _38958_ (_07470_, _07419_, word_in[26]);
  or _38959_ (_26837_[2], _07470_, _07468_);
  and _38960_ (_07472_, _07421_, word_in[19]);
  not _38961_ (_07473_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _38962_ (_07474_, _07430_, _07473_);
  and _38963_ (_07475_, _07430_, word_in[3]);
  or _38964_ (_07476_, _07475_, _07474_);
  and _38965_ (_07477_, _07476_, _07426_);
  and _38966_ (_07478_, _07424_, word_in[11]);
  or _38967_ (_07480_, _07478_, _07477_);
  and _38968_ (_07481_, _07480_, _07423_);
  or _38969_ (_07482_, _07481_, _07472_);
  and _38970_ (_07483_, _07482_, _07420_);
  and _38971_ (_07484_, _07419_, word_in[27]);
  or _38972_ (_26837_[3], _07484_, _07483_);
  and _38973_ (_07485_, _07421_, word_in[20]);
  not _38974_ (_07486_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _38975_ (_07487_, _07430_, _07486_);
  and _38976_ (_07488_, _07430_, word_in[4]);
  or _38977_ (_07489_, _07488_, _07487_);
  and _38978_ (_07490_, _07489_, _07426_);
  and _38979_ (_07491_, _07424_, word_in[12]);
  or _38980_ (_07492_, _07491_, _07490_);
  and _38981_ (_07493_, _07492_, _07423_);
  or _38982_ (_07494_, _07493_, _07485_);
  and _38983_ (_07495_, _07494_, _07420_);
  and _38984_ (_07496_, _07419_, word_in[28]);
  or _38985_ (_26837_[4], _07496_, _07495_);
  and _38986_ (_07497_, _07421_, word_in[21]);
  not _38987_ (_07498_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _38988_ (_07500_, _07430_, _07498_);
  and _38989_ (_07502_, _07430_, word_in[5]);
  or _38990_ (_07504_, _07502_, _07500_);
  and _38991_ (_07505_, _07504_, _07426_);
  and _38992_ (_07507_, _07424_, word_in[13]);
  or _38993_ (_07508_, _07507_, _07505_);
  and _38994_ (_07509_, _07508_, _07423_);
  or _38995_ (_07510_, _07509_, _07497_);
  and _38996_ (_07512_, _07510_, _07420_);
  and _38997_ (_07514_, _07419_, word_in[29]);
  or _38998_ (_26837_[5], _07514_, _07512_);
  and _38999_ (_07516_, _07421_, word_in[22]);
  not _39000_ (_07517_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _39001_ (_07518_, _07430_, _07517_);
  and _39002_ (_07519_, _07430_, word_in[6]);
  or _39003_ (_07520_, _07519_, _07518_);
  and _39004_ (_07521_, _07520_, _07426_);
  and _39005_ (_07522_, _07424_, word_in[14]);
  or _39006_ (_07523_, _07522_, _07521_);
  and _39007_ (_07524_, _07523_, _07423_);
  or _39008_ (_07525_, _07524_, _07516_);
  and _39009_ (_07526_, _07525_, _07420_);
  and _39010_ (_07527_, _07419_, word_in[30]);
  or _39011_ (_26837_[6], _07527_, _07526_);
  and _39012_ (_07529_, _07421_, word_in[23]);
  nor _39013_ (_07530_, _07430_, _05832_);
  and _39014_ (_07531_, _07430_, word_in[7]);
  or _39015_ (_07532_, _07531_, _07530_);
  and _39016_ (_07533_, _07532_, _07426_);
  and _39017_ (_07534_, _07424_, word_in[15]);
  or _39018_ (_07536_, _07534_, _07533_);
  and _39019_ (_07537_, _07536_, _07423_);
  or _39020_ (_07538_, _07537_, _07529_);
  and _39021_ (_07539_, _07538_, _07420_);
  and _39022_ (_07541_, _07419_, word_in[31]);
  or _39023_ (_26837_[7], _07541_, _07539_);
  and _39024_ (_07543_, _04920_, _23887_);
  and _39025_ (_07545_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _39026_ (_02327_, _07545_, _07543_);
  and _39027_ (_07547_, _24497_, _24219_);
  and _39028_ (_07548_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or _39029_ (_02342_, _07548_, _07547_);
  and _39030_ (_07549_, _06043_, _06105_);
  and _39031_ (_07551_, _06512_, _05885_);
  not _39032_ (_07552_, _07551_);
  or _39033_ (_07553_, _07552_, word_in[16]);
  and _39034_ (_07555_, _06515_, _05763_);
  not _39035_ (_07556_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _39036_ (_07557_, _07429_, _06521_);
  nor _39037_ (_07559_, _07557_, _07556_);
  and _39038_ (_07560_, _07557_, _06525_);
  or _39039_ (_07561_, _07560_, _07559_);
  or _39040_ (_07563_, _07561_, _07555_);
  not _39041_ (_07564_, _07555_);
  or _39042_ (_07566_, _07564_, word_in[8]);
  and _39043_ (_07567_, _07566_, _07563_);
  or _39044_ (_07568_, _07567_, _07551_);
  and _39045_ (_07569_, _07568_, _07553_);
  or _39046_ (_07570_, _07569_, _07549_);
  not _39047_ (_07571_, _07549_);
  or _39048_ (_07572_, _07571_, word_in[24]);
  and _39049_ (_26838_[0], _07572_, _07570_);
  not _39050_ (_07573_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _39051_ (_07574_, _07557_, _07573_);
  and _39052_ (_07575_, _07557_, _06548_);
  or _39053_ (_07576_, _07575_, _07574_);
  or _39054_ (_07578_, _07576_, _07555_);
  or _39055_ (_07579_, _07564_, word_in[9]);
  and _39056_ (_07581_, _07579_, _07578_);
  or _39057_ (_07582_, _07581_, _07551_);
  or _39058_ (_07583_, _07552_, word_in[17]);
  and _39059_ (_07584_, _07583_, _07571_);
  and _39060_ (_07585_, _07584_, _07582_);
  and _39061_ (_07587_, _07549_, word_in[25]);
  or _39062_ (_26838_[1], _07587_, _07585_);
  and _39063_ (_07589_, _07551_, word_in[18]);
  not _39064_ (_07590_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _39065_ (_07591_, _07557_, _07590_);
  and _39066_ (_07592_, _07557_, word_in[2]);
  nor _39067_ (_07593_, _07592_, _07591_);
  nor _39068_ (_07594_, _07593_, _07555_);
  and _39069_ (_07595_, _07555_, word_in[10]);
  or _39070_ (_07596_, _07595_, _07594_);
  and _39071_ (_07597_, _07596_, _07552_);
  or _39072_ (_07598_, _07597_, _07589_);
  and _39073_ (_07599_, _07598_, _07571_);
  and _39074_ (_07600_, _07549_, word_in[26]);
  or _39075_ (_26838_[2], _07600_, _07599_);
  and _39076_ (_07601_, _07551_, word_in[19]);
  not _39077_ (_07602_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _39078_ (_07604_, _07557_, _07602_);
  and _39079_ (_07605_, _07557_, word_in[3]);
  nor _39080_ (_07606_, _07605_, _07604_);
  nor _39081_ (_07608_, _07606_, _07555_);
  and _39082_ (_07609_, _07555_, word_in[11]);
  or _39083_ (_07610_, _07609_, _07608_);
  and _39084_ (_07611_, _07610_, _07552_);
  or _39085_ (_07612_, _07611_, _07601_);
  and _39086_ (_07613_, _07612_, _07571_);
  and _39087_ (_07615_, _07549_, word_in[27]);
  or _39088_ (_26838_[3], _07615_, _07613_);
  not _39089_ (_07616_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _39090_ (_07617_, _07557_, _07616_);
  and _39091_ (_07618_, _07557_, _06450_);
  or _39092_ (_07619_, _07618_, _07617_);
  or _39093_ (_07620_, _07619_, _07555_);
  or _39094_ (_07621_, _07564_, word_in[12]);
  and _39095_ (_07622_, _07621_, _07620_);
  or _39096_ (_07623_, _07622_, _07551_);
  or _39097_ (_07625_, _07552_, _06591_);
  and _39098_ (_07627_, _07625_, _07571_);
  and _39099_ (_07628_, _07627_, _07623_);
  and _39100_ (_07629_, _07549_, word_in[28]);
  or _39101_ (_26838_[4], _07629_, _07628_);
  or _39102_ (_07630_, _07552_, word_in[21]);
  not _39103_ (_07631_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _39104_ (_07632_, _07557_, _07631_);
  and _39105_ (_07633_, _07557_, _06469_);
  or _39106_ (_07634_, _07633_, _07632_);
  or _39107_ (_07635_, _07634_, _07555_);
  or _39108_ (_07636_, _07564_, word_in[13]);
  and _39109_ (_07637_, _07636_, _07635_);
  or _39110_ (_07638_, _07637_, _07551_);
  and _39111_ (_07640_, _07638_, _07630_);
  and _39112_ (_07641_, _07640_, _07571_);
  and _39113_ (_07642_, _07549_, word_in[29]);
  or _39114_ (_26838_[5], _07642_, _07641_);
  and _39115_ (_07643_, _07551_, word_in[22]);
  and _39116_ (_07644_, _07557_, word_in[6]);
  not _39117_ (_07647_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _39118_ (_07649_, _07557_, _07647_);
  nor _39119_ (_07650_, _07649_, _07644_);
  nor _39120_ (_07651_, _07650_, _07555_);
  and _39121_ (_07652_, _07555_, word_in[14]);
  or _39122_ (_07653_, _07652_, _07651_);
  and _39123_ (_07654_, _07653_, _07552_);
  or _39124_ (_07655_, _07654_, _07643_);
  and _39125_ (_07656_, _07655_, _07571_);
  and _39126_ (_07657_, _07549_, word_in[30]);
  or _39127_ (_26838_[6], _07657_, _07656_);
  nor _39128_ (_07658_, _07557_, _05709_);
  and _39129_ (_07659_, _07557_, _06496_);
  or _39130_ (_07660_, _07659_, _07658_);
  or _39131_ (_07661_, _07660_, _07555_);
  or _39132_ (_07662_, _07564_, word_in[15]);
  and _39133_ (_07663_, _07662_, _07661_);
  or _39134_ (_07664_, _07663_, _07551_);
  or _39135_ (_07665_, _07552_, _06047_);
  and _39136_ (_07666_, _07665_, _07571_);
  and _39137_ (_07667_, _07666_, _07664_);
  and _39138_ (_07668_, _07549_, word_in[31]);
  or _39139_ (_26838_[7], _07668_, _07667_);
  nor _39140_ (_26841_[2], _26684_, rst);
  and _39141_ (_07669_, _06647_, _05957_);
  and _39142_ (_07670_, _06649_, _05885_);
  not _39143_ (_07671_, _07670_);
  or _39144_ (_07672_, _07671_, _06538_);
  and _39145_ (_07673_, _06653_, _05763_);
  not _39146_ (_07674_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _39147_ (_07675_, _06657_, _05669_);
  nor _39148_ (_07676_, _07675_, _07674_);
  and _39149_ (_07677_, _07675_, word_in[0]);
  or _39150_ (_07678_, _07677_, _07676_);
  or _39151_ (_07679_, _07678_, _07673_);
  not _39152_ (_07680_, _07673_);
  or _39153_ (_07681_, _07680_, word_in[8]);
  and _39154_ (_07682_, _07681_, _07679_);
  or _39155_ (_07683_, _07682_, _07670_);
  and _39156_ (_07684_, _07683_, _07672_);
  or _39157_ (_07685_, _07684_, _07669_);
  not _39158_ (_07686_, _07669_);
  or _39159_ (_07687_, _07686_, word_in[24]);
  and _39160_ (_26824_[0], _07687_, _07685_);
  not _39161_ (_07688_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _39162_ (_07689_, _07675_, _07688_);
  and _39163_ (_07690_, _07675_, word_in[1]);
  or _39164_ (_07691_, _07690_, _07689_);
  or _39165_ (_07692_, _07691_, _07673_);
  or _39166_ (_07693_, _07680_, word_in[9]);
  and _39167_ (_07694_, _07693_, _07692_);
  or _39168_ (_07695_, _07694_, _07670_);
  or _39169_ (_07696_, _07671_, _06391_);
  and _39170_ (_07697_, _07696_, _07686_);
  and _39171_ (_07698_, _07697_, _07695_);
  and _39172_ (_07699_, _07669_, word_in[25]);
  or _39173_ (_26824_[1], _07699_, _07698_);
  not _39174_ (_07700_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _39175_ (_07701_, _07675_, _07700_);
  and _39176_ (_07702_, _07675_, word_in[2]);
  or _39177_ (_07704_, _07702_, _07701_);
  or _39178_ (_07705_, _07704_, _07673_);
  or _39179_ (_07706_, _07680_, word_in[10]);
  and _39180_ (_07707_, _07706_, _07705_);
  or _39181_ (_07708_, _07707_, _07670_);
  or _39182_ (_07709_, _07671_, _06572_);
  and _39183_ (_07710_, _07709_, _07686_);
  and _39184_ (_07711_, _07710_, _07708_);
  and _39185_ (_07712_, _07669_, word_in[26]);
  or _39186_ (_26824_[2], _07712_, _07711_);
  or _39187_ (_07713_, _07671_, _06586_);
  not _39188_ (_07714_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _39189_ (_07715_, _07675_, _07714_);
  and _39190_ (_07716_, _07675_, word_in[3]);
  or _39191_ (_07717_, _07716_, _07715_);
  or _39192_ (_07718_, _07717_, _07673_);
  or _39193_ (_07719_, _07680_, word_in[11]);
  and _39194_ (_07720_, _07719_, _07718_);
  or _39195_ (_07721_, _07720_, _07670_);
  and _39196_ (_07722_, _07721_, _07713_);
  or _39197_ (_07724_, _07722_, _07669_);
  or _39198_ (_07725_, _07686_, word_in[27]);
  and _39199_ (_26824_[3], _07725_, _07724_);
  not _39200_ (_07726_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _39201_ (_07727_, _07675_, _07726_);
  and _39202_ (_07728_, _07675_, word_in[4]);
  or _39203_ (_07729_, _07728_, _07727_);
  or _39204_ (_07730_, _07729_, _07673_);
  or _39205_ (_07731_, _07680_, word_in[12]);
  and _39206_ (_07732_, _07731_, _07730_);
  or _39207_ (_07733_, _07732_, _07670_);
  or _39208_ (_07734_, _07671_, _06591_);
  and _39209_ (_07735_, _07734_, _07686_);
  and _39210_ (_07736_, _07735_, _07733_);
  and _39211_ (_07737_, _07669_, word_in[28]);
  or _39212_ (_26824_[4], _07737_, _07736_);
  not _39213_ (_07738_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _39214_ (_07739_, _07675_, _07738_);
  and _39215_ (_07740_, _07675_, word_in[5]);
  or _39216_ (_07741_, _07740_, _07739_);
  or _39217_ (_07743_, _07741_, _07673_);
  or _39218_ (_07744_, _07680_, word_in[13]);
  and _39219_ (_07745_, _07744_, _07743_);
  or _39220_ (_07746_, _07745_, _07670_);
  or _39221_ (_07747_, _07671_, _06606_);
  and _39222_ (_07748_, _07747_, _07686_);
  and _39223_ (_07749_, _07748_, _07746_);
  and _39224_ (_07750_, _07669_, word_in[29]);
  or _39225_ (_26824_[5], _07750_, _07749_);
  or _39226_ (_07751_, _07671_, _06620_);
  not _39227_ (_07752_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _39228_ (_07753_, _07675_, _07752_);
  and _39229_ (_07754_, _07675_, word_in[6]);
  or _39230_ (_07755_, _07754_, _07753_);
  or _39231_ (_07756_, _07755_, _07673_);
  or _39232_ (_07757_, _07680_, word_in[14]);
  and _39233_ (_07758_, _07757_, _07756_);
  or _39234_ (_07759_, _07758_, _07670_);
  and _39235_ (_07760_, _07759_, _07751_);
  or _39236_ (_07761_, _07760_, _07669_);
  or _39237_ (_07763_, _07686_, word_in[30]);
  and _39238_ (_26824_[6], _07763_, _07761_);
  nor _39239_ (_07764_, _07675_, _05827_);
  and _39240_ (_07765_, _07675_, word_in[7]);
  or _39241_ (_07766_, _07765_, _07764_);
  or _39242_ (_07767_, _07766_, _07673_);
  or _39243_ (_07768_, _07680_, word_in[15]);
  and _39244_ (_07769_, _07768_, _07767_);
  or _39245_ (_07770_, _07769_, _07670_);
  or _39246_ (_07771_, _07671_, _06047_);
  and _39247_ (_07772_, _07771_, _07686_);
  and _39248_ (_07773_, _07772_, _07770_);
  and _39249_ (_07774_, _07669_, word_in[31]);
  or _39250_ (_26824_[7], _07774_, _07773_);
  and _39251_ (_07775_, _25414_, _23887_);
  and _39252_ (_07776_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _39253_ (_02454_, _07776_, _07775_);
  and _39254_ (_07777_, _25414_, _24219_);
  and _39255_ (_07778_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or _39256_ (_02457_, _07778_, _07777_);
  and _39257_ (_07779_, _25413_, _24140_);
  and _39258_ (_07780_, _07779_, _23996_);
  not _39259_ (_07781_, _07779_);
  and _39260_ (_07782_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or _39261_ (_27158_, _07782_, _07780_);
  and _39262_ (_07783_, _07779_, _23583_);
  and _39263_ (_07784_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  or _39264_ (_02464_, _07784_, _07783_);
  and _39265_ (_07785_, _07779_, _23548_);
  and _39266_ (_07786_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or _39267_ (_02466_, _07786_, _07785_);
  and _39268_ (_07787_, _02368_, _24089_);
  and _39269_ (_07788_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or _39270_ (_27151_, _07788_, _07787_);
  and _39271_ (_07789_, _02368_, _23887_);
  and _39272_ (_07790_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or _39273_ (_02477_, _07790_, _07789_);
  and _39274_ (_07791_, _02413_, _24051_);
  and _39275_ (_07792_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _39276_ (_02482_, _07792_, _07791_);
  and _39277_ (_07793_, _06767_, _05885_);
  and _39278_ (_07794_, _06029_, _05763_);
  not _39279_ (_07795_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _39280_ (_07796_, _07429_, _06032_);
  nor _39281_ (_07797_, _07796_, _07795_);
  and _39282_ (_07798_, _07796_, _06525_);
  or _39283_ (_07799_, _07798_, _07797_);
  or _39284_ (_07800_, _07799_, _07794_);
  not _39285_ (_07801_, word_in[8]);
  nand _39286_ (_07802_, _07794_, _07801_);
  and _39287_ (_07803_, _07802_, _07800_);
  or _39288_ (_07804_, _07803_, _07793_);
  and _39289_ (_07805_, _06044_, _05957_);
  not _39290_ (_07806_, _07805_);
  not _39291_ (_07807_, _07793_);
  or _39292_ (_07808_, _07807_, word_in[16]);
  and _39293_ (_07809_, _07808_, _07806_);
  and _39294_ (_07810_, _07809_, _07804_);
  and _39295_ (_07811_, _07805_, _06364_);
  or _39296_ (_26825_[0], _07811_, _07810_);
  and _39297_ (_07813_, _02413_, _23583_);
  and _39298_ (_07814_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _39299_ (_02487_, _07814_, _07813_);
  and _39300_ (_07815_, _07796_, word_in[1]);
  not _39301_ (_07816_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _39302_ (_07817_, _07796_, _07816_);
  nor _39303_ (_07818_, _07817_, _07815_);
  nor _39304_ (_07819_, _07818_, _07794_);
  and _39305_ (_07820_, _07794_, word_in[9]);
  or _39306_ (_07821_, _07820_, _07819_);
  and _39307_ (_07822_, _07821_, _07807_);
  and _39308_ (_07823_, _07793_, word_in[17]);
  or _39309_ (_07824_, _07823_, _07805_);
  or _39310_ (_07825_, _07824_, _07822_);
  or _39311_ (_07826_, _07806_, _06801_);
  and _39312_ (_26825_[1], _07826_, _07825_);
  and _39313_ (_07827_, _07796_, word_in[2]);
  not _39314_ (_07828_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _39315_ (_07829_, _07796_, _07828_);
  nor _39316_ (_07830_, _07829_, _07827_);
  nor _39317_ (_07831_, _07830_, _07794_);
  and _39318_ (_07832_, _07794_, word_in[10]);
  or _39319_ (_07833_, _07832_, _07831_);
  and _39320_ (_07834_, _07833_, _07807_);
  and _39321_ (_07835_, _07793_, word_in[18]);
  or _39322_ (_07836_, _07835_, _07805_);
  or _39323_ (_07837_, _07836_, _07834_);
  or _39324_ (_07838_, _07806_, _06407_);
  and _39325_ (_26825_[2], _07838_, _07837_);
  and _39326_ (_07839_, _07796_, word_in[3]);
  not _39327_ (_07840_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _39328_ (_07841_, _07796_, _07840_);
  nor _39329_ (_07842_, _07841_, _07839_);
  nor _39330_ (_07843_, _07842_, _07794_);
  and _39331_ (_07844_, _07794_, word_in[11]);
  or _39332_ (_07845_, _07844_, _07843_);
  and _39333_ (_07846_, _07845_, _07807_);
  and _39334_ (_07847_, _07793_, word_in[19]);
  or _39335_ (_07848_, _07847_, _07846_);
  and _39336_ (_07849_, _07848_, _07806_);
  and _39337_ (_07850_, _07805_, word_in[27]);
  or _39338_ (_26825_[3], _07850_, _07849_);
  and _39339_ (_07851_, _02455_, _24051_);
  and _39340_ (_07852_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _39341_ (_02493_, _07852_, _07851_);
  and _39342_ (_07853_, _07796_, word_in[4]);
  not _39343_ (_07854_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _39344_ (_07855_, _07796_, _07854_);
  nor _39345_ (_07856_, _07855_, _07853_);
  nor _39346_ (_07857_, _07856_, _07794_);
  and _39347_ (_07858_, _07794_, word_in[12]);
  or _39348_ (_07859_, _07858_, _07857_);
  and _39349_ (_07860_, _07859_, _07807_);
  and _39350_ (_07861_, _07793_, _06591_);
  or _39351_ (_07862_, _07861_, _07860_);
  and _39352_ (_07863_, _07862_, _07806_);
  and _39353_ (_07864_, _07805_, word_in[28]);
  or _39354_ (_26825_[4], _07864_, _07863_);
  and _39355_ (_07865_, _02455_, _23583_);
  and _39356_ (_07866_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _39357_ (_02496_, _07866_, _07865_);
  and _39358_ (_07867_, _07796_, word_in[5]);
  not _39359_ (_07869_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _39360_ (_07871_, _07796_, _07869_);
  nor _39361_ (_07872_, _07871_, _07867_);
  nor _39362_ (_07873_, _07872_, _07794_);
  and _39363_ (_07874_, _07794_, word_in[13]);
  or _39364_ (_07876_, _07874_, _07873_);
  and _39365_ (_07878_, _07876_, _07807_);
  and _39366_ (_07880_, _07793_, word_in[21]);
  or _39367_ (_07882_, _07880_, _07805_);
  or _39368_ (_07883_, _07882_, _07878_);
  or _39369_ (_07885_, _07806_, _06463_);
  and _39370_ (_26825_[5], _07885_, _07883_);
  and _39371_ (_07886_, _07796_, word_in[6]);
  not _39372_ (_07887_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _39373_ (_07888_, _07796_, _07887_);
  nor _39374_ (_07890_, _07888_, _07886_);
  nor _39375_ (_07892_, _07890_, _07794_);
  and _39376_ (_07893_, _07794_, word_in[14]);
  or _39377_ (_07895_, _07893_, _07892_);
  and _39378_ (_07897_, _07895_, _07807_);
  and _39379_ (_07899_, _07793_, word_in[22]);
  or _39380_ (_07900_, _07899_, _07805_);
  or _39381_ (_07901_, _07900_, _07897_);
  or _39382_ (_07903_, _07806_, _06867_);
  and _39383_ (_26825_[6], _07903_, _07901_);
  and _39384_ (_07906_, _07796_, word_in[7]);
  nor _39385_ (_07907_, _07796_, _05697_);
  nor _39386_ (_07909_, _07907_, _07906_);
  nor _39387_ (_07911_, _07909_, _07794_);
  and _39388_ (_07913_, _07794_, word_in[15]);
  or _39389_ (_07915_, _07913_, _07911_);
  and _39390_ (_07916_, _07915_, _07807_);
  and _39391_ (_07918_, _07793_, _06047_);
  or _39392_ (_07919_, _07918_, _07916_);
  and _39393_ (_07920_, _07919_, _07806_);
  and _39394_ (_07921_, _07805_, word_in[31]);
  or _39395_ (_26825_[7], _07921_, _07920_);
  and _39396_ (_07922_, _02517_, _24134_);
  and _39397_ (_07924_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or _39398_ (_02506_, _07924_, _07922_);
  and _39399_ (_07925_, _02517_, _24089_);
  and _39400_ (_07926_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or _39401_ (_02510_, _07926_, _07925_);
  and _39402_ (_07927_, _02890_, _23583_);
  and _39403_ (_07928_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or _39404_ (_02529_, _07928_, _07927_);
  and _39405_ (_07929_, _04865_, _23996_);
  and _39406_ (_07930_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or _39407_ (_02533_, _07930_, _07929_);
  and _39408_ (_07931_, _04812_, _24089_);
  and _39409_ (_07932_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _39410_ (_02538_, _07932_, _07931_);
  and _39411_ (_07933_, _05431_, _23887_);
  and _39412_ (_07934_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or _39413_ (_27129_, _07934_, _07933_);
  and _39414_ (_07935_, _05431_, _24219_);
  and _39415_ (_07936_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or _39416_ (_02547_, _07936_, _07935_);
  and _39417_ (_07937_, _05456_, _23996_);
  and _39418_ (_07938_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _39419_ (_27128_, _07938_, _07937_);
  and _39420_ (_07939_, _03360_, _23996_);
  and _39421_ (_07940_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _39422_ (_02554_, _07940_, _07939_);
  and _39423_ (_07941_, _05456_, _23583_);
  and _39424_ (_07942_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _39425_ (_27125_, _07942_, _07941_);
  and _39426_ (_07943_, _05456_, _23548_);
  and _39427_ (_07945_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _39428_ (_02559_, _07945_, _07943_);
  and _39429_ (_07946_, _06024_, _05906_);
  not _39430_ (_07947_, _07946_);
  and _39431_ (_07948_, _06028_, _06221_);
  not _39432_ (_07949_, _07948_);
  not _39433_ (_07950_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _39434_ (_07951_, _06370_, _06034_);
  nor _39435_ (_07953_, _07951_, _07950_);
  and _39436_ (_07954_, _07951_, word_in[0]);
  or _39437_ (_07955_, _07954_, _07953_);
  and _39438_ (_07956_, _07955_, _07949_);
  and _39439_ (_07957_, _07948_, word_in[8]);
  or _39440_ (_07958_, _07957_, _07956_);
  and _39441_ (_07960_, _07958_, _07947_);
  and _39442_ (_07962_, _06043_, _06008_);
  and _39443_ (_07963_, _07962_, _05751_);
  and _39444_ (_07964_, _07946_, _06538_);
  or _39445_ (_07966_, _07964_, _07963_);
  or _39446_ (_07967_, _07966_, _07960_);
  not _39447_ (_07969_, _07963_);
  or _39448_ (_07970_, _07969_, _06364_);
  and _39449_ (_26826_[0], _07970_, _07967_);
  and _39450_ (_07971_, _05491_, _24051_);
  and _39451_ (_07973_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or _39452_ (_02567_, _07973_, _07971_);
  not _39453_ (_07974_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _39454_ (_07976_, _07951_, _07974_);
  and _39455_ (_07977_, _07951_, word_in[1]);
  or _39456_ (_07978_, _07977_, _07976_);
  or _39457_ (_07979_, _07978_, _07948_);
  or _39458_ (_07980_, _07949_, word_in[9]);
  and _39459_ (_07982_, _07980_, _07979_);
  or _39460_ (_07984_, _07982_, _07946_);
  or _39461_ (_07985_, _07947_, _06391_);
  and _39462_ (_07986_, _07985_, _07984_);
  or _39463_ (_07987_, _07986_, _07963_);
  or _39464_ (_07989_, _07969_, _06801_);
  and _39465_ (_26826_[1], _07989_, _07987_);
  and _39466_ (_07991_, _07946_, _06572_);
  not _39467_ (_07992_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _39468_ (_07994_, _07951_, _07992_);
  and _39469_ (_07996_, _07951_, word_in[2]);
  or _39470_ (_07998_, _07996_, _07994_);
  and _39471_ (_07999_, _07998_, _07949_);
  and _39472_ (_08000_, _07948_, word_in[10]);
  or _39473_ (_08001_, _08000_, _07999_);
  and _39474_ (_08003_, _08001_, _07947_);
  or _39475_ (_08004_, _08003_, _07991_);
  and _39476_ (_08006_, _08004_, _07969_);
  and _39477_ (_08007_, _07963_, _06407_);
  or _39478_ (_26826_[2], _08007_, _08006_);
  not _39479_ (_08008_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _39480_ (_08009_, _07951_, _08008_);
  and _39481_ (_08010_, _07951_, word_in[3]);
  or _39482_ (_08011_, _08010_, _08009_);
  or _39483_ (_08013_, _08011_, _07948_);
  or _39484_ (_08014_, _07949_, word_in[11]);
  and _39485_ (_08015_, _08014_, _08013_);
  and _39486_ (_08016_, _08015_, _07947_);
  and _39487_ (_08018_, _07946_, _06586_);
  or _39488_ (_08019_, _08018_, _07963_);
  or _39489_ (_08021_, _08019_, _08016_);
  or _39490_ (_08022_, _07969_, _06441_);
  and _39491_ (_26826_[3], _08022_, _08021_);
  and _39492_ (_08024_, _05491_, _24219_);
  and _39493_ (_08025_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or _39494_ (_02575_, _08025_, _08024_);
  not _39495_ (_08026_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _39496_ (_08027_, _07951_, _08026_);
  and _39497_ (_08028_, _07951_, word_in[4]);
  or _39498_ (_08029_, _08028_, _08027_);
  and _39499_ (_08030_, _08029_, _07949_);
  and _39500_ (_08031_, _07948_, word_in[12]);
  or _39501_ (_08032_, _08031_, _08030_);
  and _39502_ (_08033_, _08032_, _07947_);
  and _39503_ (_08034_, _07946_, _06591_);
  or _39504_ (_08035_, _08034_, _07963_);
  or _39505_ (_08036_, _08035_, _08033_);
  or _39506_ (_08037_, _07969_, _06446_);
  and _39507_ (_26826_[4], _08037_, _08036_);
  and _39508_ (_08038_, _24409_, _24134_);
  and _39509_ (_08039_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or _39510_ (_02579_, _08039_, _08038_);
  not _39511_ (_08040_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _39512_ (_08041_, _07951_, _08040_);
  and _39513_ (_08042_, _07951_, word_in[5]);
  or _39514_ (_08043_, _08042_, _08041_);
  or _39515_ (_08044_, _08043_, _07948_);
  or _39516_ (_08045_, _07949_, word_in[13]);
  and _39517_ (_08046_, _08045_, _08044_);
  and _39518_ (_08047_, _08046_, _07947_);
  and _39519_ (_08048_, _07946_, _06606_);
  or _39520_ (_08049_, _08048_, _07963_);
  or _39521_ (_08050_, _08049_, _08047_);
  or _39522_ (_08051_, _07969_, _06463_);
  and _39523_ (_26826_[5], _08051_, _08050_);
  not _39524_ (_08052_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _39525_ (_08053_, _07951_, _08052_);
  and _39526_ (_08054_, _07951_, word_in[6]);
  or _39527_ (_08055_, _08054_, _08053_);
  or _39528_ (_08056_, _08055_, _07948_);
  or _39529_ (_08057_, _07949_, word_in[14]);
  and _39530_ (_08058_, _08057_, _08056_);
  and _39531_ (_08059_, _08058_, _07947_);
  and _39532_ (_08060_, _07946_, _06620_);
  or _39533_ (_08061_, _08060_, _07963_);
  or _39534_ (_08062_, _08061_, _08059_);
  or _39535_ (_08063_, _07969_, _06867_);
  and _39536_ (_26826_[6], _08063_, _08062_);
  nor _39537_ (_08064_, _07951_, _05818_);
  and _39538_ (_08065_, _07951_, word_in[7]);
  or _39539_ (_08066_, _08065_, _08064_);
  and _39540_ (_08067_, _08066_, _07949_);
  and _39541_ (_08068_, _07948_, word_in[15]);
  or _39542_ (_08069_, _08068_, _08067_);
  and _39543_ (_08070_, _08069_, _07947_);
  and _39544_ (_08071_, _07946_, _06047_);
  or _39545_ (_08072_, _08071_, _07963_);
  or _39546_ (_08073_, _08072_, _08070_);
  or _39547_ (_08074_, _07969_, _06052_);
  and _39548_ (_26826_[7], _08074_, _08073_);
  not _39549_ (_08075_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _39550_ (_08076_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _08075_);
  and _39551_ (_26885_, _08076_, _22731_);
  and _39552_ (_08077_, _24409_, _23548_);
  and _39553_ (_08078_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or _39554_ (_27119_, _08078_, _08077_);
  and _39555_ (_08079_, _05485_, _24089_);
  and _39556_ (_08080_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _39557_ (_27135_, _08080_, _08079_);
  and _39558_ (_08081_, _05485_, _24219_);
  and _39559_ (_08082_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _39560_ (_27133_, _08082_, _08081_);
  and _39561_ (_08083_, _05431_, _23996_);
  and _39562_ (_08084_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or _39563_ (_27132_, _08084_, _08083_);
  and _39564_ (_08085_, _05485_, _23887_);
  and _39565_ (_08086_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _39566_ (_27134_, _08086_, _08085_);
  and _39567_ (_08088_, _25414_, _24089_);
  and _39568_ (_08089_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _39569_ (_27160_, _08089_, _08088_);
  and _39570_ (_08090_, _07779_, _24051_);
  and _39571_ (_08091_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or _39572_ (_27157_, _08091_, _08090_);
  and _39573_ (_08092_, _02368_, _24134_);
  and _39574_ (_08093_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or _39575_ (_27153_, _08093_, _08092_);
  and _39576_ (_08094_, _02413_, _23996_);
  and _39577_ (_08095_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _39578_ (_27150_, _08095_, _08094_);
  and _39579_ (_08096_, _02455_, _23996_);
  and _39580_ (_08097_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _39581_ (_27146_, _08097_, _08096_);
  and _39582_ (_08098_, _06024_, _05753_);
  not _39583_ (_08099_, _08098_);
  and _39584_ (_08100_, _06515_, _05800_);
  and _39585_ (_08101_, _06521_, _06034_);
  and _39586_ (_08102_, _08101_, word_in[0]);
  not _39587_ (_08104_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _39588_ (_08105_, _08101_, _08104_);
  nor _39589_ (_08106_, _08105_, _08102_);
  nor _39590_ (_08107_, _08106_, _08100_);
  and _39591_ (_08108_, _08100_, word_in[8]);
  or _39592_ (_08109_, _08108_, _08107_);
  and _39593_ (_08110_, _08109_, _08099_);
  and _39594_ (_08111_, _07962_, _05906_);
  and _39595_ (_08112_, _08098_, _06538_);
  or _39596_ (_08113_, _08112_, _08111_);
  or _39597_ (_08114_, _08113_, _08110_);
  not _39598_ (_08115_, _08111_);
  or _39599_ (_08116_, _08115_, _06364_);
  and _39600_ (_26827_[0], _08116_, _08114_);
  not _39601_ (_08117_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _39602_ (_08118_, _08101_, _08117_);
  and _39603_ (_08119_, _08101_, _06548_);
  or _39604_ (_08120_, _08119_, _08118_);
  or _39605_ (_08121_, _08120_, _08100_);
  not _39606_ (_08122_, _08100_);
  or _39607_ (_08124_, _08122_, word_in[9]);
  and _39608_ (_08125_, _08124_, _08121_);
  or _39609_ (_08126_, _08125_, _08098_);
  or _39610_ (_08127_, _08099_, _06391_);
  and _39611_ (_08128_, _08127_, _08115_);
  and _39612_ (_08129_, _08128_, _08126_);
  and _39613_ (_08130_, _08111_, _06801_);
  or _39614_ (_26827_[1], _08130_, _08129_);
  and _39615_ (_08131_, _02517_, _24219_);
  and _39616_ (_08132_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or _39617_ (_27142_, _08132_, _08131_);
  and _39618_ (_08133_, _08101_, word_in[2]);
  not _39619_ (_08134_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _39620_ (_08135_, _08101_, _08134_);
  nor _39621_ (_08136_, _08135_, _08133_);
  nor _39622_ (_08137_, _08136_, _08100_);
  and _39623_ (_08138_, _08100_, word_in[10]);
  or _39624_ (_08139_, _08138_, _08137_);
  and _39625_ (_08140_, _08139_, _08099_);
  and _39626_ (_08141_, _08098_, _06572_);
  or _39627_ (_08143_, _08141_, _08111_);
  or _39628_ (_08144_, _08143_, _08140_);
  or _39629_ (_08145_, _08115_, _06407_);
  and _39630_ (_26827_[2], _08145_, _08144_);
  and _39631_ (_08146_, _02890_, _24051_);
  and _39632_ (_08147_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or _39633_ (_27141_, _08147_, _08146_);
  not _39634_ (_08148_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _39635_ (_08149_, _08101_, _08148_);
  and _39636_ (_08150_, _08101_, _06427_);
  or _39637_ (_08151_, _08150_, _08149_);
  or _39638_ (_08152_, _08151_, _08100_);
  or _39639_ (_08153_, _08122_, word_in[11]);
  and _39640_ (_08154_, _08153_, _08152_);
  or _39641_ (_08155_, _08154_, _08098_);
  or _39642_ (_08156_, _08099_, _06586_);
  and _39643_ (_08157_, _08156_, _08115_);
  and _39644_ (_08158_, _08157_, _08155_);
  and _39645_ (_08159_, _08111_, _06441_);
  or _39646_ (_26827_[3], _08159_, _08158_);
  and _39647_ (_08160_, _02890_, _23548_);
  and _39648_ (_08161_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or _39649_ (_27140_, _08161_, _08160_);
  not _39650_ (_08162_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _39651_ (_08163_, _08101_, _08162_);
  and _39652_ (_08164_, _08101_, _06450_);
  or _39653_ (_08165_, _08164_, _08163_);
  or _39654_ (_08166_, _08165_, _08100_);
  or _39655_ (_08167_, _08122_, word_in[12]);
  and _39656_ (_08168_, _08167_, _08166_);
  or _39657_ (_08170_, _08168_, _08098_);
  or _39658_ (_08171_, _08099_, _06591_);
  and _39659_ (_08172_, _08171_, _08115_);
  and _39660_ (_08173_, _08172_, _08170_);
  and _39661_ (_08174_, _08111_, _06446_);
  or _39662_ (_26827_[4], _08174_, _08173_);
  and _39663_ (_08175_, _04812_, _24134_);
  and _39664_ (_08176_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _39665_ (_27139_, _08176_, _08175_);
  and _39666_ (_08177_, _08098_, _06606_);
  and _39667_ (_08178_, _08101_, word_in[5]);
  not _39668_ (_08179_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _39669_ (_08180_, _08101_, _08179_);
  nor _39670_ (_08181_, _08180_, _08178_);
  nor _39671_ (_08182_, _08181_, _08100_);
  and _39672_ (_08183_, _08100_, word_in[13]);
  or _39673_ (_08184_, _08183_, _08182_);
  and _39674_ (_08185_, _08184_, _08099_);
  or _39675_ (_08186_, _08185_, _08177_);
  and _39676_ (_08187_, _08186_, _08115_);
  and _39677_ (_08188_, _08111_, _06463_);
  or _39678_ (_26827_[5], _08188_, _08187_);
  and _39679_ (_08189_, _05431_, _24089_);
  and _39680_ (_08190_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or _39681_ (_27130_, _08190_, _08189_);
  and _39682_ (_08191_, _08101_, word_in[6]);
  not _39683_ (_08192_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _39684_ (_08193_, _08101_, _08192_);
  nor _39685_ (_08194_, _08193_, _08191_);
  nor _39686_ (_08195_, _08194_, _08100_);
  and _39687_ (_08196_, _08100_, word_in[14]);
  or _39688_ (_08197_, _08196_, _08195_);
  and _39689_ (_08198_, _08197_, _08099_);
  and _39690_ (_08199_, _08098_, _06620_);
  or _39691_ (_08200_, _08199_, _08111_);
  or _39692_ (_08201_, _08200_, _08198_);
  or _39693_ (_08202_, _08115_, _06867_);
  and _39694_ (_26827_[6], _08202_, _08201_);
  nor _39695_ (_08203_, _08101_, _05704_);
  and _39696_ (_08204_, _08101_, _06496_);
  or _39697_ (_08205_, _08204_, _08203_);
  or _39698_ (_08206_, _08205_, _08100_);
  or _39699_ (_08207_, _08122_, word_in[15]);
  and _39700_ (_08208_, _08207_, _08206_);
  or _39701_ (_08209_, _08208_, _08098_);
  or _39702_ (_08210_, _08099_, _06047_);
  and _39703_ (_08211_, _08210_, _08115_);
  and _39704_ (_08212_, _08211_, _08209_);
  and _39705_ (_08213_, _08111_, _06052_);
  or _39706_ (_26827_[7], _08213_, _08212_);
  and _39707_ (_08214_, _05456_, _24051_);
  and _39708_ (_08215_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _39709_ (_27127_, _08215_, _08214_);
  nand _39710_ (_08216_, _01816_, _24126_);
  and _39711_ (_08217_, _02210_, _02320_);
  and _39712_ (_08218_, _08217_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _39713_ (_08219_, _08218_);
  nor _39714_ (_08220_, _08219_, _01814_);
  not _39715_ (_08221_, _08220_);
  nor _39716_ (_08222_, _08221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _39717_ (_08223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _39718_ (_08224_, _08223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _39719_ (_08225_, _08224_, _02210_);
  and _39720_ (_08226_, _08225_, _02196_);
  nand _39721_ (_08227_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _39722_ (_08228_, _08227_, _01814_);
  and _39723_ (_08229_, _08221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _39724_ (_08230_, _08229_, _08228_);
  or _39725_ (_08231_, _08230_, _08222_);
  or _39726_ (_08232_, _08231_, _01816_);
  and _39727_ (_08234_, _08232_, _22731_);
  and _39728_ (_02667_, _08234_, _08216_);
  and _39729_ (_08235_, _05491_, _23887_);
  and _39730_ (_08236_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or _39731_ (_27123_, _08236_, _08235_);
  and _39732_ (_08239_, _24350_, _23887_);
  and _39733_ (_08241_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _39734_ (_27058_, _08241_, _08239_);
  and _39735_ (_08243_, _24409_, _23583_);
  and _39736_ (_08244_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or _39737_ (_27120_, _08244_, _08243_);
  and _39738_ (_08245_, _04812_, _23548_);
  and _39739_ (_08246_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _39740_ (_27137_, _08246_, _08245_);
  and _39741_ (_08248_, _05485_, _24134_);
  and _39742_ (_08250_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _39743_ (_27136_, _08250_, _08248_);
  and _39744_ (_08251_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and _39745_ (_08252_, _04897_, _23887_);
  or _39746_ (_27008_, _08252_, _08251_);
  and _39747_ (_08254_, _02455_, _24219_);
  and _39748_ (_08255_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _39749_ (_27144_, _08255_, _08254_);
  and _39750_ (_08257_, _06024_, _05784_);
  not _39751_ (_08258_, _08257_);
  and _39752_ (_08260_, _06653_, _05800_);
  and _39753_ (_08262_, _06657_, _05962_);
  and _39754_ (_08263_, _08262_, word_in[0]);
  not _39755_ (_08264_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _39756_ (_08265_, _08262_, _08264_);
  nor _39757_ (_08267_, _08265_, _08263_);
  nor _39758_ (_08269_, _08267_, _08260_);
  and _39759_ (_08271_, _08260_, word_in[8]);
  or _39760_ (_08273_, _08271_, _08269_);
  and _39761_ (_08274_, _08273_, _08258_);
  and _39762_ (_08276_, _06647_, _06008_);
  and _39763_ (_08277_, _08257_, _06538_);
  or _39764_ (_08279_, _08277_, _08276_);
  or _39765_ (_08281_, _08279_, _08274_);
  not _39766_ (_08282_, _08276_);
  or _39767_ (_08283_, _08282_, _06364_);
  and _39768_ (_26828_[0], _08283_, _08281_);
  and _39769_ (_08285_, _05491_, _24134_);
  and _39770_ (_08286_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or _39771_ (_27124_, _08286_, _08285_);
  not _39772_ (_08287_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _39773_ (_08289_, _08262_, _08287_);
  and _39774_ (_08291_, _08262_, word_in[1]);
  nor _39775_ (_08292_, _08291_, _08289_);
  nor _39776_ (_08293_, _08292_, _08260_);
  and _39777_ (_08295_, _08260_, word_in[9]);
  or _39778_ (_08296_, _08295_, _08293_);
  and _39779_ (_08297_, _08296_, _08258_);
  and _39780_ (_08298_, _08257_, _06391_);
  or _39781_ (_08299_, _08298_, _08276_);
  or _39782_ (_08300_, _08299_, _08297_);
  or _39783_ (_08301_, _08282_, _06801_);
  and _39784_ (_26828_[1], _08301_, _08300_);
  and _39785_ (_08302_, _24409_, _23996_);
  and _39786_ (_08303_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or _39787_ (_27121_, _08303_, _08302_);
  not _39788_ (_08304_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _39789_ (_08305_, _08262_, _08304_);
  and _39790_ (_08306_, _08262_, word_in[2]);
  nor _39791_ (_08307_, _08306_, _08305_);
  nor _39792_ (_08308_, _08307_, _08260_);
  and _39793_ (_08309_, _08260_, word_in[10]);
  or _39794_ (_08310_, _08309_, _08308_);
  and _39795_ (_08311_, _08310_, _08258_);
  and _39796_ (_08312_, _08257_, _06572_);
  or _39797_ (_08313_, _08312_, _08276_);
  or _39798_ (_08314_, _08313_, _08311_);
  or _39799_ (_08315_, _08282_, _06407_);
  and _39800_ (_26828_[2], _08315_, _08314_);
  not _39801_ (_08316_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _39802_ (_08317_, _08262_, _08316_);
  and _39803_ (_08318_, _08262_, word_in[3]);
  nor _39804_ (_08319_, _08318_, _08317_);
  nor _39805_ (_08320_, _08319_, _08260_);
  and _39806_ (_08321_, _08260_, word_in[11]);
  or _39807_ (_08322_, _08321_, _08320_);
  and _39808_ (_08323_, _08322_, _08258_);
  and _39809_ (_08324_, _08257_, _06586_);
  or _39810_ (_08325_, _08324_, _08276_);
  or _39811_ (_08326_, _08325_, _08323_);
  or _39812_ (_08327_, _08282_, _06441_);
  and _39813_ (_26828_[3], _08327_, _08326_);
  nand _39814_ (_08328_, _25608_, _23542_);
  and _39815_ (_08329_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _39816_ (_08330_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _39817_ (_08332_, _08330_, _08329_);
  or _39818_ (_08333_, _08332_, _25608_);
  and _39819_ (_08334_, _08333_, _25617_);
  and _39820_ (_08335_, _08334_, _08328_);
  and _39821_ (_08336_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _39822_ (_08337_, _08336_, _08335_);
  and _39823_ (_02719_, _08337_, _22731_);
  not _39824_ (_08338_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _39825_ (_08339_, _08262_, _08338_);
  and _39826_ (_08340_, _08262_, word_in[4]);
  nor _39827_ (_08341_, _08340_, _08339_);
  nor _39828_ (_08342_, _08341_, _08260_);
  and _39829_ (_08343_, _08260_, word_in[12]);
  or _39830_ (_08344_, _08343_, _08342_);
  and _39831_ (_08345_, _08344_, _08258_);
  and _39832_ (_08346_, _08257_, _06591_);
  or _39833_ (_08347_, _08346_, _08276_);
  or _39834_ (_08348_, _08347_, _08345_);
  or _39835_ (_08349_, _08282_, _06446_);
  and _39836_ (_26828_[4], _08349_, _08348_);
  and _39837_ (_08350_, _25414_, _24051_);
  and _39838_ (_08351_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _39839_ (_02721_, _08351_, _08350_);
  not _39840_ (_08352_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _39841_ (_08353_, _08262_, _08352_);
  and _39842_ (_08354_, _08262_, word_in[5]);
  nor _39843_ (_08355_, _08354_, _08353_);
  nor _39844_ (_08356_, _08355_, _08260_);
  and _39845_ (_08357_, _08260_, word_in[13]);
  or _39846_ (_08358_, _08357_, _08356_);
  and _39847_ (_08359_, _08358_, _08258_);
  and _39848_ (_08360_, _08257_, _06606_);
  or _39849_ (_08361_, _08360_, _08276_);
  or _39850_ (_08362_, _08361_, _08359_);
  or _39851_ (_08363_, _08282_, _06463_);
  and _39852_ (_26828_[5], _08363_, _08362_);
  and _39853_ (_08364_, _02368_, _23996_);
  and _39854_ (_08365_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or _39855_ (_02725_, _08365_, _08364_);
  not _39856_ (_08366_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _39857_ (_08367_, _08262_, _08366_);
  and _39858_ (_08368_, _08262_, word_in[6]);
  nor _39859_ (_08370_, _08368_, _08367_);
  nor _39860_ (_08371_, _08370_, _08260_);
  and _39861_ (_08372_, _08260_, word_in[14]);
  or _39862_ (_08373_, _08372_, _08371_);
  and _39863_ (_08374_, _08373_, _08258_);
  and _39864_ (_08375_, _08257_, _06620_);
  or _39865_ (_08376_, _08375_, _08276_);
  or _39866_ (_08377_, _08376_, _08374_);
  or _39867_ (_08379_, _08282_, _06867_);
  and _39868_ (_26828_[6], _08379_, _08377_);
  nor _39869_ (_08380_, _08262_, _05811_);
  and _39870_ (_08382_, _08262_, word_in[7]);
  nor _39871_ (_08383_, _08382_, _08380_);
  nor _39872_ (_08384_, _08383_, _08260_);
  and _39873_ (_08385_, _08260_, word_in[15]);
  or _39874_ (_08386_, _08385_, _08384_);
  and _39875_ (_08387_, _08386_, _08258_);
  and _39876_ (_08388_, _08257_, _06047_);
  or _39877_ (_08389_, _08388_, _08276_);
  or _39878_ (_08390_, _08389_, _08387_);
  or _39879_ (_08391_, _08282_, _06052_);
  and _39880_ (_26828_[7], _08391_, _08390_);
  and _39881_ (_08392_, _02517_, _23548_);
  and _39882_ (_08394_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or _39883_ (_02736_, _08394_, _08392_);
  and _39884_ (_08395_, _05431_, _24051_);
  and _39885_ (_08396_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or _39886_ (_02741_, _08396_, _08395_);
  and _39887_ (_08398_, _04812_, _23887_);
  and _39888_ (_08399_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _39889_ (_02747_, _08399_, _08398_);
  not _39890_ (_08401_, _25608_);
  nor _39891_ (_08402_, _08401_, _24126_);
  and _39892_ (_08403_, _24533_, _24181_);
  and _39893_ (_08404_, _08403_, _25488_);
  and _39894_ (_08405_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _39895_ (_08406_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _39896_ (_08407_, _08406_, _08405_);
  nor _39897_ (_08409_, _08407_, _25608_);
  or _39898_ (_08411_, _08409_, _08404_);
  or _39899_ (_08412_, _08411_, _08402_);
  not _39900_ (_08413_, _08404_);
  or _39901_ (_08414_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _39902_ (_08415_, _08414_, _22731_);
  and _39903_ (_02751_, _08415_, _08412_);
  and _39904_ (_08416_, _02413_, _24219_);
  and _39905_ (_08417_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _39906_ (_27147_, _08417_, _08416_);
  nand _39907_ (_08418_, _25603_, _24082_);
  or _39908_ (_08419_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  not _39909_ (_08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand _39910_ (_08421_, _25609_, _08420_);
  and _39911_ (_08422_, _08421_, _08419_);
  or _39912_ (_08423_, _08422_, _25603_);
  and _39913_ (_08424_, _08423_, _22731_);
  and _39914_ (_02763_, _08424_, _08418_);
  or _39915_ (_08425_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _39916_ (_08426_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _39917_ (_08427_, _08426_, _08425_);
  or _39918_ (_08428_, _08427_, _25603_);
  nand _39919_ (_08429_, _25603_, _24210_);
  and _39920_ (_08430_, _08429_, _22731_);
  and _39921_ (_02766_, _08430_, _08428_);
  and _39922_ (_08431_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  and _39923_ (_08432_, _03011_, _23548_);
  or _39924_ (_02770_, _08432_, _08431_);
  and _39925_ (_08433_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and _39926_ (_08434_, _06203_, _24134_);
  or _39927_ (_02773_, _08434_, _08433_);
  and _39928_ (_08435_, _24159_, _24006_);
  and _39929_ (_08436_, _08435_, _23583_);
  not _39930_ (_08437_, _08435_);
  and _39931_ (_08438_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or _39932_ (_02781_, _08438_, _08436_);
  and _39933_ (_08439_, _25499_, _23577_);
  and _39934_ (_08440_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _39935_ (_08441_, _08440_, _25523_);
  nand _39936_ (_08442_, _25509_, _25507_);
  nor _39937_ (_08443_, _08442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _39938_ (_08444_, _08442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _39939_ (_08445_, _08444_, _25531_);
  or _39940_ (_08446_, _08445_, _08443_);
  or _39941_ (_08447_, _08446_, _08441_);
  not _39942_ (_08448_, _25531_);
  or _39943_ (_08449_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _39944_ (_08450_, _08449_, _25502_);
  and _39945_ (_08451_, _08450_, _08447_);
  and _39946_ (_08452_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _39947_ (_08453_, _08452_, _08451_);
  or _39948_ (_08454_, _08453_, _08439_);
  and _39949_ (_02788_, _08454_, _22731_);
  and _39950_ (_08455_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _39951_ (_08456_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _39952_ (_08457_, _08456_, _25523_);
  and _39953_ (_08458_, _25519_, _25507_);
  nor _39954_ (_08459_, _08458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _39955_ (_08460_, _08459_, _25543_);
  or _39956_ (_08461_, _08460_, _25531_);
  or _39957_ (_08462_, _08461_, _08457_);
  or _39958_ (_08463_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _39959_ (_08464_, _08463_, _25502_);
  and _39960_ (_08465_, _08464_, _08462_);
  or _39961_ (_08466_, _08465_, _08455_);
  and _39962_ (_08467_, _25556_, _25488_);
  and _39963_ (_08468_, _08467_, _24179_);
  and _39964_ (_08469_, _08468_, _02689_);
  or _39965_ (_08470_, _08469_, _08466_);
  and _39966_ (_02791_, _08470_, _22731_);
  and _39967_ (_08471_, _06035_, word_in[0]);
  not _39968_ (_08472_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _39969_ (_08473_, _06035_, _08472_);
  nor _39970_ (_08474_, _08473_, _08471_);
  nor _39971_ (_08475_, _08474_, _06030_);
  and _39972_ (_08476_, _06030_, word_in[8]);
  or _39973_ (_08477_, _08476_, _08475_);
  and _39974_ (_08478_, _08477_, _06027_);
  and _39975_ (_08479_, _06538_, _06026_);
  or _39976_ (_08480_, _08479_, _06046_);
  or _39977_ (_08481_, _08480_, _08478_);
  or _39978_ (_08482_, _06364_, _06051_);
  and _39979_ (_26829_[0], _08482_, _08481_);
  and _39980_ (_08483_, _06035_, word_in[1]);
  not _39981_ (_08484_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _39982_ (_08485_, _06035_, _08484_);
  nor _39983_ (_08486_, _08485_, _08483_);
  nor _39984_ (_08487_, _08486_, _06030_);
  and _39985_ (_08488_, _06030_, word_in[9]);
  or _39986_ (_08489_, _08488_, _08487_);
  and _39987_ (_08491_, _08489_, _06027_);
  and _39988_ (_08492_, _06391_, _06026_);
  or _39989_ (_08493_, _08492_, _06046_);
  or _39990_ (_08494_, _08493_, _08491_);
  or _39991_ (_08495_, _06801_, _06051_);
  and _39992_ (_26829_[1], _08495_, _08494_);
  and _39993_ (_08496_, _06763_, _23996_);
  and _39994_ (_08497_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _39995_ (_02797_, _08497_, _08496_);
  not _39996_ (_08498_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _39997_ (_08499_, _06035_, _08498_);
  and _39998_ (_08500_, _06412_, _06035_);
  or _39999_ (_08501_, _08500_, _08499_);
  or _40000_ (_08502_, _08501_, _06030_);
  not _40001_ (_08503_, _06030_);
  or _40002_ (_08504_, _08503_, word_in[10]);
  and _40003_ (_08505_, _08504_, _08502_);
  or _40004_ (_08506_, _08505_, _06026_);
  or _40005_ (_08507_, _06572_, _06027_);
  and _40006_ (_08508_, _08507_, _08506_);
  or _40007_ (_08509_, _08508_, _06046_);
  or _40008_ (_08510_, _06407_, _06051_);
  and _40009_ (_26829_[2], _08510_, _08509_);
  or _40010_ (_08511_, _08503_, word_in[11]);
  not _40011_ (_08512_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _40012_ (_08513_, _06035_, _08512_);
  and _40013_ (_08514_, _06427_, _06035_);
  or _40014_ (_08515_, _08514_, _08513_);
  or _40015_ (_08516_, _08515_, _06030_);
  and _40016_ (_08517_, _08516_, _06027_);
  and _40017_ (_08518_, _08517_, _08511_);
  and _40018_ (_08519_, _06586_, _06026_);
  or _40019_ (_08520_, _08519_, _06046_);
  or _40020_ (_08521_, _08520_, _08518_);
  or _40021_ (_08522_, _06441_, _06051_);
  and _40022_ (_26829_[3], _08522_, _08521_);
  and _40023_ (_08523_, _24474_, _24006_);
  and _40024_ (_08524_, _08523_, _23548_);
  not _40025_ (_08525_, _08523_);
  and _40026_ (_08526_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or _40027_ (_27081_, _08526_, _08524_);
  and _40028_ (_08527_, _06035_, word_in[4]);
  not _40029_ (_08528_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _40030_ (_08529_, _06035_, _08528_);
  nor _40031_ (_08530_, _08529_, _08527_);
  nor _40032_ (_08531_, _08530_, _06030_);
  and _40033_ (_08532_, _06030_, word_in[12]);
  or _40034_ (_08533_, _08532_, _08531_);
  and _40035_ (_08534_, _08533_, _06027_);
  and _40036_ (_08535_, _06591_, _06026_);
  or _40037_ (_08536_, _08535_, _06046_);
  or _40038_ (_08537_, _08536_, _08534_);
  or _40039_ (_08538_, _06446_, _06051_);
  and _40040_ (_26829_[4], _08538_, _08537_);
  and _40041_ (_08539_, _25479_, _24177_);
  nand _40042_ (_08540_, _08539_, _23504_);
  not _40043_ (_08541_, _25489_);
  or _40044_ (_08542_, _08539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _40045_ (_08543_, _08542_, _08541_);
  and _40046_ (_08544_, _08543_, _08540_);
  nor _40047_ (_08545_, _08541_, _23542_);
  or _40048_ (_08546_, _08545_, _08544_);
  and _40049_ (_02805_, _08546_, _22731_);
  not _40050_ (_08547_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _40051_ (_08548_, _06035_, _08547_);
  and _40052_ (_08549_, _06469_, _06035_);
  or _40053_ (_08550_, _08549_, _08548_);
  or _40054_ (_08551_, _08550_, _06030_);
  or _40055_ (_08552_, _08503_, word_in[13]);
  and _40056_ (_08553_, _08552_, _08551_);
  or _40057_ (_08554_, _08553_, _06026_);
  or _40058_ (_08555_, _06606_, _06027_);
  and _40059_ (_08556_, _08555_, _08554_);
  or _40060_ (_08557_, _08556_, _06046_);
  or _40061_ (_08558_, _06463_, _06051_);
  and _40062_ (_26829_[5], _08558_, _08557_);
  and _40063_ (_08559_, _24223_, _24006_);
  and _40064_ (_08560_, _08559_, _24134_);
  not _40065_ (_08561_, _08559_);
  and _40066_ (_08562_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or _40067_ (_02808_, _08562_, _08560_);
  or _40068_ (_08563_, _08503_, word_in[14]);
  not _40069_ (_08564_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _40070_ (_08565_, _06035_, _08564_);
  and _40071_ (_08566_, _06623_, _06035_);
  or _40072_ (_08567_, _08566_, _08565_);
  or _40073_ (_08568_, _08567_, _06030_);
  and _40074_ (_08569_, _08568_, _06027_);
  and _40075_ (_08570_, _08569_, _08563_);
  and _40076_ (_08571_, _06620_, _06026_);
  or _40077_ (_08573_, _08571_, _06046_);
  or _40078_ (_08574_, _08573_, _08570_);
  or _40079_ (_08575_, _06867_, _06051_);
  and _40080_ (_26829_[6], _08575_, _08574_);
  and _40081_ (_08576_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and _40082_ (_08577_, _06339_, _24134_);
  or _40083_ (_02822_, _08577_, _08576_);
  and _40084_ (_08578_, _24319_, _24006_);
  and _40085_ (_08579_, _08578_, _23996_);
  not _40086_ (_08580_, _08578_);
  and _40087_ (_08581_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or _40088_ (_02828_, _08581_, _08579_);
  and _40089_ (_08582_, _25479_, _24607_);
  nand _40090_ (_08583_, _08582_, _23504_);
  or _40091_ (_08584_, _08582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _40092_ (_08585_, _08584_, _08541_);
  and _40093_ (_08586_, _08585_, _08583_);
  nor _40094_ (_08587_, _08541_, _24043_);
  or _40095_ (_08588_, _08587_, _08586_);
  and _40096_ (_02843_, _08588_, _22731_);
  and _40097_ (_08589_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _40098_ (_08590_, _06339_, _23996_);
  or _40099_ (_02850_, _08590_, _08589_);
  and _40100_ (_08591_, _02039_, _24899_);
  not _40101_ (_08592_, _08591_);
  and _40102_ (_08593_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  and _40103_ (_08594_, _08591_, _23548_);
  or _40104_ (_02853_, _08594_, _08593_);
  and _40105_ (_08595_, _24442_, _23548_);
  and _40106_ (_08596_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or _40107_ (_02864_, _08596_, _08595_);
  and _40108_ (_08598_, _05460_, _23583_);
  and _40109_ (_08599_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _40110_ (_27073_, _08599_, _08598_);
  and _40111_ (_08600_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  and _40112_ (_08601_, _08591_, _23887_);
  or _40113_ (_02878_, _08601_, _08600_);
  and _40114_ (_08603_, _05689_, word_in[0]);
  nand _40115_ (_08604_, _05613_, _07556_);
  or _40116_ (_08605_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _40117_ (_08607_, _08605_, _08604_);
  and _40118_ (_08608_, _08607_, _05649_);
  nand _40119_ (_08609_, _05613_, _08104_);
  or _40120_ (_08610_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _40121_ (_08611_, _08610_, _08609_);
  and _40122_ (_08612_, _08611_, _05629_);
  nand _40123_ (_08613_, _05613_, _07795_);
  or _40124_ (_08614_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _40125_ (_08615_, _08614_, _08613_);
  and _40126_ (_08616_, _08615_, _05632_);
  or _40127_ (_08617_, _08616_, _08612_);
  or _40128_ (_08618_, _08617_, _08608_);
  nand _40129_ (_08619_, _05613_, _08472_);
  or _40130_ (_08620_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _40131_ (_08621_, _08620_, _08619_);
  and _40132_ (_08622_, _08621_, _05639_);
  or _40133_ (_08623_, _08622_, _05724_);
  or _40134_ (_08624_, _08623_, _08618_);
  nand _40135_ (_08625_, _05613_, _06518_);
  or _40136_ (_08626_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _40137_ (_08627_, _08626_, _08625_);
  and _40138_ (_08628_, _08627_, _05649_);
  nand _40139_ (_08630_, _05613_, _06775_);
  or _40140_ (_08631_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _40141_ (_08632_, _08631_, _08630_);
  and _40142_ (_08633_, _08632_, _05632_);
  nand _40143_ (_08635_, _05613_, _07023_);
  or _40144_ (_08636_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _40145_ (_08637_, _08636_, _08635_);
  and _40146_ (_08638_, _08637_, _05629_);
  or _40147_ (_08639_, _08638_, _08633_);
  or _40148_ (_08640_, _08639_, _08628_);
  nand _40149_ (_08641_, _05613_, _07294_);
  or _40150_ (_08642_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _40151_ (_08643_, _08642_, _08641_);
  and _40152_ (_08644_, _08643_, _05639_);
  or _40153_ (_08645_, _08644_, _05617_);
  or _40154_ (_08646_, _08645_, _08640_);
  and _40155_ (_08647_, _08646_, _08624_);
  and _40156_ (_08648_, _08647_, _05688_);
  or _40157_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _08648_, _08603_);
  and _40158_ (_08649_, _05689_, word_in[1]);
  nand _40159_ (_08651_, _05613_, _07573_);
  or _40160_ (_08652_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _40161_ (_08653_, _08652_, _08651_);
  and _40162_ (_08654_, _08653_, _05649_);
  nand _40163_ (_08656_, _05613_, _08117_);
  or _40164_ (_08657_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _40165_ (_08658_, _08657_, _08656_);
  and _40166_ (_08659_, _08658_, _05629_);
  nand _40167_ (_08660_, _05613_, _07816_);
  or _40168_ (_08661_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _40169_ (_08663_, _08661_, _08660_);
  and _40170_ (_08664_, _08663_, _05632_);
  or _40171_ (_08665_, _08664_, _08659_);
  or _40172_ (_08666_, _08665_, _08654_);
  nand _40173_ (_08668_, _05613_, _08484_);
  or _40174_ (_08669_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _40175_ (_08670_, _08669_, _08668_);
  and _40176_ (_08671_, _08670_, _05639_);
  or _40177_ (_08672_, _08671_, _05724_);
  or _40178_ (_08673_, _08672_, _08666_);
  nand _40179_ (_08674_, _05613_, _06545_);
  or _40180_ (_08675_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _40181_ (_08676_, _08675_, _08674_);
  and _40182_ (_08677_, _08676_, _05649_);
  nand _40183_ (_08678_, _05613_, _06790_);
  or _40184_ (_08679_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _40185_ (_08680_, _08679_, _08678_);
  and _40186_ (_08681_, _08680_, _05632_);
  nand _40187_ (_08682_, _05613_, _07046_);
  or _40188_ (_08683_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _40189_ (_08684_, _08683_, _08682_);
  and _40190_ (_08685_, _08684_, _05629_);
  or _40191_ (_08686_, _08685_, _08681_);
  or _40192_ (_08687_, _08686_, _08677_);
  nand _40193_ (_08688_, _05613_, _07310_);
  or _40194_ (_08689_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _40195_ (_08690_, _08689_, _08688_);
  and _40196_ (_08691_, _08690_, _05639_);
  or _40197_ (_08692_, _08691_, _05617_);
  or _40198_ (_08693_, _08692_, _08687_);
  and _40199_ (_08695_, _08693_, _08673_);
  and _40200_ (_08696_, _08695_, _05688_);
  or _40201_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _08696_, _08649_);
  and _40202_ (_08697_, _05689_, word_in[2]);
  nand _40203_ (_08698_, _05613_, _07590_);
  or _40204_ (_08699_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _40205_ (_08700_, _08699_, _08698_);
  and _40206_ (_08702_, _08700_, _05649_);
  nand _40207_ (_08703_, _05613_, _07828_);
  or _40208_ (_08704_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _40209_ (_08705_, _08704_, _08703_);
  and _40210_ (_08706_, _08705_, _05632_);
  nand _40211_ (_08707_, _05613_, _08134_);
  or _40212_ (_08708_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _40213_ (_08709_, _08708_, _08707_);
  and _40214_ (_08710_, _08709_, _05629_);
  or _40215_ (_08712_, _08710_, _08706_);
  or _40216_ (_08713_, _08712_, _08702_);
  nand _40217_ (_08714_, _05613_, _08498_);
  or _40218_ (_08715_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _40219_ (_08716_, _08715_, _08714_);
  and _40220_ (_08717_, _08716_, _05639_);
  or _40221_ (_08718_, _08717_, _05724_);
  or _40222_ (_08719_, _08718_, _08713_);
  nand _40223_ (_08720_, _05613_, _06562_);
  or _40224_ (_08721_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _40225_ (_08722_, _08721_, _08720_);
  and _40226_ (_08723_, _08722_, _05649_);
  nand _40227_ (_08725_, _05613_, _06804_);
  or _40228_ (_08726_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _40229_ (_08727_, _08726_, _08725_);
  and _40230_ (_08729_, _08727_, _05632_);
  nand _40231_ (_08730_, _05613_, _07063_);
  or _40232_ (_08731_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _40233_ (_08732_, _08731_, _08730_);
  and _40234_ (_08733_, _08732_, _05629_);
  or _40235_ (_08734_, _08733_, _08729_);
  or _40236_ (_08735_, _08734_, _08723_);
  nand _40237_ (_08736_, _05613_, _07329_);
  or _40238_ (_08737_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _40239_ (_08739_, _08737_, _08736_);
  and _40240_ (_08740_, _08739_, _05639_);
  or _40241_ (_08741_, _08740_, _05617_);
  or _40242_ (_08742_, _08741_, _08735_);
  and _40243_ (_08743_, _08742_, _08719_);
  and _40244_ (_08744_, _08743_, _05688_);
  or _40245_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _08744_, _08697_);
  and _40246_ (_08745_, _05689_, word_in[3]);
  nand _40247_ (_08747_, _05613_, _07840_);
  or _40248_ (_08748_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _40249_ (_08749_, _08748_, _08747_);
  and _40250_ (_08750_, _08749_, _05632_);
  nand _40251_ (_08751_, _05613_, _08148_);
  or _40252_ (_08752_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _40253_ (_08753_, _08752_, _08751_);
  and _40254_ (_08754_, _08753_, _05629_);
  nand _40255_ (_08755_, _05613_, _07602_);
  or _40256_ (_08756_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _40257_ (_08757_, _08756_, _08755_);
  and _40258_ (_08758_, _08757_, _05649_);
  or _40259_ (_08759_, _08758_, _08754_);
  or _40260_ (_08760_, _08759_, _08750_);
  nand _40261_ (_08761_, _05613_, _08512_);
  or _40262_ (_08762_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _40263_ (_08763_, _08762_, _08761_);
  and _40264_ (_08764_, _08763_, _05639_);
  or _40265_ (_08765_, _08764_, _05724_);
  or _40266_ (_08766_, _08765_, _08760_);
  nand _40267_ (_08768_, _05613_, _06818_);
  or _40268_ (_08769_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _40269_ (_08770_, _08769_, _08768_);
  and _40270_ (_08771_, _08770_, _05632_);
  nand _40271_ (_08772_, _05613_, _06578_);
  or _40272_ (_08773_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _40273_ (_08774_, _08773_, _08772_);
  and _40274_ (_08775_, _08774_, _05649_);
  nand _40275_ (_08776_, _05613_, _07078_);
  or _40276_ (_08777_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _40277_ (_08778_, _08777_, _08776_);
  and _40278_ (_08779_, _08778_, _05629_);
  or _40279_ (_08781_, _08779_, _08775_);
  or _40280_ (_08783_, _08781_, _08771_);
  nand _40281_ (_08784_, _05613_, _07339_);
  or _40282_ (_08785_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _40283_ (_08786_, _08785_, _08784_);
  and _40284_ (_08787_, _08786_, _05639_);
  or _40285_ (_08788_, _08787_, _05617_);
  or _40286_ (_08789_, _08788_, _08783_);
  and _40287_ (_08790_, _08789_, _08766_);
  and _40288_ (_08791_, _08790_, _05688_);
  or _40289_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _08791_, _08745_);
  and _40290_ (_08792_, _05689_, word_in[4]);
  nand _40291_ (_08793_, _05613_, _07854_);
  or _40292_ (_08794_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _40293_ (_08795_, _08794_, _08793_);
  and _40294_ (_08796_, _08795_, _05632_);
  nand _40295_ (_08797_, _05613_, _08162_);
  or _40296_ (_08798_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _40297_ (_08800_, _08798_, _08797_);
  and _40298_ (_08801_, _08800_, _05629_);
  nand _40299_ (_08803_, _05613_, _07616_);
  or _40300_ (_08804_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _40301_ (_08805_, _08804_, _08803_);
  and _40302_ (_08806_, _08805_, _05649_);
  or _40303_ (_08807_, _08806_, _08801_);
  or _40304_ (_08808_, _08807_, _08796_);
  nand _40305_ (_08810_, _05613_, _08528_);
  or _40306_ (_08811_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _40307_ (_08813_, _08811_, _08810_);
  and _40308_ (_08815_, _08813_, _05639_);
  or _40309_ (_08816_, _08815_, _05724_);
  or _40310_ (_08818_, _08816_, _08808_);
  nand _40311_ (_08819_, _05613_, _06832_);
  or _40312_ (_08820_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _40313_ (_08821_, _08820_, _08819_);
  and _40314_ (_08822_, _08821_, _05632_);
  nand _40315_ (_08823_, _05613_, _06594_);
  or _40316_ (_08824_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _40317_ (_08826_, _08824_, _08823_);
  and _40318_ (_08827_, _08826_, _05649_);
  nand _40319_ (_08828_, _05613_, _07096_);
  or _40320_ (_08829_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _40321_ (_08830_, _08829_, _08828_);
  and _40322_ (_08831_, _08830_, _05629_);
  or _40323_ (_08832_, _08831_, _08827_);
  or _40324_ (_08833_, _08832_, _08822_);
  nand _40325_ (_08834_, _05613_, _07357_);
  or _40326_ (_08835_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _40327_ (_08836_, _08835_, _08834_);
  and _40328_ (_08837_, _08836_, _05639_);
  or _40329_ (_08838_, _08837_, _05617_);
  or _40330_ (_08839_, _08838_, _08833_);
  and _40331_ (_08840_, _08839_, _08818_);
  and _40332_ (_08841_, _08840_, _05688_);
  or _40333_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _08841_, _08792_);
  and _40334_ (_08842_, _05689_, word_in[5]);
  nand _40335_ (_08843_, _05613_, _07631_);
  or _40336_ (_08844_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _40337_ (_08846_, _08844_, _08843_);
  and _40338_ (_08848_, _08846_, _05649_);
  nand _40339_ (_08849_, _05613_, _07869_);
  or _40340_ (_08850_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _40341_ (_08852_, _08850_, _08849_);
  and _40342_ (_08853_, _08852_, _05632_);
  nand _40343_ (_08854_, _05613_, _08179_);
  or _40344_ (_08856_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _40345_ (_08857_, _08856_, _08854_);
  and _40346_ (_08858_, _08857_, _05629_);
  or _40347_ (_08859_, _08858_, _08853_);
  or _40348_ (_08860_, _08859_, _08848_);
  nand _40349_ (_08861_, _05613_, _08547_);
  or _40350_ (_08863_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _40351_ (_08864_, _08863_, _08861_);
  and _40352_ (_08866_, _08864_, _05639_);
  or _40353_ (_08867_, _08866_, _05724_);
  or _40354_ (_08868_, _08867_, _08860_);
  nand _40355_ (_08869_, _05613_, _06609_);
  or _40356_ (_08870_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _40357_ (_08871_, _08870_, _08869_);
  and _40358_ (_08872_, _08871_, _05649_);
  nand _40359_ (_08874_, _05613_, _06845_);
  or _40360_ (_08875_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _40361_ (_08876_, _08875_, _08874_);
  and _40362_ (_08877_, _08876_, _05632_);
  nand _40363_ (_08878_, _05613_, _07112_);
  or _40364_ (_08879_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _40365_ (_08880_, _08879_, _08878_);
  and _40366_ (_08881_, _08880_, _05629_);
  or _40367_ (_08882_, _08881_, _08877_);
  or _40368_ (_08883_, _08882_, _08872_);
  nand _40369_ (_08884_, _05613_, _07375_);
  or _40370_ (_08885_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _40371_ (_08886_, _08885_, _08884_);
  and _40372_ (_08888_, _08886_, _05639_);
  or _40373_ (_08889_, _08888_, _05617_);
  or _40374_ (_08890_, _08889_, _08883_);
  and _40375_ (_08891_, _08890_, _08868_);
  and _40376_ (_08893_, _08891_, _05688_);
  or _40377_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _08893_, _08842_);
  and _40378_ (_08894_, _05689_, word_in[6]);
  nand _40379_ (_08895_, _05613_, _07647_);
  or _40380_ (_08897_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _40381_ (_08898_, _08897_, _08895_);
  and _40382_ (_08899_, _08898_, _05649_);
  nand _40383_ (_08900_, _05613_, _08192_);
  or _40384_ (_08901_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _40385_ (_08902_, _08901_, _08900_);
  and _40386_ (_08904_, _08902_, _05629_);
  nand _40387_ (_08906_, _05613_, _07887_);
  or _40388_ (_08908_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _40389_ (_08909_, _08908_, _08906_);
  and _40390_ (_08910_, _08909_, _05632_);
  or _40391_ (_08911_, _08910_, _08904_);
  or _40392_ (_08913_, _08911_, _08899_);
  nand _40393_ (_08914_, _05613_, _08564_);
  or _40394_ (_08915_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _40395_ (_08916_, _08915_, _08914_);
  and _40396_ (_08917_, _08916_, _05639_);
  or _40397_ (_08918_, _08917_, _05724_);
  or _40398_ (_08919_, _08918_, _08913_);
  nand _40399_ (_08920_, _05613_, _06625_);
  or _40400_ (_08921_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _40401_ (_08922_, _08921_, _08920_);
  and _40402_ (_08924_, _08922_, _05649_);
  nand _40403_ (_08926_, _05613_, _06857_);
  or _40404_ (_08927_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _40405_ (_08928_, _08927_, _08926_);
  and _40406_ (_08929_, _08928_, _05632_);
  nand _40407_ (_08930_, _05613_, _07127_);
  or _40408_ (_08931_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _40409_ (_08933_, _08931_, _08930_);
  and _40410_ (_08934_, _08933_, _05629_);
  or _40411_ (_08935_, _08934_, _08929_);
  or _40412_ (_08936_, _08935_, _08924_);
  nand _40413_ (_08937_, _05613_, _07384_);
  or _40414_ (_08938_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _40415_ (_08939_, _08938_, _08937_);
  and _40416_ (_08940_, _08939_, _05639_);
  or _40417_ (_08941_, _08940_, _05617_);
  or _40418_ (_08942_, _08941_, _08936_);
  and _40419_ (_08943_, _08942_, _08919_);
  and _40420_ (_08944_, _08943_, _05688_);
  or _40421_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _08944_, _08894_);
  and _40422_ (_08945_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and _40423_ (_08946_, _08591_, _24051_);
  or _40424_ (_27018_, _08946_, _08945_);
  and _40425_ (_08948_, _05810_, word_in[8]);
  nand _40426_ (_08950_, _05613_, _07674_);
  or _40427_ (_08951_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _40428_ (_08952_, _08951_, _08950_);
  and _40429_ (_08953_, _08952_, _05787_);
  nand _40430_ (_08954_, _05613_, _07428_);
  or _40431_ (_08955_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _40432_ (_08956_, _08955_, _08954_);
  and _40433_ (_08957_, _08956_, _05785_);
  or _40434_ (_08958_, _08957_, _08953_);
  and _40435_ (_08959_, _08958_, _05763_);
  nand _40436_ (_08960_, _05613_, _06655_);
  or _40437_ (_08961_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _40438_ (_08962_, _08961_, _08960_);
  and _40439_ (_08963_, _08962_, _05787_);
  nand _40440_ (_08964_, _05613_, _06375_);
  or _40441_ (_08965_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _40442_ (_08966_, _08965_, _08964_);
  and _40443_ (_08967_, _08966_, _05785_);
  or _40444_ (_08968_, _08967_, _08963_);
  and _40445_ (_08969_, _08968_, _05767_);
  nand _40446_ (_08970_, _05613_, _07170_);
  or _40447_ (_08972_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _40448_ (_08973_, _08972_, _08970_);
  and _40449_ (_08974_, _08973_, _05787_);
  nand _40450_ (_08975_, _05613_, _06892_);
  or _40451_ (_08976_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _40452_ (_08977_, _08976_, _08975_);
  and _40453_ (_08978_, _08977_, _05785_);
  or _40454_ (_08979_, _08978_, _08974_);
  and _40455_ (_08980_, _08979_, _05797_);
  or _40456_ (_08981_, _08980_, _08969_);
  nand _40457_ (_08982_, _05613_, _08264_);
  or _40458_ (_08983_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _40459_ (_08984_, _08983_, _08982_);
  and _40460_ (_08985_, _08984_, _05787_);
  nand _40461_ (_08987_, _05613_, _07950_);
  or _40462_ (_08988_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _40463_ (_08990_, _08988_, _08987_);
  and _40464_ (_08991_, _08990_, _05785_);
  or _40465_ (_08993_, _08991_, _08985_);
  and _40466_ (_08994_, _08993_, _05800_);
  or _40467_ (_08996_, _08994_, _08981_);
  nor _40468_ (_08997_, _08996_, _08959_);
  nor _40469_ (_08998_, _08997_, _05810_);
  or _40470_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _08998_, _08948_);
  and _40471_ (_09000_, _05810_, word_in[9]);
  nand _40472_ (_09001_, _05613_, _07688_);
  or _40473_ (_09003_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _40474_ (_09005_, _09003_, _09001_);
  and _40475_ (_09006_, _09005_, _05787_);
  nand _40476_ (_09007_, _05613_, _07443_);
  or _40477_ (_09010_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _40478_ (_09011_, _09010_, _09007_);
  and _40479_ (_09012_, _09011_, _05785_);
  or _40480_ (_09013_, _09012_, _09006_);
  and _40481_ (_09015_, _09013_, _05763_);
  nand _40482_ (_09016_, _05613_, _06674_);
  or _40483_ (_09018_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _40484_ (_09019_, _09018_, _09016_);
  and _40485_ (_09020_, _09019_, _05787_);
  nand _40486_ (_09021_, _05613_, _06393_);
  or _40487_ (_09022_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _40488_ (_09023_, _09022_, _09021_);
  and _40489_ (_09024_, _09023_, _05785_);
  or _40490_ (_09025_, _09024_, _09020_);
  and _40491_ (_09026_, _09025_, _05767_);
  nand _40492_ (_09027_, _05613_, _07183_);
  or _40493_ (_09028_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _40494_ (_09029_, _09028_, _09027_);
  and _40495_ (_09030_, _09029_, _05787_);
  nand _40496_ (_09031_, _05613_, _06908_);
  or _40497_ (_09033_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _40498_ (_09035_, _09033_, _09031_);
  and _40499_ (_09036_, _09035_, _05785_);
  or _40500_ (_09037_, _09036_, _09030_);
  and _40501_ (_09039_, _09037_, _05797_);
  or _40502_ (_09040_, _09039_, _09026_);
  nand _40503_ (_09041_, _05613_, _08287_);
  or _40504_ (_09043_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _40505_ (_09044_, _09043_, _09041_);
  and _40506_ (_09045_, _09044_, _05787_);
  nand _40507_ (_09046_, _05613_, _07974_);
  or _40508_ (_09047_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _40509_ (_09049_, _09047_, _09046_);
  and _40510_ (_09050_, _09049_, _05785_);
  or _40511_ (_09051_, _09050_, _09045_);
  and _40512_ (_09052_, _09051_, _05800_);
  or _40513_ (_09053_, _09052_, _09040_);
  nor _40514_ (_09054_, _09053_, _09015_);
  nor _40515_ (_09055_, _09054_, _05810_);
  or _40516_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _09055_, _09000_);
  and _40517_ (_09058_, _05810_, word_in[10]);
  nand _40518_ (_09060_, _05613_, _07700_);
  or _40519_ (_09062_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _40520_ (_09064_, _09062_, _09060_);
  and _40521_ (_09065_, _09064_, _05787_);
  nand _40522_ (_09066_, _05613_, _07458_);
  or _40523_ (_09067_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _40524_ (_09068_, _09067_, _09066_);
  and _40525_ (_09070_, _09068_, _05785_);
  or _40526_ (_09071_, _09070_, _09065_);
  and _40527_ (_09072_, _09071_, _05763_);
  nand _40528_ (_09073_, _05613_, _06686_);
  or _40529_ (_09074_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _40530_ (_09075_, _09074_, _09073_);
  and _40531_ (_09076_, _09075_, _05787_);
  nand _40532_ (_09077_, _05613_, _06410_);
  or _40533_ (_09078_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _40534_ (_09080_, _09078_, _09077_);
  and _40535_ (_09081_, _09080_, _05785_);
  or _40536_ (_09082_, _09081_, _09076_);
  and _40537_ (_09083_, _09082_, _05767_);
  nand _40538_ (_09084_, _05613_, _07203_);
  or _40539_ (_09085_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _40540_ (_09086_, _09085_, _09084_);
  and _40541_ (_09087_, _09086_, _05787_);
  nand _40542_ (_09088_, _05613_, _06920_);
  or _40543_ (_09089_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _40544_ (_09090_, _09089_, _09088_);
  and _40545_ (_09091_, _09090_, _05785_);
  or _40546_ (_09092_, _09091_, _09087_);
  and _40547_ (_09094_, _09092_, _05797_);
  or _40548_ (_09095_, _09094_, _09083_);
  nand _40549_ (_09097_, _05613_, _08304_);
  or _40550_ (_09098_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _40551_ (_09099_, _09098_, _09097_);
  and _40552_ (_09100_, _09099_, _05787_);
  nand _40553_ (_09101_, _05613_, _07992_);
  or _40554_ (_09102_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _40555_ (_09104_, _09102_, _09101_);
  and _40556_ (_09105_, _09104_, _05785_);
  or _40557_ (_09106_, _09105_, _09100_);
  and _40558_ (_09107_, _09106_, _05800_);
  or _40559_ (_09109_, _09107_, _09095_);
  nor _40560_ (_09110_, _09109_, _09072_);
  nor _40561_ (_09111_, _09110_, _05810_);
  or _40562_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _09111_, _09058_);
  and _40563_ (_09114_, _05810_, word_in[11]);
  nand _40564_ (_09115_, _05613_, _07714_);
  or _40565_ (_09116_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _40566_ (_09117_, _09116_, _09115_);
  and _40567_ (_09120_, _09117_, _05787_);
  nand _40568_ (_09121_, _05613_, _07473_);
  or _40569_ (_09123_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _40570_ (_09124_, _09123_, _09121_);
  and _40571_ (_09125_, _09124_, _05785_);
  or _40572_ (_09126_, _09125_, _09120_);
  and _40573_ (_09127_, _09126_, _05763_);
  nand _40574_ (_09128_, _05613_, _06699_);
  or _40575_ (_09129_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _40576_ (_09131_, _09129_, _09128_);
  and _40577_ (_09132_, _09131_, _05787_);
  nand _40578_ (_09134_, _05613_, _06425_);
  or _40579_ (_09135_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _40580_ (_09137_, _09135_, _09134_);
  and _40581_ (_09138_, _09137_, _05785_);
  or _40582_ (_09140_, _09138_, _09132_);
  and _40583_ (_09142_, _09140_, _05767_);
  nand _40584_ (_09143_, _05613_, _07218_);
  or _40585_ (_09144_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _40586_ (_09146_, _09144_, _09143_);
  and _40587_ (_09149_, _09146_, _05787_);
  nand _40588_ (_09150_, _05613_, _06934_);
  or _40589_ (_09151_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _40590_ (_09153_, _09151_, _09150_);
  and _40591_ (_09154_, _09153_, _05785_);
  or _40592_ (_09155_, _09154_, _09149_);
  and _40593_ (_09156_, _09155_, _05797_);
  or _40594_ (_09158_, _09156_, _09142_);
  nand _40595_ (_09160_, _05613_, _08316_);
  or _40596_ (_09161_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _40597_ (_09162_, _09161_, _09160_);
  and _40598_ (_09163_, _09162_, _05787_);
  nand _40599_ (_09164_, _05613_, _08008_);
  or _40600_ (_09165_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _40601_ (_09166_, _09165_, _09164_);
  and _40602_ (_09167_, _09166_, _05785_);
  or _40603_ (_09168_, _09167_, _09163_);
  and _40604_ (_09169_, _09168_, _05800_);
  or _40605_ (_09170_, _09169_, _09158_);
  nor _40606_ (_09171_, _09170_, _09127_);
  nor _40607_ (_09172_, _09171_, _05810_);
  or _40608_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _09172_, _09114_);
  and _40609_ (_09173_, _05810_, word_in[12]);
  nand _40610_ (_09174_, _05613_, _07726_);
  or _40611_ (_09175_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _40612_ (_09176_, _09175_, _09174_);
  and _40613_ (_09178_, _09176_, _05787_);
  nand _40614_ (_09179_, _05613_, _07486_);
  or _40615_ (_09181_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _40616_ (_09182_, _09181_, _09179_);
  and _40617_ (_09184_, _09182_, _05785_);
  or _40618_ (_09185_, _09184_, _09178_);
  and _40619_ (_09186_, _09185_, _05763_);
  nand _40620_ (_09187_, _05613_, _08338_);
  or _40621_ (_09189_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _40622_ (_09190_, _09189_, _09187_);
  and _40623_ (_09192_, _09190_, _05787_);
  nand _40624_ (_09193_, _05613_, _08026_);
  or _40625_ (_09194_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _40626_ (_09195_, _09194_, _09193_);
  and _40627_ (_09197_, _09195_, _05785_);
  or _40628_ (_09199_, _09197_, _09192_);
  and _40629_ (_09200_, _09199_, _05800_);
  nand _40630_ (_09202_, _05613_, _07234_);
  or _40631_ (_09203_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _40632_ (_09204_, _09203_, _09202_);
  and _40633_ (_09205_, _09204_, _05787_);
  nand _40634_ (_09206_, _05613_, _06946_);
  or _40635_ (_09208_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _40636_ (_09210_, _09208_, _09206_);
  and _40637_ (_09212_, _09210_, _05785_);
  or _40638_ (_09213_, _09212_, _09205_);
  and _40639_ (_09215_, _09213_, _05797_);
  nand _40640_ (_09217_, _05613_, _06711_);
  or _40641_ (_09219_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _40642_ (_09221_, _09219_, _09217_);
  and _40643_ (_09222_, _09221_, _05787_);
  nand _40644_ (_09223_, _05613_, _06448_);
  or _40645_ (_09225_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _40646_ (_09227_, _09225_, _09223_);
  and _40647_ (_09229_, _09227_, _05785_);
  or _40648_ (_09231_, _09229_, _09222_);
  and _40649_ (_09233_, _09231_, _05767_);
  or _40650_ (_09234_, _09233_, _09215_);
  or _40651_ (_09235_, _09234_, _09200_);
  nor _40652_ (_09236_, _09235_, _09186_);
  nor _40653_ (_09237_, _09236_, _05810_);
  or _40654_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _09237_, _09173_);
  and _40655_ (_09238_, _05810_, word_in[13]);
  nand _40656_ (_09239_, _05613_, _07738_);
  or _40657_ (_09240_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _40658_ (_09241_, _09240_, _09239_);
  and _40659_ (_09242_, _09241_, _05787_);
  nand _40660_ (_09243_, _05613_, _07498_);
  or _40661_ (_09244_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _40662_ (_09245_, _09244_, _09243_);
  and _40663_ (_09246_, _09245_, _05785_);
  or _40664_ (_09247_, _09246_, _09242_);
  and _40665_ (_09248_, _09247_, _05763_);
  nand _40666_ (_09249_, _05613_, _08352_);
  or _40667_ (_09250_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _40668_ (_09251_, _09250_, _09249_);
  and _40669_ (_09252_, _09251_, _05787_);
  nand _40670_ (_09253_, _05613_, _08040_);
  or _40671_ (_09254_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _40672_ (_09255_, _09254_, _09253_);
  and _40673_ (_09257_, _09255_, _05785_);
  or _40674_ (_09258_, _09257_, _09252_);
  and _40675_ (_09259_, _09258_, _05800_);
  nand _40676_ (_09260_, _05613_, _07247_);
  or _40677_ (_09261_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _40678_ (_09262_, _09261_, _09260_);
  and _40679_ (_09263_, _09262_, _05787_);
  nand _40680_ (_09264_, _05613_, _06961_);
  or _40681_ (_09265_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _40682_ (_09266_, _09265_, _09264_);
  and _40683_ (_09267_, _09266_, _05785_);
  or _40684_ (_09269_, _09267_, _09263_);
  and _40685_ (_09271_, _09269_, _05797_);
  nand _40686_ (_09272_, _05613_, _06726_);
  or _40687_ (_09273_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _40688_ (_09274_, _09273_, _09272_);
  and _40689_ (_09275_, _09274_, _05787_);
  nand _40690_ (_09277_, _05613_, _06466_);
  or _40691_ (_09278_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _40692_ (_09279_, _09278_, _09277_);
  and _40693_ (_09280_, _09279_, _05785_);
  or _40694_ (_09281_, _09280_, _09275_);
  and _40695_ (_09282_, _09281_, _05767_);
  or _40696_ (_09283_, _09282_, _09271_);
  or _40697_ (_09284_, _09283_, _09259_);
  nor _40698_ (_09285_, _09284_, _09248_);
  nor _40699_ (_09286_, _09285_, _05810_);
  or _40700_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _09286_, _09238_);
  and _40701_ (_09288_, _05810_, word_in[14]);
  nand _40702_ (_09289_, _05613_, _07752_);
  or _40703_ (_09290_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _40704_ (_09291_, _09290_, _09289_);
  and _40705_ (_09292_, _09291_, _05787_);
  nand _40706_ (_09293_, _05613_, _07517_);
  or _40707_ (_09294_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _40708_ (_09295_, _09294_, _09293_);
  and _40709_ (_09296_, _09295_, _05785_);
  or _40710_ (_09297_, _09296_, _09292_);
  and _40711_ (_09298_, _09297_, _05763_);
  nand _40712_ (_09299_, _05613_, _08366_);
  or _40713_ (_09300_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _40714_ (_09301_, _09300_, _09299_);
  and _40715_ (_09302_, _09301_, _05787_);
  nand _40716_ (_09303_, _05613_, _08052_);
  or _40717_ (_09304_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _40718_ (_09305_, _09304_, _09303_);
  and _40719_ (_09306_, _09305_, _05785_);
  or _40720_ (_09307_, _09306_, _09302_);
  and _40721_ (_09308_, _09307_, _05800_);
  nand _40722_ (_09309_, _05613_, _07260_);
  or _40723_ (_09310_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _40724_ (_09311_, _09310_, _09309_);
  and _40725_ (_09312_, _09311_, _05787_);
  nand _40726_ (_09313_, _05613_, _06976_);
  or _40727_ (_09314_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _40728_ (_09315_, _09314_, _09313_);
  and _40729_ (_09316_, _09315_, _05785_);
  or _40730_ (_09318_, _09316_, _09312_);
  and _40731_ (_09319_, _09318_, _05797_);
  nand _40732_ (_09320_, _05613_, _06738_);
  or _40733_ (_09321_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _40734_ (_09322_, _09321_, _09320_);
  and _40735_ (_09323_, _09322_, _05787_);
  nand _40736_ (_09324_, _05613_, _06481_);
  or _40737_ (_09325_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _40738_ (_09326_, _09325_, _09324_);
  and _40739_ (_09327_, _09326_, _05785_);
  or _40740_ (_09329_, _09327_, _09323_);
  and _40741_ (_09330_, _09329_, _05767_);
  or _40742_ (_09332_, _09330_, _09319_);
  or _40743_ (_09333_, _09332_, _09308_);
  nor _40744_ (_09334_, _09333_, _09298_);
  nor _40745_ (_09335_, _09334_, _05810_);
  or _40746_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _09335_, _09288_);
  and _40747_ (_09336_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and _40748_ (_09337_, _08591_, _23996_);
  or _40749_ (_02933_, _09337_, _09336_);
  and _40750_ (_09338_, _05918_, word_in[16]);
  and _40751_ (_09339_, _08627_, _05639_);
  and _40752_ (_09340_, _08643_, _05629_);
  or _40753_ (_09341_, _09340_, _09339_);
  and _40754_ (_09342_, _08637_, _05632_);
  and _40755_ (_09343_, _08632_, _05649_);
  or _40756_ (_09344_, _09343_, _09342_);
  or _40757_ (_09345_, _09344_, _09341_);
  or _40758_ (_09346_, _09345_, _05921_);
  and _40759_ (_09348_, _08611_, _05632_);
  and _40760_ (_09349_, _08607_, _05639_);
  or _40761_ (_09350_, _09349_, _09348_);
  and _40762_ (_09351_, _08621_, _05629_);
  and _40763_ (_09352_, _08615_, _05649_);
  or _40764_ (_09353_, _09352_, _09351_);
  nor _40765_ (_09354_, _09353_, _09350_);
  nand _40766_ (_09355_, _09354_, _05921_);
  nand _40767_ (_09356_, _09355_, _09346_);
  nor _40768_ (_09358_, _09356_, _05918_);
  or _40769_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _09358_, _09338_);
  and _40770_ (_09359_, _05918_, word_in[17]);
  and _40771_ (_09360_, _08684_, _05632_);
  and _40772_ (_09361_, _08676_, _05639_);
  or _40773_ (_09362_, _09361_, _09360_);
  and _40774_ (_09363_, _08690_, _05629_);
  and _40775_ (_09364_, _08680_, _05649_);
  or _40776_ (_09365_, _09364_, _09363_);
  or _40777_ (_09366_, _09365_, _09362_);
  or _40778_ (_09368_, _09366_, _05921_);
  and _40779_ (_09369_, _08653_, _05639_);
  and _40780_ (_09370_, _08670_, _05629_);
  or _40781_ (_09371_, _09370_, _09369_);
  and _40782_ (_09372_, _08658_, _05632_);
  and _40783_ (_09373_, _08663_, _05649_);
  or _40784_ (_09374_, _09373_, _09372_);
  nor _40785_ (_09375_, _09374_, _09371_);
  nand _40786_ (_09376_, _09375_, _05921_);
  nand _40787_ (_09377_, _09376_, _09368_);
  nor _40788_ (_09378_, _09377_, _05918_);
  or _40789_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _09378_, _09359_);
  and _40790_ (_09379_, _05918_, word_in[18]);
  and _40791_ (_09380_, _08722_, _05639_);
  and _40792_ (_09381_, _08739_, _05629_);
  or _40793_ (_09382_, _09381_, _09380_);
  and _40794_ (_09383_, _08732_, _05632_);
  and _40795_ (_09384_, _08727_, _05649_);
  or _40796_ (_09385_, _09384_, _09383_);
  or _40797_ (_09386_, _09385_, _09382_);
  or _40798_ (_09387_, _09386_, _05921_);
  and _40799_ (_09388_, _08700_, _05639_);
  and _40800_ (_09389_, _08716_, _05629_);
  or _40801_ (_09390_, _09389_, _09388_);
  and _40802_ (_09392_, _08709_, _05632_);
  and _40803_ (_09393_, _08705_, _05649_);
  or _40804_ (_09394_, _09393_, _09392_);
  nor _40805_ (_09395_, _09394_, _09390_);
  nand _40806_ (_09396_, _09395_, _05921_);
  nand _40807_ (_09397_, _09396_, _09387_);
  nor _40808_ (_09398_, _09397_, _05918_);
  or _40809_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _09398_, _09379_);
  and _40810_ (_09399_, _05918_, word_in[19]);
  and _40811_ (_09400_, _08778_, _05632_);
  and _40812_ (_09401_, _08774_, _05639_);
  or _40813_ (_09403_, _09401_, _09400_);
  and _40814_ (_09404_, _08786_, _05629_);
  and _40815_ (_09405_, _08770_, _05649_);
  or _40816_ (_09406_, _09405_, _09404_);
  or _40817_ (_09407_, _09406_, _09403_);
  or _40818_ (_09408_, _09407_, _05921_);
  and _40819_ (_09409_, _08757_, _05639_);
  and _40820_ (_09410_, _08763_, _05629_);
  or _40821_ (_09411_, _09410_, _09409_);
  and _40822_ (_09413_, _08753_, _05632_);
  and _40823_ (_09414_, _08749_, _05649_);
  or _40824_ (_09415_, _09414_, _09413_);
  nor _40825_ (_09417_, _09415_, _09411_);
  nand _40826_ (_09418_, _09417_, _05921_);
  nand _40827_ (_09419_, _09418_, _09408_);
  nor _40828_ (_09420_, _09419_, _05918_);
  or _40829_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _09420_, _09399_);
  and _40830_ (_09421_, _05918_, word_in[20]);
  and _40831_ (_09422_, _08826_, _05639_);
  and _40832_ (_09423_, _08836_, _05629_);
  or _40833_ (_09424_, _09423_, _09422_);
  and _40834_ (_09425_, _08830_, _05632_);
  and _40835_ (_09426_, _08821_, _05649_);
  or _40836_ (_09428_, _09426_, _09425_);
  or _40837_ (_09429_, _09428_, _09424_);
  or _40838_ (_09430_, _09429_, _05921_);
  and _40839_ (_09431_, _08805_, _05639_);
  and _40840_ (_09432_, _08813_, _05629_);
  or _40841_ (_09433_, _09432_, _09431_);
  and _40842_ (_09434_, _08800_, _05632_);
  and _40843_ (_09435_, _08795_, _05649_);
  or _40844_ (_09436_, _09435_, _09434_);
  nor _40845_ (_09437_, _09436_, _09433_);
  nand _40846_ (_09438_, _09437_, _05921_);
  nand _40847_ (_09439_, _09438_, _09430_);
  nor _40848_ (_09440_, _09439_, _05918_);
  or _40849_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _09440_, _09421_);
  and _40850_ (_09441_, _05918_, word_in[21]);
  and _40851_ (_09442_, _08871_, _05639_);
  and _40852_ (_09443_, _08886_, _05629_);
  or _40853_ (_09444_, _09443_, _09442_);
  and _40854_ (_09445_, _08880_, _05632_);
  and _40855_ (_09446_, _08876_, _05649_);
  or _40856_ (_09447_, _09446_, _09445_);
  or _40857_ (_09449_, _09447_, _09444_);
  or _40858_ (_09450_, _09449_, _05921_);
  and _40859_ (_09451_, _08857_, _05632_);
  and _40860_ (_09452_, _08846_, _05639_);
  or _40861_ (_09453_, _09452_, _09451_);
  and _40862_ (_09454_, _08864_, _05629_);
  and _40863_ (_09455_, _08852_, _05649_);
  or _40864_ (_09456_, _09455_, _09454_);
  nor _40865_ (_09457_, _09456_, _09453_);
  nand _40866_ (_09458_, _09457_, _05921_);
  nand _40867_ (_09459_, _09458_, _09450_);
  nor _40868_ (_09460_, _09459_, _05918_);
  or _40869_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _09460_, _09441_);
  and _40870_ (_09461_, _05918_, word_in[22]);
  and _40871_ (_09463_, _08933_, _05632_);
  and _40872_ (_09464_, _08922_, _05639_);
  or _40873_ (_09465_, _09464_, _09463_);
  and _40874_ (_09466_, _08939_, _05629_);
  and _40875_ (_09467_, _08928_, _05649_);
  or _40876_ (_09468_, _09467_, _09466_);
  or _40877_ (_09469_, _09468_, _09465_);
  or _40878_ (_09470_, _09469_, _05921_);
  and _40879_ (_09471_, _08902_, _05632_);
  and _40880_ (_09472_, _08898_, _05639_);
  or _40881_ (_09473_, _09472_, _09471_);
  and _40882_ (_09474_, _08916_, _05629_);
  and _40883_ (_09475_, _08909_, _05649_);
  or _40884_ (_09476_, _09475_, _09474_);
  nor _40885_ (_09477_, _09476_, _09473_);
  nand _40886_ (_09478_, _09477_, _05921_);
  nand _40887_ (_09480_, _09478_, _09470_);
  nor _40888_ (_09481_, _09480_, _05918_);
  or _40889_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _09481_, _09461_);
  and _40890_ (_09482_, _05991_, word_in[24]);
  and _40891_ (_09483_, _08956_, _05787_);
  and _40892_ (_09484_, _08952_, _05785_);
  or _40893_ (_09485_, _09484_, _09483_);
  and _40894_ (_09486_, _09485_, _05957_);
  and _40895_ (_09487_, _08966_, _05787_);
  and _40896_ (_09488_, _08962_, _05785_);
  or _40897_ (_09489_, _09488_, _09487_);
  and _40898_ (_09490_, _09489_, _05996_);
  and _40899_ (_09491_, _08977_, _05787_);
  and _40900_ (_09492_, _08973_, _05785_);
  or _40901_ (_09493_, _09492_, _09491_);
  and _40902_ (_09494_, _09493_, _06003_);
  and _40903_ (_09495_, _08990_, _05787_);
  and _40904_ (_09496_, _08984_, _05785_);
  or _40905_ (_09497_, _09496_, _09495_);
  and _40906_ (_09498_, _09497_, _06008_);
  or _40907_ (_09500_, _09498_, _09494_);
  or _40908_ (_09501_, _09500_, _09490_);
  nor _40909_ (_09502_, _09501_, _09486_);
  nor _40910_ (_09503_, _09502_, _05991_);
  or _40911_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _09503_, _09482_);
  and _40912_ (_09504_, _05991_, word_in[25]);
  and _40913_ (_09505_, _09011_, _05787_);
  and _40914_ (_09506_, _09005_, _05785_);
  or _40915_ (_09507_, _09506_, _09505_);
  and _40916_ (_09508_, _09507_, _05957_);
  and _40917_ (_09509_, _09023_, _05787_);
  and _40918_ (_09510_, _09019_, _05785_);
  or _40919_ (_09511_, _09510_, _09509_);
  and _40920_ (_09512_, _09511_, _05996_);
  and _40921_ (_09514_, _09035_, _05787_);
  and _40922_ (_09515_, _09029_, _05785_);
  or _40923_ (_09516_, _09515_, _09514_);
  and _40924_ (_09517_, _09516_, _06003_);
  and _40925_ (_09518_, _09049_, _05787_);
  and _40926_ (_09519_, _09044_, _05785_);
  or _40927_ (_09520_, _09519_, _09518_);
  and _40928_ (_09521_, _09520_, _06008_);
  or _40929_ (_09522_, _09521_, _09517_);
  or _40930_ (_09523_, _09522_, _09512_);
  nor _40931_ (_09524_, _09523_, _09508_);
  nor _40932_ (_09525_, _09524_, _05991_);
  or _40933_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _09525_, _09504_);
  and _40934_ (_09526_, _05991_, word_in[26]);
  and _40935_ (_09527_, _09068_, _05787_);
  and _40936_ (_09528_, _09064_, _05785_);
  or _40937_ (_09529_, _09528_, _09527_);
  and _40938_ (_09530_, _09529_, _05957_);
  and _40939_ (_09531_, _09080_, _05787_);
  and _40940_ (_09532_, _09075_, _05785_);
  or _40941_ (_09533_, _09532_, _09531_);
  and _40942_ (_09534_, _09533_, _05996_);
  and _40943_ (_09535_, _09090_, _05787_);
  and _40944_ (_09536_, _09086_, _05785_);
  or _40945_ (_09537_, _09536_, _09535_);
  and _40946_ (_09538_, _09537_, _06003_);
  and _40947_ (_09540_, _09104_, _05787_);
  and _40948_ (_09541_, _09099_, _05785_);
  or _40949_ (_09542_, _09541_, _09540_);
  and _40950_ (_09543_, _09542_, _06008_);
  or _40951_ (_09545_, _09543_, _09538_);
  or _40952_ (_09546_, _09545_, _09534_);
  nor _40953_ (_09547_, _09546_, _09530_);
  nor _40954_ (_09548_, _09547_, _05991_);
  or _40955_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _09548_, _09526_);
  and _40956_ (_09549_, _05991_, word_in[27]);
  and _40957_ (_09550_, _09137_, _05787_);
  and _40958_ (_09551_, _09131_, _05785_);
  or _40959_ (_09552_, _09551_, _09550_);
  and _40960_ (_09553_, _09552_, _05996_);
  and _40961_ (_09554_, _09124_, _05787_);
  and _40962_ (_09555_, _09117_, _05785_);
  or _40963_ (_09556_, _09555_, _09554_);
  and _40964_ (_09557_, _09556_, _05957_);
  and _40965_ (_09558_, _09153_, _05787_);
  and _40966_ (_09559_, _09146_, _05785_);
  or _40967_ (_09561_, _09559_, _09558_);
  and _40968_ (_09562_, _09561_, _06003_);
  and _40969_ (_09563_, _09166_, _05787_);
  and _40970_ (_09564_, _09162_, _05785_);
  or _40971_ (_09565_, _09564_, _09563_);
  and _40972_ (_09566_, _09565_, _06008_);
  or _40973_ (_09567_, _09566_, _09562_);
  or _40974_ (_09568_, _09567_, _09557_);
  nor _40975_ (_09569_, _09568_, _09553_);
  nor _40976_ (_09570_, _09569_, _05991_);
  or _40977_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _09570_, _09549_);
  and _40978_ (_09571_, _05991_, word_in[28]);
  and _40979_ (_09572_, _09227_, _05787_);
  and _40980_ (_09573_, _09221_, _05785_);
  or _40981_ (_09574_, _09573_, _09572_);
  and _40982_ (_09575_, _09574_, _05996_);
  and _40983_ (_09576_, _09182_, _05787_);
  and _40984_ (_09577_, _09176_, _05785_);
  or _40985_ (_09578_, _09577_, _09576_);
  and _40986_ (_09579_, _09578_, _05957_);
  and _40987_ (_09581_, _09210_, _05787_);
  and _40988_ (_09582_, _09204_, _05785_);
  or _40989_ (_09583_, _09582_, _09581_);
  and _40990_ (_09584_, _09583_, _06003_);
  and _40991_ (_09585_, _09195_, _05787_);
  and _40992_ (_09586_, _09190_, _05785_);
  or _40993_ (_09587_, _09586_, _09585_);
  and _40994_ (_09588_, _09587_, _06008_);
  or _40995_ (_09589_, _09588_, _09584_);
  or _40996_ (_09590_, _09589_, _09579_);
  nor _40997_ (_09591_, _09590_, _09575_);
  nor _40998_ (_09592_, _09591_, _05991_);
  or _40999_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _09592_, _09571_);
  and _41000_ (_09593_, _05991_, word_in[29]);
  and _41001_ (_09594_, _09245_, _05787_);
  and _41002_ (_09595_, _09241_, _05785_);
  or _41003_ (_09596_, _09595_, _09594_);
  and _41004_ (_09597_, _09596_, _05957_);
  and _41005_ (_09598_, _09279_, _05787_);
  and _41006_ (_09599_, _09274_, _05785_);
  or _41007_ (_09601_, _09599_, _09598_);
  and _41008_ (_09602_, _09601_, _05996_);
  and _41009_ (_09603_, _09266_, _05787_);
  and _41010_ (_09604_, _09262_, _05785_);
  or _41011_ (_09605_, _09604_, _09603_);
  and _41012_ (_09606_, _09605_, _06003_);
  and _41013_ (_09607_, _09255_, _05787_);
  and _41014_ (_09608_, _09251_, _05785_);
  or _41015_ (_09609_, _09608_, _09607_);
  and _41016_ (_09610_, _09609_, _06008_);
  or _41017_ (_09611_, _09610_, _09606_);
  or _41018_ (_09612_, _09611_, _09602_);
  nor _41019_ (_09614_, _09612_, _09597_);
  nor _41020_ (_09615_, _09614_, _05991_);
  or _41021_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _09615_, _09593_);
  and _41022_ (_09616_, _05991_, word_in[30]);
  and _41023_ (_09617_, _09295_, _05787_);
  and _41024_ (_09618_, _09291_, _05785_);
  or _41025_ (_09619_, _09618_, _09617_);
  and _41026_ (_09620_, _09619_, _05957_);
  and _41027_ (_09622_, _09326_, _05787_);
  and _41028_ (_09623_, _09322_, _05785_);
  or _41029_ (_09624_, _09623_, _09622_);
  and _41030_ (_09625_, _09624_, _05996_);
  and _41031_ (_09626_, _09315_, _05787_);
  and _41032_ (_09627_, _09311_, _05785_);
  or _41033_ (_09628_, _09627_, _09626_);
  and _41034_ (_09629_, _09628_, _06003_);
  and _41035_ (_09631_, _09305_, _05787_);
  and _41036_ (_09632_, _09301_, _05785_);
  or _41037_ (_09633_, _09632_, _09631_);
  and _41038_ (_09634_, _09633_, _06008_);
  or _41039_ (_09635_, _09634_, _09629_);
  or _41040_ (_09636_, _09635_, _09625_);
  nor _41041_ (_09637_, _09636_, _09620_);
  nor _41042_ (_09638_, _09637_, _05991_);
  or _41043_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _09638_, _09616_);
  and _41044_ (_09639_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _41045_ (_09640_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _41046_ (_09641_, _22740_, _09640_);
  or _41047_ (_09642_, _09641_, _09639_);
  and _41048_ (_26862_[1], _09642_, _22731_);
  and _41049_ (_09643_, _24350_, _24134_);
  and _41050_ (_09644_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _41051_ (_27062_, _09644_, _09643_);
  and _41052_ (_09645_, _02039_, _23941_);
  not _41053_ (_09646_, _09645_);
  and _41054_ (_09647_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and _41055_ (_09648_, _09645_, _24219_);
  or _41056_ (_03000_, _09648_, _09647_);
  and _41057_ (_09651_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and _41058_ (_09652_, _09645_, _23887_);
  or _41059_ (_03012_, _09652_, _09651_);
  and _41060_ (_09653_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and _41061_ (_09654_, _09645_, _24089_);
  or _41062_ (_03027_, _09654_, _09653_);
  and _41063_ (_09655_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and _41064_ (_09656_, _09645_, _24134_);
  or _41065_ (_03047_, _09656_, _09655_);
  and _41066_ (_09657_, _24415_, _24089_);
  and _41067_ (_09658_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or _41068_ (_03051_, _09658_, _09657_);
  and _41069_ (_09659_, _24485_, _24134_);
  and _41070_ (_09660_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or _41071_ (_03053_, _09660_, _09659_);
  and _41072_ (_09661_, _25206_, _23583_);
  and _41073_ (_09663_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _41074_ (_03056_, _09663_, _09661_);
  and _41075_ (_09665_, _25442_, _23996_);
  and _41076_ (_09667_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _41077_ (_27035_, _09667_, _09665_);
  and _41078_ (_09668_, _25648_, _24134_);
  and _41079_ (_09669_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or _41080_ (_27032_, _09669_, _09668_);
  and _41081_ (_09670_, _24365_, _24236_);
  and _41082_ (_09671_, _09670_, _23996_);
  not _41083_ (_09672_, _09670_);
  and _41084_ (_09673_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or _41085_ (_03063_, _09673_, _09671_);
  and _41086_ (_09674_, _25648_, _23887_);
  and _41087_ (_09675_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or _41088_ (_03064_, _09675_, _09674_);
  and _41089_ (_09676_, _02039_, _24349_);
  not _41090_ (_09677_, _09676_);
  and _41091_ (_09678_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _41092_ (_09679_, _09676_, _23548_);
  or _41093_ (_03069_, _09679_, _09678_);
  and _41094_ (_09680_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _41095_ (_09681_, _09676_, _24089_);
  or _41096_ (_03076_, _09681_, _09680_);
  and _41097_ (_09682_, _24442_, _24134_);
  and _41098_ (_09683_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or _41099_ (_03079_, _09683_, _09682_);
  and _41100_ (_09684_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and _41101_ (_09685_, _02338_, _24219_);
  or _41102_ (_03092_, _09685_, _09684_);
  and _41103_ (_09687_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and _41104_ (_09689_, _02836_, _24051_);
  or _41105_ (_03095_, _09689_, _09687_);
  and _41106_ (_09690_, _02990_, _23583_);
  and _41107_ (_09692_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or _41108_ (_03099_, _09692_, _09690_);
  and _41109_ (_09693_, _02990_, _24219_);
  and _41110_ (_09694_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or _41111_ (_27053_, _09694_, _09693_);
  and _41112_ (_09695_, _03186_, _24089_);
  and _41113_ (_09696_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or _41114_ (_03103_, _09696_, _09695_);
  and _41115_ (_09697_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _41116_ (_09698_, _09676_, _24051_);
  or _41117_ (_27022_, _09698_, _09697_);
  and _41118_ (_09699_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _41119_ (_09700_, _09676_, _23996_);
  or _41120_ (_03112_, _09700_, _09699_);
  and _41121_ (_09701_, _02065_, _23583_);
  and _41122_ (_09702_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or _41123_ (_03116_, _09702_, _09701_);
  and _41124_ (_09703_, _24051_, _24008_);
  and _41125_ (_09704_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _41126_ (_03117_, _09704_, _09703_);
  and _41127_ (_09705_, _02039_, _24236_);
  not _41128_ (_09706_, _09705_);
  and _41129_ (_09707_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _41130_ (_09708_, _09705_, _24219_);
  or _41131_ (_03123_, _09708_, _09707_);
  and _41132_ (_09709_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _41133_ (_09710_, _09705_, _23583_);
  or _41134_ (_03125_, _09710_, _09709_);
  and _41135_ (_09711_, _24889_, _24051_);
  and _41136_ (_09712_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _41137_ (_03130_, _09712_, _09711_);
  and _41138_ (_09713_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _41139_ (_09714_, _09705_, _24089_);
  or _41140_ (_03154_, _09714_, _09713_);
  and _41141_ (_09715_, _04920_, _23583_);
  and _41142_ (_09716_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _41143_ (_03156_, _09716_, _09715_);
  and _41144_ (_09717_, _24159_, _23945_);
  and _41145_ (_09718_, _09717_, _24089_);
  not _41146_ (_09719_, _09717_);
  and _41147_ (_09720_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _41148_ (_03160_, _09720_, _09718_);
  and _41149_ (_09722_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and _41150_ (_09723_, _09705_, _24134_);
  or _41151_ (_03163_, _09723_, _09722_);
  and _41152_ (_09724_, _24237_, _23583_);
  and _41153_ (_09725_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _41154_ (_27063_, _09725_, _09724_);
  and _41155_ (_09726_, _24330_, _24134_);
  and _41156_ (_09727_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _41157_ (_03177_, _09727_, _09726_);
  and _41158_ (_09728_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and _41159_ (_09729_, _09705_, _23996_);
  or _41160_ (_03179_, _09729_, _09728_);
  and _41161_ (_09730_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _41162_ (_09731_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _41163_ (_09732_, _22740_, _09731_);
  or _41164_ (_09733_, _09732_, _09730_);
  and _41165_ (_26862_[0], _09733_, _22731_);
  and _41166_ (_09734_, _02478_, _24219_);
  and _41167_ (_09736_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _41168_ (_03196_, _09736_, _09734_);
  and _41169_ (_09737_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and _41170_ (_09738_, _04853_, _24134_);
  or _41171_ (_03206_, _09738_, _09737_);
  and _41172_ (_09739_, _25442_, _23887_);
  and _41173_ (_09740_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _41174_ (_03216_, _09740_, _09739_);
  and _41175_ (_09742_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  and _41176_ (_09744_, _04853_, _24051_);
  or _41177_ (_03223_, _09744_, _09742_);
  and _41178_ (_09746_, _02990_, _23996_);
  and _41179_ (_09747_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or _41180_ (_03240_, _09747_, _09746_);
  and _41181_ (_09749_, _23890_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _41182_ (_09750_, _23845_, _26578_);
  and _41183_ (_09751_, _23909_, _23800_);
  or _41184_ (_09752_, _03899_, _09751_);
  or _41185_ (_09753_, _09752_, _09750_);
  not _41186_ (_09754_, _26736_);
  or _41187_ (_09756_, _24253_, _23913_);
  or _41188_ (_09757_, _09756_, _09754_);
  or _41189_ (_09758_, _09757_, _09753_);
  or _41190_ (_09759_, _23916_, _23839_);
  or _41191_ (_09760_, _26739_, _23901_);
  or _41192_ (_09761_, _09760_, _09759_);
  and _41193_ (_09762_, _23841_, _23708_);
  and _41194_ (_09763_, _24247_, _23896_);
  or _41195_ (_09764_, _09763_, _24248_);
  or _41196_ (_09765_, _09764_, _09762_);
  or _41197_ (_09767_, _09765_, _23906_);
  or _41198_ (_09769_, _09767_, _09761_);
  or _41199_ (_09771_, _09769_, _23934_);
  or _41200_ (_09772_, _09771_, _09758_);
  and _41201_ (_09773_, _09772_, _23855_);
  or _41202_ (_26850_[0], _09773_, _09749_);
  and _41203_ (_09774_, _24496_, _24319_);
  and _41204_ (_09775_, _09774_, _24051_);
  not _41205_ (_09777_, _09774_);
  and _41206_ (_09778_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or _41207_ (_03262_, _09778_, _09775_);
  and _41208_ (_09779_, _23944_, _22977_);
  and _41209_ (_09780_, _09779_, _24159_);
  and _41210_ (_09781_, _09780_, _23996_);
  not _41211_ (_09782_, _09780_);
  and _41212_ (_09783_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _41213_ (_27006_, _09783_, _09781_);
  and _41214_ (_09784_, _07013_, _24219_);
  and _41215_ (_09785_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or _41216_ (_03268_, _09785_, _09784_);
  and _41217_ (_09787_, _09780_, _24134_);
  and _41218_ (_09789_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _41219_ (_27005_, _09789_, _09787_);
  not _41220_ (_09790_, _05520_);
  not _41221_ (_09791_, _05535_);
  and _41222_ (_09792_, _05548_, _05547_);
  and _41223_ (_09793_, _05513_, _05511_);
  and _41224_ (_09794_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and _41225_ (_09795_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _41226_ (_09796_, _09795_, _09794_);
  and _41227_ (_09797_, _09796_, _09792_);
  and _41228_ (_09798_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and _41229_ (_09799_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _41230_ (_09801_, _09799_, _09798_);
  and _41231_ (_09802_, _09801_, _05549_);
  or _41232_ (_09803_, _09802_, _09797_);
  or _41233_ (_09804_, _09803_, _09791_);
  not _41234_ (_09805_, _05542_);
  and _41235_ (_09806_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and _41236_ (_09808_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _41237_ (_09811_, _09808_, _09806_);
  and _41238_ (_09812_, _09811_, _09792_);
  and _41239_ (_09813_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and _41240_ (_09814_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _41241_ (_09815_, _09814_, _09813_);
  and _41242_ (_09816_, _09815_, _05549_);
  or _41243_ (_09817_, _09816_, _09812_);
  or _41244_ (_09818_, _09817_, _05535_);
  and _41245_ (_09819_, _09818_, _09805_);
  and _41246_ (_09820_, _09819_, _09804_);
  or _41247_ (_09821_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _41248_ (_09822_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and _41249_ (_09823_, _09822_, _09821_);
  and _41250_ (_09824_, _09823_, _09792_);
  or _41251_ (_09825_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _41252_ (_09827_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and _41253_ (_09828_, _09827_, _09825_);
  and _41254_ (_09829_, _09828_, _05549_);
  or _41255_ (_09830_, _09829_, _09824_);
  or _41256_ (_09831_, _09830_, _09791_);
  or _41257_ (_09832_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _41258_ (_09833_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and _41259_ (_09834_, _09833_, _09832_);
  and _41260_ (_09836_, _09834_, _09792_);
  or _41261_ (_09838_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _41262_ (_09839_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and _41263_ (_09840_, _09839_, _09838_);
  and _41264_ (_09841_, _09840_, _05549_);
  or _41265_ (_09842_, _09841_, _09836_);
  or _41266_ (_09843_, _09842_, _05535_);
  and _41267_ (_09845_, _09843_, _05542_);
  and _41268_ (_09847_, _09845_, _09831_);
  or _41269_ (_09848_, _09847_, _09820_);
  and _41270_ (_09849_, _09848_, _05518_);
  not _41271_ (_09850_, _05518_);
  and _41272_ (_09851_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and _41273_ (_09852_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _41274_ (_09853_, _09852_, _09851_);
  and _41275_ (_09855_, _09853_, _09792_);
  and _41276_ (_09856_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and _41277_ (_09857_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _41278_ (_09858_, _09857_, _09856_);
  and _41279_ (_09859_, _09858_, _05549_);
  or _41280_ (_09860_, _09859_, _09855_);
  or _41281_ (_09861_, _09860_, _09791_);
  and _41282_ (_09862_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and _41283_ (_09863_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _41284_ (_09865_, _09863_, _09862_);
  and _41285_ (_09866_, _09865_, _09792_);
  and _41286_ (_09867_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and _41287_ (_09869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _41288_ (_09870_, _09869_, _09867_);
  and _41289_ (_09871_, _09870_, _05549_);
  or _41290_ (_09872_, _09871_, _09866_);
  or _41291_ (_09873_, _09872_, _05535_);
  and _41292_ (_09874_, _09873_, _09805_);
  and _41293_ (_09876_, _09874_, _09861_);
  or _41294_ (_09877_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _41295_ (_09878_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and _41296_ (_09879_, _09878_, _05549_);
  and _41297_ (_09880_, _09879_, _09877_);
  or _41298_ (_09882_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _41299_ (_09883_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and _41300_ (_09885_, _09883_, _09792_);
  and _41301_ (_09887_, _09885_, _09882_);
  or _41302_ (_09888_, _09887_, _09880_);
  or _41303_ (_09889_, _09888_, _09791_);
  or _41304_ (_09890_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _41305_ (_09892_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and _41306_ (_09893_, _09892_, _05549_);
  and _41307_ (_09895_, _09893_, _09890_);
  or _41308_ (_09897_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _41309_ (_09898_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and _41310_ (_09899_, _09898_, _09792_);
  and _41311_ (_09900_, _09899_, _09897_);
  or _41312_ (_09901_, _09900_, _09895_);
  or _41313_ (_09902_, _09901_, _05535_);
  and _41314_ (_09903_, _09902_, _05542_);
  and _41315_ (_09904_, _09903_, _09889_);
  or _41316_ (_09905_, _09904_, _09876_);
  and _41317_ (_09906_, _09905_, _09850_);
  or _41318_ (_09907_, _09906_, _09849_);
  and _41319_ (_09909_, _09907_, _09790_);
  and _41320_ (_09910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _41321_ (_09912_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _41322_ (_09913_, _09912_, _09910_);
  and _41323_ (_09915_, _09913_, _09792_);
  and _41324_ (_09917_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _41325_ (_09919_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _41326_ (_09921_, _09919_, _09917_);
  and _41327_ (_09923_, _09921_, _05549_);
  or _41328_ (_09924_, _09923_, _09915_);
  and _41329_ (_09925_, _09924_, _05535_);
  and _41330_ (_09926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _41331_ (_09927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _41332_ (_09928_, _09927_, _09926_);
  and _41333_ (_09930_, _09928_, _09792_);
  and _41334_ (_09931_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _41335_ (_09932_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _41336_ (_09933_, _09932_, _09931_);
  and _41337_ (_09934_, _09933_, _05549_);
  or _41338_ (_09935_, _09934_, _09930_);
  and _41339_ (_09936_, _09935_, _09791_);
  or _41340_ (_09937_, _09936_, _09925_);
  and _41341_ (_09938_, _09937_, _09805_);
  or _41342_ (_09940_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _41343_ (_09941_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _41344_ (_09942_, _09941_, _05549_);
  and _41345_ (_09943_, _09942_, _09940_);
  or _41346_ (_09944_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _41347_ (_09945_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _41348_ (_09946_, _09945_, _09792_);
  and _41349_ (_09947_, _09946_, _09944_);
  or _41350_ (_09948_, _09947_, _09943_);
  and _41351_ (_09949_, _09948_, _05535_);
  or _41352_ (_09951_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _41353_ (_09952_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _41354_ (_09954_, _09952_, _05549_);
  and _41355_ (_09956_, _09954_, _09951_);
  or _41356_ (_09957_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _41357_ (_09958_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and _41358_ (_09960_, _09958_, _09792_);
  and _41359_ (_09962_, _09960_, _09957_);
  or _41360_ (_09963_, _09962_, _09956_);
  and _41361_ (_09964_, _09963_, _09791_);
  or _41362_ (_09965_, _09964_, _09949_);
  and _41363_ (_09967_, _09965_, _05542_);
  or _41364_ (_09968_, _09967_, _09938_);
  and _41365_ (_09969_, _09968_, _09850_);
  and _41366_ (_09971_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and _41367_ (_09973_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _41368_ (_09975_, _09973_, _09971_);
  and _41369_ (_09976_, _09975_, _09792_);
  and _41370_ (_09978_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and _41371_ (_09979_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _41372_ (_09981_, _09979_, _09978_);
  and _41373_ (_09982_, _09981_, _05549_);
  or _41374_ (_09983_, _09982_, _09976_);
  and _41375_ (_09984_, _09983_, _05535_);
  and _41376_ (_09985_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and _41377_ (_09987_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _41378_ (_09988_, _09987_, _09985_);
  and _41379_ (_09989_, _09988_, _09792_);
  and _41380_ (_09990_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and _41381_ (_09991_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _41382_ (_09992_, _09991_, _09990_);
  and _41383_ (_09993_, _09992_, _05549_);
  or _41384_ (_09994_, _09993_, _09989_);
  and _41385_ (_09995_, _09994_, _09791_);
  or _41386_ (_09997_, _09995_, _09984_);
  and _41387_ (_09998_, _09997_, _09805_);
  or _41388_ (_09999_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _41389_ (_10000_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and _41390_ (_10002_, _10000_, _09999_);
  and _41391_ (_10004_, _10002_, _09792_);
  or _41392_ (_10005_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _41393_ (_10007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and _41394_ (_10009_, _10007_, _10005_);
  and _41395_ (_10010_, _10009_, _05549_);
  or _41396_ (_10011_, _10010_, _10004_);
  and _41397_ (_10013_, _10011_, _05535_);
  or _41398_ (_10014_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _41399_ (_10015_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and _41400_ (_10016_, _10015_, _10014_);
  and _41401_ (_10017_, _10016_, _09792_);
  or _41402_ (_10019_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _41403_ (_10020_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and _41404_ (_10021_, _10020_, _10019_);
  and _41405_ (_10022_, _10021_, _05549_);
  or _41406_ (_10023_, _10022_, _10017_);
  and _41407_ (_10024_, _10023_, _09791_);
  or _41408_ (_10025_, _10024_, _10013_);
  and _41409_ (_10026_, _10025_, _05542_);
  or _41410_ (_10027_, _10026_, _09998_);
  and _41411_ (_10028_, _10027_, _05518_);
  or _41412_ (_10029_, _10028_, _09969_);
  and _41413_ (_10030_, _10029_, _05520_);
  or _41414_ (_10031_, _10030_, _09909_);
  or _41415_ (_10032_, _10031_, _05526_);
  not _41416_ (_10033_, _05526_);
  and _41417_ (_10034_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and _41418_ (_10035_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _41419_ (_10036_, _10035_, _10034_);
  and _41420_ (_10037_, _10036_, _09792_);
  and _41421_ (_10038_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and _41422_ (_10039_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _41423_ (_10041_, _10039_, _10038_);
  and _41424_ (_10042_, _10041_, _05549_);
  or _41425_ (_10044_, _10042_, _10037_);
  or _41426_ (_10046_, _10044_, _09791_);
  and _41427_ (_10047_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and _41428_ (_10049_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _41429_ (_10051_, _10049_, _10047_);
  and _41430_ (_10052_, _10051_, _09792_);
  and _41431_ (_10053_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and _41432_ (_10054_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _41433_ (_10056_, _10054_, _10053_);
  and _41434_ (_10057_, _10056_, _05549_);
  or _41435_ (_10058_, _10057_, _10052_);
  or _41436_ (_10060_, _10058_, _05535_);
  and _41437_ (_10062_, _10060_, _09805_);
  and _41438_ (_10063_, _10062_, _10046_);
  or _41439_ (_10064_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _41440_ (_10065_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and _41441_ (_10066_, _10065_, _05549_);
  and _41442_ (_10067_, _10066_, _10064_);
  or _41443_ (_10068_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _41444_ (_10069_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and _41445_ (_10071_, _10069_, _09792_);
  and _41446_ (_10072_, _10071_, _10068_);
  or _41447_ (_10073_, _10072_, _10067_);
  or _41448_ (_10074_, _10073_, _09791_);
  or _41449_ (_10075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _41450_ (_10076_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and _41451_ (_10077_, _10076_, _05549_);
  and _41452_ (_10078_, _10077_, _10075_);
  or _41453_ (_10079_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _41454_ (_10080_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and _41455_ (_10081_, _10080_, _09792_);
  and _41456_ (_10082_, _10081_, _10079_);
  or _41457_ (_10083_, _10082_, _10078_);
  or _41458_ (_10084_, _10083_, _05535_);
  and _41459_ (_10085_, _10084_, _05542_);
  and _41460_ (_10086_, _10085_, _10074_);
  or _41461_ (_10087_, _10086_, _10063_);
  and _41462_ (_10088_, _10087_, _09850_);
  and _41463_ (_10089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and _41464_ (_10091_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _41465_ (_10092_, _10091_, _10089_);
  and _41466_ (_10094_, _10092_, _09792_);
  and _41467_ (_10095_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and _41468_ (_10096_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _41469_ (_10098_, _10096_, _10095_);
  and _41470_ (_10099_, _10098_, _05549_);
  or _41471_ (_10100_, _10099_, _10094_);
  or _41472_ (_10101_, _10100_, _09791_);
  and _41473_ (_10103_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and _41474_ (_10104_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _41475_ (_10105_, _10104_, _10103_);
  and _41476_ (_10106_, _10105_, _09792_);
  and _41477_ (_10108_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _41478_ (_10109_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _41479_ (_10110_, _10109_, _10108_);
  and _41480_ (_10112_, _10110_, _05549_);
  or _41481_ (_10114_, _10112_, _10106_);
  or _41482_ (_10116_, _10114_, _05535_);
  and _41483_ (_10117_, _10116_, _09805_);
  and _41484_ (_10119_, _10117_, _10101_);
  or _41485_ (_10121_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _41486_ (_10122_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and _41487_ (_10123_, _10122_, _10121_);
  and _41488_ (_10124_, _10123_, _09792_);
  or _41489_ (_10125_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _41490_ (_10127_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and _41491_ (_10128_, _10127_, _10125_);
  and _41492_ (_10129_, _10128_, _05549_);
  or _41493_ (_10131_, _10129_, _10124_);
  or _41494_ (_10133_, _10131_, _09791_);
  or _41495_ (_10134_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _41496_ (_10135_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and _41497_ (_10137_, _10135_, _10134_);
  and _41498_ (_10138_, _10137_, _09792_);
  or _41499_ (_10139_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _41500_ (_10141_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _41501_ (_10142_, _10141_, _10139_);
  and _41502_ (_10143_, _10142_, _05549_);
  or _41503_ (_10145_, _10143_, _10138_);
  or _41504_ (_10146_, _10145_, _05535_);
  and _41505_ (_10148_, _10146_, _05542_);
  and _41506_ (_10149_, _10148_, _10133_);
  or _41507_ (_10150_, _10149_, _10119_);
  and _41508_ (_10152_, _10150_, _05518_);
  or _41509_ (_10153_, _10152_, _10088_);
  and _41510_ (_10155_, _10153_, _09790_);
  or _41511_ (_10156_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _41512_ (_10157_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and _41513_ (_10158_, _10157_, _10156_);
  and _41514_ (_10159_, _10158_, _09792_);
  or _41515_ (_10160_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _41516_ (_10162_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and _41517_ (_10163_, _10162_, _10160_);
  and _41518_ (_10164_, _10163_, _05549_);
  or _41519_ (_10165_, _10164_, _10159_);
  and _41520_ (_10167_, _10165_, _09791_);
  or _41521_ (_10168_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _41522_ (_10169_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and _41523_ (_10171_, _10169_, _10168_);
  and _41524_ (_10172_, _10171_, _09792_);
  or _41525_ (_10174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _41526_ (_10176_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and _41527_ (_10178_, _10176_, _10174_);
  and _41528_ (_10180_, _10178_, _05549_);
  or _41529_ (_10182_, _10180_, _10172_);
  and _41530_ (_10183_, _10182_, _05535_);
  or _41531_ (_10184_, _10183_, _10167_);
  and _41532_ (_10185_, _10184_, _05542_);
  and _41533_ (_10187_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and _41534_ (_10188_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _41535_ (_10189_, _10188_, _10187_);
  and _41536_ (_10191_, _10189_, _09792_);
  and _41537_ (_10192_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and _41538_ (_10193_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _41539_ (_10195_, _10193_, _10192_);
  and _41540_ (_10197_, _10195_, _05549_);
  or _41541_ (_10199_, _10197_, _10191_);
  and _41542_ (_10200_, _10199_, _09791_);
  and _41543_ (_10202_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and _41544_ (_10203_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _41545_ (_10204_, _10203_, _10202_);
  and _41546_ (_10205_, _10204_, _09792_);
  and _41547_ (_10206_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and _41548_ (_10207_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _41549_ (_10208_, _10207_, _10206_);
  and _41550_ (_10209_, _10208_, _05549_);
  or _41551_ (_10210_, _10209_, _10205_);
  and _41552_ (_10211_, _10210_, _05535_);
  or _41553_ (_10212_, _10211_, _10200_);
  and _41554_ (_10213_, _10212_, _09805_);
  or _41555_ (_10215_, _10213_, _10185_);
  and _41556_ (_10216_, _10215_, _05518_);
  or _41557_ (_10217_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _41558_ (_10218_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and _41559_ (_10219_, _10218_, _05549_);
  and _41560_ (_10221_, _10219_, _10217_);
  or _41561_ (_10222_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _41562_ (_10223_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _41563_ (_10224_, _10223_, _09792_);
  and _41564_ (_10225_, _10224_, _10222_);
  or _41565_ (_10226_, _10225_, _10221_);
  and _41566_ (_10227_, _10226_, _09791_);
  or _41567_ (_10228_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _41568_ (_10229_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and _41569_ (_10230_, _10229_, _05549_);
  and _41570_ (_10231_, _10230_, _10228_);
  or _41571_ (_10232_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _41572_ (_10233_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and _41573_ (_10234_, _10233_, _09792_);
  and _41574_ (_10235_, _10234_, _10232_);
  or _41575_ (_10236_, _10235_, _10231_);
  and _41576_ (_10237_, _10236_, _05535_);
  or _41577_ (_10238_, _10237_, _10227_);
  and _41578_ (_10239_, _10238_, _05542_);
  and _41579_ (_10240_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and _41580_ (_10241_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _41581_ (_10243_, _10241_, _10240_);
  and _41582_ (_10245_, _10243_, _09792_);
  and _41583_ (_10246_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and _41584_ (_10247_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _41585_ (_10248_, _10247_, _10246_);
  and _41586_ (_10249_, _10248_, _05549_);
  or _41587_ (_10251_, _10249_, _10245_);
  and _41588_ (_10252_, _10251_, _09791_);
  and _41589_ (_10253_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and _41590_ (_10254_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _41591_ (_10255_, _10254_, _10253_);
  and _41592_ (_10256_, _10255_, _09792_);
  and _41593_ (_10257_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and _41594_ (_10258_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _41595_ (_10259_, _10258_, _10257_);
  and _41596_ (_10261_, _10259_, _05549_);
  or _41597_ (_10262_, _10261_, _10256_);
  and _41598_ (_10263_, _10262_, _05535_);
  or _41599_ (_10264_, _10263_, _10252_);
  and _41600_ (_10265_, _10264_, _09805_);
  or _41601_ (_10267_, _10265_, _10239_);
  and _41602_ (_10268_, _10267_, _09850_);
  or _41603_ (_10269_, _10268_, _10216_);
  and _41604_ (_10270_, _10269_, _05520_);
  or _41605_ (_10271_, _10270_, _10155_);
  or _41606_ (_10272_, _10271_, _10033_);
  and _41607_ (_10273_, _10272_, _10032_);
  or _41608_ (_10274_, _10273_, _00143_);
  and _41609_ (_10275_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _41610_ (_10276_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or _41611_ (_10277_, _10276_, _10275_);
  and _41612_ (_10278_, _10277_, _05549_);
  and _41613_ (_10279_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and _41614_ (_10280_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _41615_ (_10281_, _10280_, _10279_);
  and _41616_ (_10282_, _10281_, _09792_);
  or _41617_ (_10283_, _10282_, _10278_);
  or _41618_ (_10284_, _10283_, _09791_);
  and _41619_ (_10285_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _41620_ (_10286_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or _41621_ (_10287_, _10286_, _10285_);
  and _41622_ (_10288_, _10287_, _05549_);
  and _41623_ (_10289_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _41624_ (_10290_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _41625_ (_10291_, _10290_, _10289_);
  and _41626_ (_10292_, _10291_, _09792_);
  or _41627_ (_10294_, _10292_, _10288_);
  or _41628_ (_10295_, _10294_, _05535_);
  and _41629_ (_10296_, _10295_, _09805_);
  and _41630_ (_10297_, _10296_, _10284_);
  or _41631_ (_10298_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or _41632_ (_10299_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and _41633_ (_10300_, _10299_, _09792_);
  and _41634_ (_10301_, _10300_, _10298_);
  or _41635_ (_10302_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _41636_ (_10303_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _41637_ (_10305_, _10303_, _05549_);
  and _41638_ (_10306_, _10305_, _10302_);
  or _41639_ (_10307_, _10306_, _10301_);
  or _41640_ (_10308_, _10307_, _09791_);
  or _41641_ (_10309_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or _41642_ (_10310_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and _41643_ (_10311_, _10310_, _09792_);
  and _41644_ (_10312_, _10311_, _10309_);
  or _41645_ (_10313_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _41646_ (_10314_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _41647_ (_10315_, _10314_, _05549_);
  and _41648_ (_10316_, _10315_, _10313_);
  or _41649_ (_10317_, _10316_, _10312_);
  or _41650_ (_10318_, _10317_, _05535_);
  and _41651_ (_10319_, _10318_, _05542_);
  and _41652_ (_10320_, _10319_, _10308_);
  or _41653_ (_10321_, _10320_, _10297_);
  and _41654_ (_10322_, _10321_, _09850_);
  and _41655_ (_10323_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and _41656_ (_10325_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _41657_ (_10326_, _10325_, _09792_);
  or _41658_ (_10327_, _10326_, _10323_);
  and _41659_ (_10328_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and _41660_ (_10329_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _41661_ (_10330_, _10329_, _05549_);
  or _41662_ (_10331_, _10330_, _10328_);
  and _41663_ (_10332_, _10331_, _10327_);
  or _41664_ (_10333_, _10332_, _09791_);
  and _41665_ (_10334_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and _41666_ (_10335_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _41667_ (_10336_, _10335_, _09792_);
  or _41668_ (_10338_, _10336_, _10334_);
  and _41669_ (_10339_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and _41670_ (_10340_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _41671_ (_10341_, _10340_, _05549_);
  or _41672_ (_10342_, _10341_, _10339_);
  and _41673_ (_10343_, _10342_, _10338_);
  or _41674_ (_10344_, _10343_, _05535_);
  and _41675_ (_10345_, _10344_, _09805_);
  and _41676_ (_10346_, _10345_, _10333_);
  or _41677_ (_10348_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _41678_ (_10349_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and _41679_ (_10350_, _10349_, _10348_);
  or _41680_ (_10351_, _10350_, _05549_);
  or _41681_ (_10352_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _41682_ (_10353_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and _41683_ (_10354_, _10353_, _10352_);
  or _41684_ (_10355_, _10354_, _09792_);
  and _41685_ (_10356_, _10355_, _10351_);
  or _41686_ (_10357_, _10356_, _09791_);
  or _41687_ (_10359_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _41688_ (_10360_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and _41689_ (_10361_, _10360_, _10359_);
  or _41690_ (_10362_, _10361_, _05549_);
  or _41691_ (_10363_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _41692_ (_10364_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and _41693_ (_10365_, _10364_, _10363_);
  or _41694_ (_10367_, _10365_, _09792_);
  and _41695_ (_10368_, _10367_, _10362_);
  or _41696_ (_10369_, _10368_, _05535_);
  and _41697_ (_10370_, _10369_, _05542_);
  and _41698_ (_10371_, _10370_, _10357_);
  or _41699_ (_10372_, _10371_, _10346_);
  and _41700_ (_10373_, _10372_, _05518_);
  or _41701_ (_10374_, _10373_, _10322_);
  and _41702_ (_10376_, _10374_, _09790_);
  and _41703_ (_10377_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and _41704_ (_10378_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or _41705_ (_10380_, _10378_, _10377_);
  and _41706_ (_10381_, _10380_, _09792_);
  and _41707_ (_10383_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  and _41708_ (_10384_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or _41709_ (_10385_, _10384_, _10383_);
  and _41710_ (_10386_, _10385_, _05549_);
  or _41711_ (_10387_, _10386_, _10381_);
  and _41712_ (_10388_, _10387_, _05535_);
  and _41713_ (_10389_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  and _41714_ (_10390_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or _41715_ (_10391_, _10390_, _10389_);
  and _41716_ (_10392_, _10391_, _09792_);
  and _41717_ (_10393_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and _41718_ (_10394_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or _41719_ (_10395_, _10394_, _10393_);
  and _41720_ (_10396_, _10395_, _05549_);
  or _41721_ (_10397_, _10396_, _10392_);
  and _41722_ (_10398_, _10397_, _09791_);
  or _41723_ (_10399_, _10398_, _10388_);
  and _41724_ (_10400_, _10399_, _09805_);
  or _41725_ (_10401_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or _41726_ (_10402_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  and _41727_ (_10403_, _10402_, _10401_);
  and _41728_ (_10404_, _10403_, _09792_);
  or _41729_ (_10405_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or _41730_ (_10406_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and _41731_ (_10407_, _10406_, _10405_);
  and _41732_ (_10408_, _10407_, _05549_);
  or _41733_ (_10409_, _10408_, _10404_);
  and _41734_ (_10410_, _10409_, _05535_);
  or _41735_ (_10411_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or _41736_ (_10412_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  and _41737_ (_10413_, _10412_, _10411_);
  and _41738_ (_10414_, _10413_, _09792_);
  or _41739_ (_10415_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or _41740_ (_10416_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  and _41741_ (_10417_, _10416_, _10415_);
  and _41742_ (_10418_, _10417_, _05549_);
  or _41743_ (_10419_, _10418_, _10414_);
  and _41744_ (_10421_, _10419_, _09791_);
  or _41745_ (_10422_, _10421_, _10410_);
  and _41746_ (_10423_, _10422_, _05542_);
  or _41747_ (_10424_, _10423_, _10400_);
  and _41748_ (_10425_, _10424_, _09850_);
  and _41749_ (_10426_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _41750_ (_10427_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _41751_ (_10429_, _10427_, _10426_);
  and _41752_ (_10430_, _10429_, _09792_);
  and _41753_ (_10432_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and _41754_ (_10433_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _41755_ (_10435_, _10433_, _10432_);
  and _41756_ (_10436_, _10435_, _05549_);
  or _41757_ (_10437_, _10436_, _10430_);
  and _41758_ (_10438_, _10437_, _05535_);
  and _41759_ (_10439_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _41760_ (_10440_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _41761_ (_10441_, _10440_, _10439_);
  and _41762_ (_10443_, _10441_, _09792_);
  and _41763_ (_10444_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and _41764_ (_10445_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _41765_ (_10447_, _10445_, _10444_);
  and _41766_ (_10448_, _10447_, _05549_);
  or _41767_ (_10449_, _10448_, _10443_);
  and _41768_ (_10450_, _10449_, _09791_);
  or _41769_ (_10451_, _10450_, _10438_);
  and _41770_ (_10452_, _10451_, _09805_);
  or _41771_ (_10453_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _41772_ (_10455_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and _41773_ (_10456_, _10455_, _10453_);
  and _41774_ (_10457_, _10456_, _09792_);
  or _41775_ (_10458_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _41776_ (_10459_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and _41777_ (_10462_, _10459_, _10458_);
  and _41778_ (_10463_, _10462_, _05549_);
  or _41779_ (_10464_, _10463_, _10457_);
  and _41780_ (_10465_, _10464_, _05535_);
  or _41781_ (_10466_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _41782_ (_10467_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and _41783_ (_10468_, _10467_, _10466_);
  and _41784_ (_10469_, _10468_, _09792_);
  or _41785_ (_10470_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _41786_ (_10471_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and _41787_ (_10472_, _10471_, _10470_);
  and _41788_ (_10473_, _10472_, _05549_);
  or _41789_ (_10474_, _10473_, _10469_);
  and _41790_ (_10475_, _10474_, _09791_);
  or _41791_ (_10476_, _10475_, _10465_);
  and _41792_ (_10477_, _10476_, _05542_);
  or _41793_ (_10478_, _10477_, _10452_);
  and _41794_ (_10479_, _10478_, _05518_);
  or _41795_ (_10480_, _10479_, _10425_);
  and _41796_ (_10481_, _10480_, _05520_);
  or _41797_ (_10483_, _10481_, _10376_);
  or _41798_ (_10484_, _10483_, _05526_);
  and _41799_ (_10485_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and _41800_ (_10486_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _41801_ (_10487_, _10486_, _10485_);
  and _41802_ (_10488_, _10487_, _09792_);
  and _41803_ (_10489_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and _41804_ (_10490_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _41805_ (_10491_, _10490_, _10489_);
  and _41806_ (_10492_, _10491_, _05549_);
  or _41807_ (_10493_, _10492_, _10488_);
  or _41808_ (_10494_, _10493_, _09791_);
  and _41809_ (_10495_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and _41810_ (_10496_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _41811_ (_10497_, _10496_, _10495_);
  and _41812_ (_10498_, _10497_, _09792_);
  and _41813_ (_10499_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and _41814_ (_10500_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _41815_ (_10501_, _10500_, _10499_);
  and _41816_ (_10502_, _10501_, _05549_);
  or _41817_ (_10503_, _10502_, _10498_);
  or _41818_ (_10504_, _10503_, _05535_);
  and _41819_ (_10505_, _10504_, _09805_);
  and _41820_ (_10507_, _10505_, _10494_);
  or _41821_ (_10509_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _41822_ (_10510_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and _41823_ (_10511_, _10510_, _05549_);
  and _41824_ (_10512_, _10511_, _10509_);
  or _41825_ (_10514_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _41826_ (_10515_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and _41827_ (_10517_, _10515_, _09792_);
  and _41828_ (_10518_, _10517_, _10514_);
  or _41829_ (_10519_, _10518_, _10512_);
  or _41830_ (_10520_, _10519_, _09791_);
  or _41831_ (_10521_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _41832_ (_10522_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and _41833_ (_10524_, _10522_, _05549_);
  and _41834_ (_10525_, _10524_, _10521_);
  or _41835_ (_10526_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _41836_ (_10527_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and _41837_ (_10529_, _10527_, _09792_);
  and _41838_ (_10530_, _10529_, _10526_);
  or _41839_ (_10531_, _10530_, _10525_);
  or _41840_ (_10532_, _10531_, _05535_);
  and _41841_ (_10533_, _10532_, _05542_);
  and _41842_ (_10535_, _10533_, _10520_);
  or _41843_ (_10536_, _10535_, _10507_);
  and _41844_ (_10537_, _10536_, _09850_);
  and _41845_ (_10538_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _41846_ (_10540_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _41847_ (_10542_, _10540_, _10538_);
  and _41848_ (_10543_, _10542_, _09792_);
  and _41849_ (_10544_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and _41850_ (_10545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or _41851_ (_10546_, _10545_, _10544_);
  and _41852_ (_10547_, _10546_, _05549_);
  or _41853_ (_10548_, _10547_, _10543_);
  or _41854_ (_10549_, _10548_, _09791_);
  and _41855_ (_10550_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _41856_ (_10552_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or _41857_ (_10553_, _10552_, _10550_);
  and _41858_ (_10554_, _10553_, _09792_);
  and _41859_ (_10555_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _41860_ (_10556_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _41861_ (_10557_, _10556_, _10555_);
  and _41862_ (_10558_, _10557_, _05549_);
  or _41863_ (_10559_, _10558_, _10554_);
  or _41864_ (_10561_, _10559_, _05535_);
  and _41865_ (_10563_, _10561_, _09805_);
  and _41866_ (_10564_, _10563_, _10549_);
  or _41867_ (_10566_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or _41868_ (_10567_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and _41869_ (_10568_, _10567_, _10566_);
  and _41870_ (_10570_, _10568_, _09792_);
  or _41871_ (_10571_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _41872_ (_10573_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _41873_ (_10575_, _10573_, _10571_);
  and _41874_ (_10576_, _10575_, _05549_);
  or _41875_ (_10578_, _10576_, _10570_);
  or _41876_ (_10579_, _10578_, _09791_);
  or _41877_ (_10580_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or _41878_ (_10581_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _41879_ (_10582_, _10581_, _10580_);
  and _41880_ (_10584_, _10582_, _09792_);
  or _41881_ (_10585_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _41882_ (_10586_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _41883_ (_10587_, _10586_, _10585_);
  and _41884_ (_10588_, _10587_, _05549_);
  or _41885_ (_10590_, _10588_, _10584_);
  or _41886_ (_10591_, _10590_, _05535_);
  and _41887_ (_10593_, _10591_, _05542_);
  and _41888_ (_10594_, _10593_, _10579_);
  or _41889_ (_10595_, _10594_, _10564_);
  and _41890_ (_10596_, _10595_, _05518_);
  or _41891_ (_10597_, _10596_, _10537_);
  and _41892_ (_10598_, _10597_, _09790_);
  or _41893_ (_10600_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _41894_ (_10602_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and _41895_ (_10603_, _10602_, _10600_);
  and _41896_ (_10604_, _10603_, _09792_);
  or _41897_ (_10605_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or _41898_ (_10606_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _41899_ (_10608_, _10606_, _10605_);
  and _41900_ (_10610_, _10608_, _05549_);
  or _41901_ (_10611_, _10610_, _10604_);
  and _41902_ (_10612_, _10611_, _09791_);
  or _41903_ (_10614_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or _41904_ (_10615_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and _41905_ (_10616_, _10615_, _10614_);
  and _41906_ (_10617_, _10616_, _09792_);
  or _41907_ (_10619_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or _41908_ (_10621_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _41909_ (_10623_, _10621_, _10619_);
  and _41910_ (_10625_, _10623_, _05549_);
  or _41911_ (_10626_, _10625_, _10617_);
  and _41912_ (_10627_, _10626_, _05535_);
  or _41913_ (_10628_, _10627_, _10612_);
  and _41914_ (_10629_, _10628_, _05542_);
  and _41915_ (_10631_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _41916_ (_10632_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _41917_ (_10633_, _10632_, _10631_);
  and _41918_ (_10634_, _10633_, _09792_);
  and _41919_ (_10635_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and _41920_ (_10636_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or _41921_ (_10637_, _10636_, _10635_);
  and _41922_ (_10638_, _10637_, _05549_);
  or _41923_ (_10640_, _10638_, _10634_);
  and _41924_ (_10641_, _10640_, _09791_);
  and _41925_ (_10642_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and _41926_ (_10643_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or _41927_ (_10644_, _10643_, _10642_);
  and _41928_ (_10646_, _10644_, _09792_);
  and _41929_ (_10647_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _41930_ (_10649_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _41931_ (_10651_, _10649_, _10647_);
  and _41932_ (_10652_, _10651_, _05549_);
  or _41933_ (_10654_, _10652_, _10646_);
  and _41934_ (_10655_, _10654_, _05535_);
  or _41935_ (_10657_, _10655_, _10641_);
  and _41936_ (_10659_, _10657_, _09805_);
  or _41937_ (_10660_, _10659_, _10629_);
  and _41938_ (_10661_, _10660_, _05518_);
  or _41939_ (_10662_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _41940_ (_10663_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _41941_ (_10664_, _10663_, _05549_);
  and _41942_ (_10665_, _10664_, _10662_);
  or _41943_ (_10666_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _41944_ (_10667_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and _41945_ (_10669_, _10667_, _09792_);
  and _41946_ (_10670_, _10669_, _10666_);
  or _41947_ (_10672_, _10670_, _10665_);
  and _41948_ (_10673_, _10672_, _09791_);
  or _41949_ (_10674_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _41950_ (_10676_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and _41951_ (_10677_, _10676_, _05549_);
  and _41952_ (_10678_, _10677_, _10674_);
  or _41953_ (_10679_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _41954_ (_10680_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _41955_ (_10682_, _10680_, _09792_);
  and _41956_ (_10683_, _10682_, _10679_);
  or _41957_ (_10684_, _10683_, _10678_);
  and _41958_ (_10685_, _10684_, _05535_);
  or _41959_ (_10687_, _10685_, _10673_);
  and _41960_ (_10689_, _10687_, _05542_);
  and _41961_ (_10691_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and _41962_ (_10693_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _41963_ (_10695_, _10693_, _10691_);
  and _41964_ (_10697_, _10695_, _09792_);
  and _41965_ (_10698_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and _41966_ (_10699_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _41967_ (_10700_, _10699_, _10698_);
  and _41968_ (_10701_, _10700_, _05549_);
  or _41969_ (_10702_, _10701_, _10697_);
  and _41970_ (_10704_, _10702_, _09791_);
  and _41971_ (_10706_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and _41972_ (_10707_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _41973_ (_10708_, _10707_, _10706_);
  and _41974_ (_10709_, _10708_, _09792_);
  and _41975_ (_10710_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and _41976_ (_10712_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _41977_ (_10714_, _10712_, _10710_);
  and _41978_ (_10715_, _10714_, _05549_);
  or _41979_ (_10717_, _10715_, _10709_);
  and _41980_ (_10718_, _10717_, _05535_);
  or _41981_ (_10719_, _10718_, _10704_);
  and _41982_ (_10721_, _10719_, _09805_);
  or _41983_ (_10722_, _10721_, _10689_);
  and _41984_ (_10724_, _10722_, _09850_);
  or _41985_ (_10725_, _10724_, _10661_);
  and _41986_ (_10726_, _10725_, _05520_);
  or _41987_ (_10728_, _10726_, _10598_);
  or _41988_ (_10729_, _10728_, _10033_);
  and _41989_ (_10730_, _10729_, _10484_);
  or _41990_ (_10731_, _10730_, _04413_);
  and _41991_ (_10732_, _10731_, _10274_);
  or _41992_ (_10733_, _10732_, _05563_);
  not _41993_ (_10735_, _05563_);
  or _41994_ (_10737_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _41995_ (_10738_, _10737_, _22731_);
  and _41996_ (_27313_[6], _10738_, _10733_);
  and _41997_ (_10740_, _09774_, _24089_);
  and _41998_ (_10741_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or _41999_ (_03297_, _10741_, _10740_);
  and _42000_ (_10742_, _03026_, _23548_);
  and _42001_ (_10743_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _42002_ (_03300_, _10743_, _10742_);
  and _42003_ (_10744_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and _42004_ (_10745_, _04853_, _23548_);
  or _42005_ (_03321_, _10745_, _10744_);
  and _42006_ (_10746_, _24408_, _24372_);
  and _42007_ (_10748_, _10746_, _24219_);
  not _42008_ (_10749_, _10746_);
  and _42009_ (_10750_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or _42010_ (_03336_, _10750_, _10748_);
  and _42011_ (_10751_, _24408_, _24146_);
  and _42012_ (_10752_, _10751_, _23996_);
  not _42013_ (_10754_, _10751_);
  and _42014_ (_10755_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or _42015_ (_03339_, _10755_, _10752_);
  and _42016_ (_10756_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and _42017_ (_10757_, _04853_, _24219_);
  or _42018_ (_03342_, _10757_, _10756_);
  and _42019_ (_10758_, _10751_, _24089_);
  and _42020_ (_10759_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or _42021_ (_03345_, _10759_, _10758_);
  and _42022_ (_10760_, _10751_, _24219_);
  and _42023_ (_10761_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or _42024_ (_03352_, _10761_, _10760_);
  and _42025_ (_10762_, _24408_, _24140_);
  and _42026_ (_10763_, _10762_, _24134_);
  not _42027_ (_10765_, _10762_);
  and _42028_ (_10766_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _42029_ (_27113_, _10766_, _10763_);
  and _42030_ (_10767_, _10762_, _23548_);
  and _42031_ (_10768_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _42032_ (_27111_, _10768_, _10767_);
  and _42033_ (_10769_, _02512_, _24159_);
  not _42034_ (_10770_, _10769_);
  and _42035_ (_10771_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and _42036_ (_10772_, _10769_, _24219_);
  or _42037_ (_03389_, _10772_, _10771_);
  and _42038_ (_10773_, _02512_, _24297_);
  not _42039_ (_10774_, _10773_);
  and _42040_ (_10775_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and _42041_ (_10776_, _10773_, _23996_);
  or _42042_ (_03399_, _10776_, _10775_);
  and _42043_ (_10777_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _42044_ (_10778_, _10773_, _23583_);
  or _42045_ (_03401_, _10778_, _10777_);
  and _42046_ (_10779_, _09780_, _23548_);
  and _42047_ (_10781_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _42048_ (_03415_, _10781_, _10779_);
  and _42049_ (_10782_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _42050_ (_10783_, _04897_, _23583_);
  or _42051_ (_03418_, _10783_, _10782_);
  and _42052_ (_10784_, _09780_, _24219_);
  and _42053_ (_10785_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _42054_ (_03422_, _10785_, _10784_);
  and _42055_ (_10786_, _05465_, _24134_);
  and _42056_ (_10787_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or _42057_ (_03426_, _10787_, _10786_);
  and _42058_ (_10788_, _02512_, _24016_);
  not _42059_ (_10789_, _10788_);
  and _42060_ (_10790_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and _42061_ (_10791_, _10788_, _23583_);
  or _42062_ (_03427_, _10791_, _10790_);
  and _42063_ (_10792_, _02512_, _24236_);
  not _42064_ (_10793_, _10792_);
  and _42065_ (_10794_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  and _42066_ (_10795_, _10792_, _23996_);
  or _42067_ (_27105_, _10795_, _10794_);
  and _42068_ (_10797_, _09779_, _24297_);
  and _42069_ (_10798_, _10797_, _23996_);
  not _42070_ (_10799_, _10797_);
  and _42071_ (_10800_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or _42072_ (_03440_, _10800_, _10798_);
  and _42073_ (_10801_, _24451_, _23887_);
  and _42074_ (_10802_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _42075_ (_03443_, _10802_, _10801_);
  and _42076_ (_10803_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  and _42077_ (_10804_, _10792_, _24089_);
  or _42078_ (_27104_, _10804_, _10803_);
  and _42079_ (_10805_, _02512_, _23941_);
  not _42080_ (_10806_, _10805_);
  and _42081_ (_10807_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _42082_ (_10808_, _10805_, _23996_);
  or _42083_ (_03456_, _10808_, _10807_);
  and _42084_ (_10809_, _02512_, _24899_);
  not _42085_ (_10811_, _10809_);
  and _42086_ (_10813_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _42087_ (_10815_, _10809_, _23996_);
  or _42088_ (_03467_, _10815_, _10813_);
  and _42089_ (_10816_, _09780_, _24089_);
  and _42090_ (_10817_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _42091_ (_03472_, _10817_, _10816_);
  and _42092_ (_10819_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _42093_ (_10821_, _10809_, _23887_);
  or _42094_ (_03475_, _10821_, _10819_);
  and _42095_ (_10822_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _42096_ (_10823_, _10809_, _24219_);
  or _42097_ (_03477_, _10823_, _10822_);
  and _42098_ (_10824_, _09780_, _23583_);
  and _42099_ (_10825_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _42100_ (_03480_, _10825_, _10824_);
  and _42101_ (_10827_, _02512_, _24474_);
  not _42102_ (_10829_, _10827_);
  and _42103_ (_10830_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  and _42104_ (_10832_, _10827_, _23996_);
  or _42105_ (_03483_, _10832_, _10830_);
  and _42106_ (_10834_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  and _42107_ (_10835_, _10827_, _23548_);
  or _42108_ (_03486_, _10835_, _10834_);
  and _42109_ (_10836_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  and _42110_ (_10837_, _10792_, _23548_);
  or _42111_ (_27101_, _10837_, _10836_);
  and _42112_ (_10839_, _02512_, _24349_);
  not _42113_ (_10840_, _10839_);
  and _42114_ (_10841_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  and _42115_ (_10843_, _10839_, _24134_);
  or _42116_ (_03498_, _10843_, _10841_);
  and _42117_ (_10845_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  and _42118_ (_10846_, _10839_, _23583_);
  or _42119_ (_03507_, _10846_, _10845_);
  and _42120_ (_10847_, _10746_, _23887_);
  and _42121_ (_10848_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or _42122_ (_03509_, _10848_, _10847_);
  and _42123_ (_10849_, _09774_, _23583_);
  and _42124_ (_10850_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or _42125_ (_03511_, _10850_, _10849_);
  and _42126_ (_10851_, _10762_, _23583_);
  and _42127_ (_10852_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _42128_ (_03519_, _10852_, _10851_);
  and _42129_ (_10854_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  and _42130_ (_10855_, _10769_, _24051_);
  or _42131_ (_03529_, _10855_, _10854_);
  and _42132_ (_10856_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  and _42133_ (_10858_, _10769_, _23887_);
  or _42134_ (_03533_, _10858_, _10856_);
  and _42135_ (_10859_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _42136_ (_10860_, _10773_, _24219_);
  or _42137_ (_27108_, _10860_, _10859_);
  and _42138_ (_10861_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and _42139_ (_10862_, _10788_, _24051_);
  or _42140_ (_03539_, _10862_, _10861_);
  and _42141_ (_10863_, _10797_, _23583_);
  and _42142_ (_10865_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  or _42143_ (_27002_, _10865_, _10863_);
  and _42144_ (_10867_, _24140_, _22982_);
  and _42145_ (_10868_, _10867_, _24089_);
  not _42146_ (_10869_, _10867_);
  and _42147_ (_10871_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or _42148_ (_03548_, _10871_, _10868_);
  and _42149_ (_10872_, _10797_, _23887_);
  and _42150_ (_10873_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  or _42151_ (_03553_, _10873_, _10872_);
  and _42152_ (_10874_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and _42153_ (_10875_, _10805_, _23887_);
  or _42154_ (_03560_, _10875_, _10874_);
  and _42155_ (_10876_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  and _42156_ (_10877_, _10827_, _23583_);
  or _42157_ (_03573_, _10877_, _10876_);
  and _42158_ (_10878_, _24302_, _23583_);
  and _42159_ (_10879_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or _42160_ (_03576_, _10879_, _10878_);
  and _42161_ (_10880_, _09670_, _23583_);
  and _42162_ (_10882_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or _42163_ (_03584_, _10882_, _10880_);
  and _42164_ (_10884_, _10762_, _23996_);
  and _42165_ (_10885_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _42166_ (_03598_, _10885_, _10884_);
  and _42167_ (_10887_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and _42168_ (_10888_, _10773_, _24089_);
  or _42169_ (_03605_, _10888_, _10887_);
  and _42170_ (_10889_, _06763_, _24134_);
  and _42171_ (_10890_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _42172_ (_03609_, _10890_, _10889_);
  and _42173_ (_10892_, _10797_, _24134_);
  and _42174_ (_10894_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or _42175_ (_27004_, _10894_, _10892_);
  and _42176_ (_10895_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and _42177_ (_10896_, _10809_, _24089_);
  or _42178_ (_03627_, _10896_, _10895_);
  and _42179_ (_10898_, _10797_, _24051_);
  and _42180_ (_10900_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or _42181_ (_27003_, _10900_, _10898_);
  and _42182_ (_10902_, _10797_, _24089_);
  and _42183_ (_10903_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  or _42184_ (_03631_, _10903_, _10902_);
  and _42185_ (_10904_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _42186_ (_10905_, _06203_, _24051_);
  or _42187_ (_03648_, _10905_, _10904_);
  and _42188_ (_10906_, _09779_, _24016_);
  and _42189_ (_10907_, _10906_, _24089_);
  not _42190_ (_10908_, _10906_);
  and _42191_ (_10909_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or _42192_ (_03659_, _10909_, _10907_);
  and _42193_ (_10911_, _03026_, _24219_);
  and _42194_ (_10912_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _42195_ (_03664_, _10912_, _10911_);
  and _42196_ (_10913_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  and _42197_ (_10914_, _10839_, _23887_);
  or _42198_ (_03671_, _10914_, _10913_);
  and _42199_ (_10916_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and _42200_ (_10917_, _10839_, _24219_);
  or _42201_ (_03673_, _10917_, _10916_);
  and _42202_ (_10919_, _03186_, _23548_);
  and _42203_ (_10920_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or _42204_ (_03675_, _10920_, _10919_);
  and _42205_ (_10922_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  and _42206_ (_10924_, _10839_, _23548_);
  or _42207_ (_27098_, _10924_, _10922_);
  and _42208_ (_10926_, _03186_, _23887_);
  and _42209_ (_10927_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or _42210_ (_27050_, _10927_, _10926_);
  and _42211_ (_10929_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  and _42212_ (_10930_, _10839_, _24089_);
  or _42213_ (_03695_, _10930_, _10929_);
  and _42214_ (_10931_, _10906_, _24134_);
  and _42215_ (_10932_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  or _42216_ (_03697_, _10932_, _10931_);
  and _42217_ (_10935_, _03026_, _24089_);
  and _42218_ (_10937_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _42219_ (_03701_, _10937_, _10935_);
  and _42220_ (_10939_, _03026_, _23887_);
  and _42221_ (_10940_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _42222_ (_03704_, _10940_, _10939_);
  and _42223_ (_10943_, _10906_, _24051_);
  and _42224_ (_10945_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  or _42225_ (_03716_, _10945_, _10943_);
  and _42226_ (_10947_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  and _42227_ (_10949_, _10839_, _24051_);
  or _42228_ (_03718_, _10949_, _10947_);
  and _42229_ (_26841_[1], _26769_, _22731_);
  and _42230_ (_10952_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and _42231_ (_10954_, _10839_, _23996_);
  or _42232_ (_03726_, _10954_, _10952_);
  and _42233_ (_10956_, _02990_, _23887_);
  and _42234_ (_10957_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or _42235_ (_27054_, _10957_, _10956_);
  or _42236_ (_10959_, _02351_, _04800_);
  and _42237_ (_10961_, _10959_, _22737_);
  and _42238_ (_10962_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _42239_ (_10963_, _10962_, _02360_);
  or _42240_ (_10965_, _10963_, _02010_);
  or _42241_ (_10966_, _10965_, _10961_);
  and _42242_ (_26849_[2], _10966_, _22731_);
  and _42243_ (_10969_, _02990_, _24134_);
  and _42244_ (_10971_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or _42245_ (_03741_, _10971_, _10969_);
  and _42246_ (_10972_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and _42247_ (_10973_, _10792_, _24219_);
  or _42248_ (_03749_, _10973_, _10972_);
  and _42249_ (_10975_, _02990_, _24051_);
  and _42250_ (_10977_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or _42251_ (_03753_, _10977_, _10975_);
  and _42252_ (_10979_, _23890_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and _42253_ (_10981_, _23892_, _23779_);
  or _42254_ (_10983_, _09762_, _23923_);
  or _42255_ (_10985_, _10983_, _10981_);
  or _42256_ (_10986_, _23839_, _23793_);
  or _42257_ (_10988_, _10986_, _26739_);
  or _42258_ (_10989_, _10988_, _10985_);
  or _42259_ (_10990_, _10989_, _09753_);
  and _42260_ (_10991_, _10990_, _23855_);
  or _42261_ (_26850_[1], _10991_, _10979_);
  and _42262_ (_10992_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and _42263_ (_10994_, _10827_, _24219_);
  or _42264_ (_03761_, _10994_, _10992_);
  and _42265_ (_10996_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _42266_ (_10997_, _06203_, _24089_);
  or _42267_ (_03766_, _10997_, _10996_);
  and _42268_ (_10998_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and _42269_ (_11000_, _10827_, _23887_);
  or _42270_ (_03768_, _11000_, _10998_);
  and _42271_ (_11002_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  and _42272_ (_11003_, _10827_, _24089_);
  or _42273_ (_03780_, _11003_, _11002_);
  and _42274_ (_11004_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and _42275_ (_11006_, _02338_, _24051_);
  or _42276_ (_27027_, _11006_, _11004_);
  and _42277_ (_11007_, _09717_, _24219_);
  and _42278_ (_11008_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _42279_ (_27070_, _11008_, _11007_);
  and _42280_ (_11009_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  and _42281_ (_11010_, _10827_, _24051_);
  or _42282_ (_03800_, _11010_, _11009_);
  and _42283_ (_11012_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _42284_ (_11013_, _02040_, _24219_);
  or _42285_ (_03804_, _11013_, _11012_);
  and _42286_ (_11015_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _42287_ (_11016_, _02040_, _24134_);
  or _42288_ (_03812_, _11016_, _11015_);
  and _42289_ (_11018_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and _42290_ (_11019_, _10827_, _24134_);
  or _42291_ (_03817_, _11019_, _11018_);
  and _42292_ (_11020_, _10797_, _24219_);
  and _42293_ (_11022_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  or _42294_ (_03820_, _11022_, _11020_);
  and _42295_ (_11025_, _25648_, _24219_);
  and _42296_ (_11026_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or _42297_ (_03827_, _11026_, _11025_);
  and _42298_ (_11028_, _10906_, _23996_);
  and _42299_ (_11029_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  or _42300_ (_03836_, _11029_, _11028_);
  and _42301_ (_11031_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _42302_ (_11032_, _10809_, _23548_);
  or _42303_ (_03848_, _11032_, _11031_);
  and _42304_ (_11033_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _42305_ (_11034_, _06203_, _23583_);
  or _42306_ (_27088_, _11034_, _11033_);
  and _42307_ (_11037_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and _42308_ (_11038_, _10809_, _23583_);
  or _42309_ (_03854_, _11038_, _11037_);
  and _42310_ (_11040_, _25442_, _23548_);
  and _42311_ (_11041_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _42312_ (_03856_, _11041_, _11040_);
  and _42313_ (_11044_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and _42314_ (_11045_, _10809_, _24051_);
  or _42315_ (_03864_, _11045_, _11044_);
  and _42316_ (_11046_, _09779_, _24236_);
  and _42317_ (_11047_, _11046_, _24134_);
  not _42318_ (_11049_, _11046_);
  and _42319_ (_11051_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _42320_ (_03867_, _11051_, _11047_);
  and _42321_ (_11052_, _11046_, _23996_);
  and _42322_ (_11053_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _42323_ (_03900_, _11053_, _11052_);
  and _42324_ (_11054_, _25442_, _24051_);
  and _42325_ (_11055_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _42326_ (_03907_, _11055_, _11054_);
  and _42327_ (_11057_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and _42328_ (_11058_, _10809_, _24134_);
  or _42329_ (_03918_, _11058_, _11057_);
  and _42330_ (_11059_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _42331_ (_11060_, _10805_, _24219_);
  or _42332_ (_03921_, _11060_, _11059_);
  and _42333_ (_11061_, _25206_, _23996_);
  and _42334_ (_11062_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _42335_ (_03924_, _11062_, _11061_);
  and _42336_ (_11063_, _09717_, _23548_);
  and _42337_ (_11064_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _42338_ (_03932_, _11064_, _11063_);
  and _42339_ (_11065_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _42340_ (_11066_, _10805_, _23548_);
  or _42341_ (_03948_, _11066_, _11065_);
  and _42342_ (_11067_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _42343_ (_11069_, _10805_, _23583_);
  or _42344_ (_27097_, _11069_, _11067_);
  and _42345_ (_11070_, _10867_, _24051_);
  and _42346_ (_11072_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or _42347_ (_27262_, _11072_, _11070_);
  and _42348_ (_11073_, _24415_, _23548_);
  and _42349_ (_11075_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or _42350_ (_03961_, _11075_, _11073_);
  and _42351_ (_11078_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _42352_ (_11079_, _10805_, _24089_);
  or _42353_ (_03969_, _11079_, _11078_);
  and _42354_ (_11080_, _24381_, _23548_);
  and _42355_ (_11082_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _42356_ (_03971_, _11082_, _11080_);
  and _42357_ (_11083_, _10906_, _23887_);
  and _42358_ (_11084_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or _42359_ (_03974_, _11084_, _11083_);
  and _42360_ (_11086_, _24415_, _23996_);
  and _42361_ (_11087_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or _42362_ (_03986_, _11087_, _11086_);
  and _42363_ (_11089_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _42364_ (_11090_, _10805_, _24051_);
  or _42365_ (_03989_, _11090_, _11089_);
  or _42366_ (_11092_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and _42367_ (_03992_, _11092_, _03428_);
  and _42368_ (_11093_, _24381_, _23996_);
  and _42369_ (_11094_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _42370_ (_03994_, _11094_, _11093_);
  and _42371_ (_11095_, _10906_, _23548_);
  and _42372_ (_11096_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  or _42373_ (_27001_, _11096_, _11095_);
  and _42374_ (_11097_, _24381_, _24089_);
  and _42375_ (_11098_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _42376_ (_03999_, _11098_, _11097_);
  not _42377_ (_11099_, _02294_);
  or _42378_ (_11100_, _11099_, _23577_);
  and _42379_ (_11101_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _42380_ (_11102_, _02257_, _02248_);
  nor _42381_ (_11104_, _11102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _42382_ (_11105_, _11104_, _06159_);
  and _42383_ (_11107_, _11105_, _06158_);
  and _42384_ (_11108_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _42385_ (_11110_, _11108_, _11107_);
  nor _42386_ (_11112_, _11110_, _02616_);
  or _42387_ (_11114_, _11112_, _11101_);
  or _42388_ (_11116_, _11114_, _02294_);
  and _42389_ (_11118_, _11116_, _22731_);
  and _42390_ (_04002_, _11118_, _11100_);
  and _42391_ (_11119_, _24330_, _24051_);
  and _42392_ (_11120_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _42393_ (_04005_, _11120_, _11119_);
  and _42394_ (_11122_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _42395_ (_11123_, _10805_, _24134_);
  or _42396_ (_04007_, _11123_, _11122_);
  nor _42397_ (_11125_, _24210_, rst);
  or _42398_ (_11127_, _11125_, _02295_);
  and _42399_ (_11129_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _42400_ (_11130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _42401_ (_11131_, _11130_, _02283_);
  and _42402_ (_11132_, _11131_, _02263_);
  and _42403_ (_11134_, _02248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _42404_ (_11136_, _02248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _42405_ (_11137_, _11136_, _11134_);
  and _42406_ (_11138_, _11137_, _06158_);
  nor _42407_ (_11139_, _11138_, _11132_);
  nor _42408_ (_11140_, _11139_, _02616_);
  or _42409_ (_11141_, _11140_, _02294_);
  or _42410_ (_11143_, _11141_, _11129_);
  and _42411_ (_04010_, _11143_, _11127_);
  and _42412_ (_11145_, _10906_, _24219_);
  and _42413_ (_11147_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or _42414_ (_04013_, _11147_, _11145_);
  not _42415_ (_11148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _42416_ (_11149_, _02620_, _02237_);
  and _42417_ (_11150_, _06162_, _02271_);
  nor _42418_ (_11151_, _11150_, _11149_);
  and _42419_ (_11152_, _11151_, _11148_);
  nor _42420_ (_11153_, _11151_, _11148_);
  nor _42421_ (_11154_, _11153_, _11152_);
  or _42422_ (_11155_, _11154_, _02616_);
  nand _42423_ (_11157_, _02616_, _24210_);
  and _42424_ (_11158_, _11157_, _11155_);
  and _42425_ (_11159_, _11158_, _02295_);
  and _42426_ (_11160_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _42427_ (_04015_, _11160_, _11159_);
  and _42428_ (_11163_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  and _42429_ (_11164_, _10792_, _23887_);
  or _42430_ (_27102_, _11164_, _11163_);
  and _42431_ (_11165_, _24350_, _24219_);
  and _42432_ (_11166_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _42433_ (_04026_, _11166_, _11165_);
  or _42434_ (_11168_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _42435_ (_26894_, _11168_, _03087_);
  and _42436_ (_11169_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and _42437_ (_11171_, _10792_, _23583_);
  or _42438_ (_27103_, _11171_, _11169_);
  and _42439_ (_11174_, _24134_, _23946_);
  and _42440_ (_11175_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or _42441_ (_04037_, _11175_, _11174_);
  and _42442_ (_11177_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and _42443_ (_11179_, _10792_, _24051_);
  or _42444_ (_04040_, _11179_, _11177_);
  or _42445_ (_11181_, _02300_, _23577_);
  nand _42446_ (_11182_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _42447_ (_11183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _42448_ (_11184_, _02206_, _02205_);
  and _42449_ (_11185_, _11184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand _42450_ (_11186_, _11185_, _11183_);
  and _42451_ (_11187_, _11186_, _11182_);
  nor _42452_ (_11189_, _11187_, _01814_);
  and _42453_ (_11191_, _02207_, _11184_);
  nand _42454_ (_11193_, _11191_, _02193_);
  and _42455_ (_11194_, _11193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _42456_ (_11195_, _11194_, _11189_);
  or _42457_ (_11196_, _11195_, _01816_);
  and _42458_ (_11198_, _11196_, _22731_);
  and _42459_ (_04044_, _11198_, _11181_);
  or _42460_ (_11201_, _02193_, _23880_);
  and _42461_ (_11203_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _42462_ (_11205_, _11203_, _08224_);
  and _42463_ (_11206_, _11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _42464_ (_11207_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _42465_ (_11208_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _42466_ (_11209_, _11208_, _02197_);
  and _42467_ (_11210_, _11209_, _11207_);
  and _42468_ (_11211_, _02210_, _01820_);
  or _42469_ (_11212_, _11211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _42470_ (_11214_, _11211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _42471_ (_11216_, _11214_, _02320_);
  and _42472_ (_11217_, _11216_, _11212_);
  and _42473_ (_11218_, _01821_, _01818_);
  nand _42474_ (_11219_, _11218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _42475_ (_11221_, _01820_, _01818_);
  and _42476_ (_11223_, _11221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _42477_ (_11225_, _11223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _42478_ (_11226_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _42479_ (_11227_, _11226_, _11219_);
  or _42480_ (_11229_, _11227_, _11217_);
  or _42481_ (_11230_, _11229_, _11210_);
  or _42482_ (_11231_, _11230_, _01814_);
  and _42483_ (_11233_, _11231_, _11201_);
  or _42484_ (_11235_, _11233_, _01816_);
  or _42485_ (_11236_, _02300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _42486_ (_11238_, _11236_, _22731_);
  and _42487_ (_04046_, _11238_, _11235_);
  and _42488_ (_11239_, _24237_, _23887_);
  and _42489_ (_11241_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _42490_ (_04050_, _11241_, _11239_);
  and _42491_ (_11243_, _11046_, _24219_);
  and _42492_ (_11244_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _42493_ (_04055_, _11244_, _11243_);
  and _42494_ (_11245_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  and _42495_ (_11246_, _10792_, _24134_);
  or _42496_ (_04068_, _11246_, _11245_);
  and _42497_ (_11247_, _24237_, _24219_);
  and _42498_ (_11248_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _42499_ (_04072_, _11248_, _11247_);
  and _42500_ (_11250_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _42501_ (_11251_, _10788_, _24219_);
  or _42502_ (_27106_, _11251_, _11250_);
  or _42503_ (_11252_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _42504_ (_04075_, _11252_, _03414_);
  or _42505_ (_11253_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _42506_ (_11254_, _11253_, _22731_);
  not _42507_ (_11256_, _24189_);
  or _42508_ (_11257_, _11256_, _23880_);
  and _42509_ (_04077_, _11257_, _11254_);
  and _42510_ (_11259_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and _42511_ (_11260_, _10788_, _23548_);
  or _42512_ (_04087_, _11260_, _11259_);
  and _42513_ (_11261_, _24017_, _23996_);
  and _42514_ (_11263_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or _42515_ (_04089_, _11263_, _11261_);
  and _42516_ (_11264_, _09779_, _24349_);
  and _42517_ (_11265_, _11264_, _23996_);
  not _42518_ (_11266_, _11264_);
  and _42519_ (_11267_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _42520_ (_04092_, _11267_, _11265_);
  and _42521_ (_11269_, _24089_, _24017_);
  and _42522_ (_11270_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or _42523_ (_04097_, _11270_, _11269_);
  or _42524_ (_11271_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and _42525_ (_04101_, _11271_, _03419_);
  and _42526_ (_11272_, _05465_, _24051_);
  and _42527_ (_11273_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or _42528_ (_04107_, _11273_, _11272_);
  and _42529_ (_11274_, _11264_, _24134_);
  and _42530_ (_11275_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _42531_ (_04109_, _11275_, _11274_);
  and _42532_ (_11276_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _42533_ (_11277_, _10788_, _23887_);
  or _42534_ (_04112_, _11277_, _11276_);
  and _42535_ (_11278_, _05465_, _23583_);
  and _42536_ (_11279_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or _42537_ (_27068_, _11279_, _11278_);
  and _42538_ (_11280_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _42539_ (_11281_, _10788_, _24089_);
  or _42540_ (_04116_, _11281_, _11280_);
  and _42541_ (_11282_, _09717_, _23583_);
  and _42542_ (_11284_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _42543_ (_27071_, _11284_, _11282_);
  and _42544_ (_11286_, _04865_, _23887_);
  and _42545_ (_11288_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or _42546_ (_04126_, _11288_, _11286_);
  and _42547_ (_11290_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and _42548_ (_11291_, _10788_, _24134_);
  or _42549_ (_27107_, _11291_, _11290_);
  and _42550_ (_11293_, _11046_, _23583_);
  and _42551_ (_11295_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _42552_ (_04159_, _11295_, _11293_);
  and _42553_ (_11297_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _42554_ (_11299_, _10788_, _23996_);
  or _42555_ (_04162_, _11299_, _11297_);
  and _42556_ (_11301_, _11046_, _23887_);
  and _42557_ (_11302_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _42558_ (_04165_, _11302_, _11301_);
  and _42559_ (_11304_, _05460_, _24051_);
  and _42560_ (_11306_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _42561_ (_04168_, _11306_, _11304_);
  and _42562_ (_11307_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _42563_ (_11308_, _10773_, _23548_);
  or _42564_ (_04171_, _11308_, _11307_);
  or _42565_ (_11309_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _42566_ (_04174_, _11309_, _03408_);
  and _42567_ (_11311_, _24372_, _24006_);
  and _42568_ (_11312_, _11311_, _24219_);
  not _42569_ (_11313_, _11311_);
  and _42570_ (_11314_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or _42571_ (_04177_, _11314_, _11312_);
  and _42572_ (_11316_, _24442_, _24051_);
  and _42573_ (_11317_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or _42574_ (_27075_, _11317_, _11316_);
  and _42575_ (_11318_, _11046_, _23548_);
  and _42576_ (_11319_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _42577_ (_04185_, _11319_, _11318_);
  and _42578_ (_11320_, _11311_, _23996_);
  and _42579_ (_11321_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or _42580_ (_04187_, _11321_, _11320_);
  and _42581_ (_11323_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _42582_ (_11324_, _10773_, _23887_);
  or _42583_ (_04189_, _11324_, _11323_);
  and _42584_ (_11325_, _11311_, _24089_);
  and _42585_ (_11327_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or _42586_ (_04191_, _11327_, _11325_);
  and _42587_ (_11329_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _42588_ (_11330_, _10773_, _24051_);
  or _42589_ (_04194_, _11330_, _11329_);
  and _42590_ (_11333_, _09717_, _23887_);
  and _42591_ (_11335_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _42592_ (_04198_, _11335_, _11333_);
  and _42593_ (_11337_, _07013_, _24089_);
  and _42594_ (_11338_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _42595_ (_04200_, _11338_, _11337_);
  and _42596_ (_11339_, _24889_, _24089_);
  and _42597_ (_11340_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _42598_ (_04205_, _11340_, _11339_);
  and _42599_ (_11341_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _42600_ (_11342_, _10773_, _24134_);
  or _42601_ (_04208_, _11342_, _11341_);
  and _42602_ (_11343_, _24889_, _23887_);
  and _42603_ (_11344_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _42604_ (_04218_, _11344_, _11343_);
  and _42605_ (_11345_, _09774_, _23996_);
  and _42606_ (_11346_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or _42607_ (_27242_, _11346_, _11345_);
  and _42608_ (_11348_, _08578_, _23548_);
  and _42609_ (_11349_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or _42610_ (_27076_, _11349_, _11348_);
  and _42611_ (_11350_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  and _42612_ (_11351_, _10769_, _23548_);
  or _42613_ (_27109_, _11351_, _11350_);
  and _42614_ (_11353_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  and _42615_ (_11354_, _10769_, _23583_);
  or _42616_ (_04254_, _11354_, _11353_);
  and _42617_ (_11358_, _09774_, _24134_);
  and _42618_ (_11359_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or _42619_ (_04262_, _11359_, _11358_);
  and _42620_ (_11360_, _24056_, _24006_);
  and _42621_ (_11361_, _11360_, _23583_);
  not _42622_ (_11362_, _11360_);
  and _42623_ (_11363_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _42624_ (_04269_, _11363_, _11361_);
  and _42625_ (_11364_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  and _42626_ (_11365_, _10769_, _24089_);
  or _42627_ (_04271_, _11365_, _11364_);
  and _42628_ (_11367_, _11264_, _23548_);
  and _42629_ (_11368_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _42630_ (_04273_, _11368_, _11367_);
  and _42631_ (_11370_, _11264_, _24219_);
  and _42632_ (_11371_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _42633_ (_04279_, _11371_, _11370_);
  and _42634_ (_11373_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and _42635_ (_11374_, _10769_, _24134_);
  or _42636_ (_04282_, _11374_, _11373_);
  and _42637_ (_11376_, _02964_, _23548_);
  and _42638_ (_11377_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _42639_ (_04284_, _11377_, _11376_);
  and _42640_ (_11378_, _11360_, _24134_);
  and _42641_ (_11379_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _42642_ (_04294_, _11379_, _11378_);
  and _42643_ (_11381_, _02964_, _24219_);
  and _42644_ (_11382_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _42645_ (_04296_, _11382_, _11381_);
  and _42646_ (_11384_, _08523_, _23996_);
  and _42647_ (_11385_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or _42648_ (_04299_, _11385_, _11384_);
  and _42649_ (_11386_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  and _42650_ (_11387_, _10769_, _23996_);
  or _42651_ (_27110_, _11387_, _11386_);
  and _42652_ (_11388_, _08523_, _24089_);
  and _42653_ (_11389_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or _42654_ (_04307_, _11389_, _11388_);
  and _42655_ (_11391_, _10762_, _24219_);
  and _42656_ (_11392_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _42657_ (_04310_, _11392_, _11391_);
  and _42658_ (_11393_, _06763_, _23583_);
  and _42659_ (_11394_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _42660_ (_04313_, _11394_, _11393_);
  and _42661_ (_11395_, _10762_, _23887_);
  and _42662_ (_11396_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _42663_ (_04316_, _11396_, _11395_);
  and _42664_ (_11397_, _24089_, _24008_);
  and _42665_ (_11398_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _42666_ (_04318_, _11398_, _11397_);
  and _42667_ (_11399_, _24008_, _23548_);
  and _42668_ (_11400_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _42669_ (_04321_, _11400_, _11399_);
  and _42670_ (_11401_, _10762_, _24089_);
  and _42671_ (_11402_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _42672_ (_04324_, _11402_, _11401_);
  and _42673_ (_11403_, _02488_, _23583_);
  and _42674_ (_11404_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or _42675_ (_04346_, _11404_, _11403_);
  and _42676_ (_11405_, _02964_, _24134_);
  and _42677_ (_11406_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _42678_ (_04351_, _11406_, _11405_);
  and _42679_ (_11409_, _02065_, _23887_);
  and _42680_ (_11410_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or _42681_ (_04354_, _11410_, _11409_);
  and _42682_ (_11412_, _10762_, _24051_);
  and _42683_ (_11413_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _42684_ (_27112_, _11413_, _11412_);
  and _42685_ (_11414_, _02488_, _23996_);
  and _42686_ (_11415_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or _42687_ (_04359_, _11415_, _11414_);
  and _42688_ (_11417_, _05442_, _23887_);
  and _42689_ (_11418_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _42690_ (_04365_, _11418_, _11417_);
  and _42691_ (_11419_, _24016_, _24006_);
  and _42692_ (_11420_, _11419_, _23548_);
  not _42693_ (_11421_, _11419_);
  and _42694_ (_11422_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _42695_ (_04369_, _11422_, _11420_);
  and _42696_ (_11423_, _05442_, _24089_);
  and _42697_ (_11424_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _42698_ (_04371_, _11424_, _11423_);
  and _42699_ (_11426_, _10751_, _23548_);
  and _42700_ (_11427_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or _42701_ (_04381_, _11427_, _11426_);
  and _42702_ (_11428_, _11264_, _24089_);
  and _42703_ (_11429_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _42704_ (_04386_, _11429_, _11428_);
  and _42705_ (_11430_, _02964_, _24089_);
  and _42706_ (_11431_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _42707_ (_04391_, _11431_, _11430_);
  and _42708_ (_11432_, _11264_, _23583_);
  and _42709_ (_11433_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _42710_ (_26999_, _11433_, _11432_);
  and _42711_ (_11434_, _11419_, _24051_);
  and _42712_ (_11435_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _42713_ (_04398_, _11435_, _11434_);
  and _42714_ (_11437_, _10751_, _23887_);
  and _42715_ (_11438_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or _42716_ (_27114_, _11438_, _11437_);
  and _42717_ (_11441_, _24297_, _24006_);
  and _42718_ (_11443_, _11441_, _24089_);
  not _42719_ (_11444_, _11441_);
  and _42720_ (_11445_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _42721_ (_04408_, _11445_, _11443_);
  and _42722_ (_11447_, _02964_, _23583_);
  and _42723_ (_11448_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _42724_ (_04411_, _11448_, _11447_);
  and _42725_ (_11449_, _02964_, _23887_);
  and _42726_ (_11451_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _42727_ (_04415_, _11451_, _11449_);
  and _42728_ (_11453_, _11441_, _23548_);
  and _42729_ (_11454_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _42730_ (_04417_, _11454_, _11453_);
  and _42731_ (_11456_, _23922_, _22737_);
  and _42732_ (_11457_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _42733_ (_11458_, _11457_, _26680_);
  or _42734_ (_11459_, _11458_, _11456_);
  and _42735_ (_26852_[1], _11459_, _22731_);
  and _42736_ (_11460_, _06763_, _24051_);
  and _42737_ (_11461_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or _42738_ (_04422_, _11461_, _11460_);
  and _42739_ (_11464_, _10751_, _23583_);
  and _42740_ (_11465_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or _42741_ (_04424_, _11465_, _11464_);
  and _42742_ (_11467_, _11264_, _23887_);
  and _42743_ (_11468_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _42744_ (_26998_, _11468_, _11467_);
  and _42745_ (_11469_, _08435_, _24219_);
  and _42746_ (_11470_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or _42747_ (_04432_, _11470_, _11469_);
  and _42748_ (_11471_, _23890_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or _42749_ (_11472_, _23819_, _23809_);
  or _42750_ (_11473_, _04789_, _23929_);
  or _42751_ (_11474_, _11473_, _23836_);
  or _42752_ (_11476_, _11474_, _23828_);
  or _42753_ (_11477_, _11476_, _03919_);
  or _42754_ (_11478_, _04796_, _26731_);
  or _42755_ (_11479_, _11478_, _24276_);
  or _42756_ (_11480_, _11479_, _24262_);
  or _42757_ (_11481_, _11480_, _11477_);
  or _42758_ (_11482_, _11481_, _11472_);
  and _42759_ (_11483_, _11482_, _23855_);
  or _42760_ (_26851_[3], _11483_, _11471_);
  and _42761_ (_11484_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _42762_ (_11485_, _06203_, _24219_);
  or _42763_ (_04445_, _11485_, _11484_);
  and _42764_ (_11488_, _10751_, _24051_);
  and _42765_ (_11489_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or _42766_ (_27115_, _11489_, _11488_);
  and _42767_ (_11490_, _05438_, _23548_);
  and _42768_ (_11491_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _42769_ (_04453_, _11491_, _11490_);
  and _42770_ (_11492_, _10751_, _24134_);
  and _42771_ (_11493_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or _42772_ (_04455_, _11493_, _11492_);
  and _42773_ (_11494_, _05438_, _23887_);
  and _42774_ (_11495_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _42775_ (_04457_, _11495_, _11494_);
  and _42776_ (_11497_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and _42777_ (_11498_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _42778_ (_11499_, _11498_, _11497_);
  and _42779_ (_11500_, _11499_, _09792_);
  and _42780_ (_11501_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and _42781_ (_11502_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _42782_ (_11503_, _11502_, _11501_);
  and _42783_ (_11504_, _11503_, _05549_);
  or _42784_ (_11505_, _11504_, _11500_);
  or _42785_ (_11506_, _11505_, _09791_);
  and _42786_ (_11507_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and _42787_ (_11508_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _42788_ (_11509_, _11508_, _11507_);
  and _42789_ (_11511_, _11509_, _09792_);
  and _42790_ (_11513_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and _42791_ (_11515_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _42792_ (_11516_, _11515_, _11513_);
  and _42793_ (_11518_, _11516_, _05549_);
  or _42794_ (_11520_, _11518_, _11511_);
  or _42795_ (_11521_, _11520_, _05535_);
  and _42796_ (_11522_, _11521_, _09805_);
  and _42797_ (_11523_, _11522_, _11506_);
  or _42798_ (_11524_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _42799_ (_11525_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and _42800_ (_11527_, _11525_, _11524_);
  and _42801_ (_11529_, _11527_, _09792_);
  or _42802_ (_11530_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _42803_ (_11531_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and _42804_ (_11532_, _11531_, _11530_);
  and _42805_ (_11533_, _11532_, _05549_);
  or _42806_ (_11534_, _11533_, _11529_);
  or _42807_ (_11535_, _11534_, _09791_);
  or _42808_ (_11536_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _42809_ (_11537_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and _42810_ (_11538_, _11537_, _11536_);
  and _42811_ (_11540_, _11538_, _09792_);
  or _42812_ (_11541_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _42813_ (_11542_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and _42814_ (_11543_, _11542_, _11541_);
  and _42815_ (_11544_, _11543_, _05549_);
  or _42816_ (_11545_, _11544_, _11540_);
  or _42817_ (_11546_, _11545_, _05535_);
  and _42818_ (_11547_, _11546_, _05542_);
  and _42819_ (_11548_, _11547_, _11535_);
  or _42820_ (_11549_, _11548_, _11523_);
  and _42821_ (_11551_, _11549_, _05518_);
  and _42822_ (_11552_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and _42823_ (_11554_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _42824_ (_11555_, _11554_, _11552_);
  and _42825_ (_11556_, _11555_, _09792_);
  and _42826_ (_11557_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and _42827_ (_11558_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _42828_ (_11559_, _11558_, _11557_);
  and _42829_ (_11560_, _11559_, _05549_);
  or _42830_ (_11561_, _11560_, _11556_);
  or _42831_ (_11562_, _11561_, _09791_);
  and _42832_ (_11564_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and _42833_ (_11565_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _42834_ (_11566_, _11565_, _11564_);
  and _42835_ (_11567_, _11566_, _09792_);
  and _42836_ (_11568_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and _42837_ (_11569_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _42838_ (_11570_, _11569_, _11568_);
  and _42839_ (_11571_, _11570_, _05549_);
  or _42840_ (_11572_, _11571_, _11567_);
  or _42841_ (_11573_, _11572_, _05535_);
  and _42842_ (_11574_, _11573_, _09805_);
  and _42843_ (_11575_, _11574_, _11562_);
  or _42844_ (_11576_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _42845_ (_11577_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and _42846_ (_11578_, _11577_, _05549_);
  and _42847_ (_11579_, _11578_, _11576_);
  or _42848_ (_11580_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _42849_ (_11581_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and _42850_ (_11582_, _11581_, _09792_);
  and _42851_ (_11583_, _11582_, _11580_);
  or _42852_ (_11584_, _11583_, _11579_);
  or _42853_ (_11585_, _11584_, _09791_);
  or _42854_ (_11586_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _42855_ (_11587_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and _42856_ (_11588_, _11587_, _05549_);
  and _42857_ (_11590_, _11588_, _11586_);
  or _42858_ (_11591_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _42859_ (_11593_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and _42860_ (_11595_, _11593_, _09792_);
  and _42861_ (_11597_, _11595_, _11591_);
  or _42862_ (_11598_, _11597_, _11590_);
  or _42863_ (_11599_, _11598_, _05535_);
  and _42864_ (_11600_, _11599_, _05542_);
  and _42865_ (_11602_, _11600_, _11585_);
  or _42866_ (_11604_, _11602_, _11575_);
  and _42867_ (_11606_, _11604_, _09850_);
  or _42868_ (_11607_, _11606_, _11551_);
  and _42869_ (_11608_, _11607_, _09790_);
  and _42870_ (_11609_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and _42871_ (_11610_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _42872_ (_11612_, _11610_, _11609_);
  and _42873_ (_11613_, _11612_, _09792_);
  and _42874_ (_11615_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _42875_ (_11616_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _42876_ (_11617_, _11616_, _11615_);
  and _42877_ (_11619_, _11617_, _05549_);
  or _42878_ (_11620_, _11619_, _11613_);
  and _42879_ (_11621_, _11620_, _05535_);
  and _42880_ (_11622_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _42881_ (_11623_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _42882_ (_11624_, _11623_, _11622_);
  and _42883_ (_11625_, _11624_, _09792_);
  and _42884_ (_11626_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and _42885_ (_11628_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _42886_ (_11629_, _11628_, _11626_);
  and _42887_ (_11631_, _11629_, _05549_);
  or _42888_ (_11633_, _11631_, _11625_);
  and _42889_ (_11634_, _11633_, _09791_);
  or _42890_ (_11635_, _11634_, _11621_);
  and _42891_ (_11636_, _11635_, _09805_);
  or _42892_ (_11637_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _42893_ (_11639_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _42894_ (_11640_, _11639_, _05549_);
  and _42895_ (_11642_, _11640_, _11637_);
  or _42896_ (_11643_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _42897_ (_11645_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _42898_ (_11646_, _11645_, _09792_);
  and _42899_ (_11647_, _11646_, _11643_);
  or _42900_ (_11648_, _11647_, _11642_);
  and _42901_ (_11649_, _11648_, _05535_);
  or _42902_ (_11650_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _42903_ (_11651_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _42904_ (_11652_, _11651_, _05549_);
  and _42905_ (_11653_, _11652_, _11650_);
  or _42906_ (_11655_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _42907_ (_11657_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _42908_ (_11659_, _11657_, _09792_);
  and _42909_ (_11660_, _11659_, _11655_);
  or _42910_ (_11662_, _11660_, _11653_);
  and _42911_ (_11663_, _11662_, _09791_);
  or _42912_ (_11664_, _11663_, _11649_);
  and _42913_ (_11665_, _11664_, _05542_);
  or _42914_ (_11666_, _11665_, _11636_);
  and _42915_ (_11667_, _11666_, _09850_);
  and _42916_ (_11668_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and _42917_ (_11670_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _42918_ (_11671_, _11670_, _11668_);
  and _42919_ (_11672_, _11671_, _09792_);
  and _42920_ (_11673_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and _42921_ (_11674_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _42922_ (_11675_, _11674_, _11673_);
  and _42923_ (_11676_, _11675_, _05549_);
  or _42924_ (_11677_, _11676_, _11672_);
  and _42925_ (_11678_, _11677_, _05535_);
  and _42926_ (_11679_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and _42927_ (_11680_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _42928_ (_11681_, _11680_, _11679_);
  and _42929_ (_11682_, _11681_, _09792_);
  and _42930_ (_11683_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and _42931_ (_11684_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _42932_ (_11686_, _11684_, _11683_);
  and _42933_ (_11687_, _11686_, _05549_);
  or _42934_ (_11689_, _11687_, _11682_);
  and _42935_ (_11690_, _11689_, _09791_);
  or _42936_ (_11692_, _11690_, _11678_);
  and _42937_ (_11693_, _11692_, _09805_);
  or _42938_ (_11695_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _42939_ (_11697_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and _42940_ (_11698_, _11697_, _11695_);
  and _42941_ (_11700_, _11698_, _09792_);
  or _42942_ (_11701_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _42943_ (_11702_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and _42944_ (_11703_, _11702_, _11701_);
  and _42945_ (_11704_, _11703_, _05549_);
  or _42946_ (_11705_, _11704_, _11700_);
  and _42947_ (_11706_, _11705_, _05535_);
  or _42948_ (_11707_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _42949_ (_11709_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and _42950_ (_11710_, _11709_, _11707_);
  and _42951_ (_11712_, _11710_, _09792_);
  or _42952_ (_11713_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _42953_ (_11715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and _42954_ (_11717_, _11715_, _11713_);
  and _42955_ (_11718_, _11717_, _05549_);
  or _42956_ (_11719_, _11718_, _11712_);
  and _42957_ (_11720_, _11719_, _09791_);
  or _42958_ (_11722_, _11720_, _11706_);
  and _42959_ (_11724_, _11722_, _05542_);
  or _42960_ (_11725_, _11724_, _11693_);
  and _42961_ (_11727_, _11725_, _05518_);
  or _42962_ (_11729_, _11727_, _11667_);
  and _42963_ (_11731_, _11729_, _05520_);
  or _42964_ (_11732_, _11731_, _11608_);
  or _42965_ (_11733_, _11732_, _05526_);
  and _42966_ (_11735_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and _42967_ (_11737_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _42968_ (_11739_, _11737_, _11735_);
  and _42969_ (_11741_, _11739_, _09792_);
  and _42970_ (_11743_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and _42971_ (_11744_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _42972_ (_11745_, _11744_, _11743_);
  and _42973_ (_11747_, _11745_, _05549_);
  or _42974_ (_11748_, _11747_, _11741_);
  or _42975_ (_11749_, _11748_, _09791_);
  and _42976_ (_11751_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and _42977_ (_11753_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _42978_ (_11755_, _11753_, _11751_);
  and _42979_ (_11756_, _11755_, _09792_);
  and _42980_ (_11758_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and _42981_ (_11760_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _42982_ (_11762_, _11760_, _11758_);
  and _42983_ (_11763_, _11762_, _05549_);
  or _42984_ (_11764_, _11763_, _11756_);
  or _42985_ (_11765_, _11764_, _05535_);
  and _42986_ (_11766_, _11765_, _09805_);
  and _42987_ (_11767_, _11766_, _11749_);
  or _42988_ (_11768_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _42989_ (_11769_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and _42990_ (_11770_, _11769_, _05549_);
  and _42991_ (_11771_, _11770_, _11768_);
  or _42992_ (_11772_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _42993_ (_11773_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and _42994_ (_11774_, _11773_, _09792_);
  and _42995_ (_11775_, _11774_, _11772_);
  or _42996_ (_11777_, _11775_, _11771_);
  or _42997_ (_11779_, _11777_, _09791_);
  or _42998_ (_11780_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _42999_ (_11781_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and _43000_ (_11782_, _11781_, _05549_);
  and _43001_ (_11783_, _11782_, _11780_);
  or _43002_ (_11784_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _43003_ (_11785_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and _43004_ (_11786_, _11785_, _09792_);
  and _43005_ (_11787_, _11786_, _11784_);
  or _43006_ (_11788_, _11787_, _11783_);
  or _43007_ (_11789_, _11788_, _05535_);
  and _43008_ (_11790_, _11789_, _05542_);
  and _43009_ (_11791_, _11790_, _11779_);
  or _43010_ (_11793_, _11791_, _11767_);
  and _43011_ (_11794_, _11793_, _09850_);
  and _43012_ (_11796_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _43013_ (_11797_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _43014_ (_11798_, _11797_, _11796_);
  and _43015_ (_11799_, _11798_, _09792_);
  and _43016_ (_11800_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and _43017_ (_11801_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _43018_ (_11802_, _11801_, _11800_);
  and _43019_ (_11803_, _11802_, _05549_);
  or _43020_ (_11804_, _11803_, _11799_);
  or _43021_ (_11805_, _11804_, _09791_);
  and _43022_ (_11806_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and _43023_ (_11807_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _43024_ (_11808_, _11807_, _11806_);
  and _43025_ (_11809_, _11808_, _09792_);
  and _43026_ (_11810_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and _43027_ (_11811_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _43028_ (_11812_, _11811_, _11810_);
  and _43029_ (_11813_, _11812_, _05549_);
  or _43030_ (_11814_, _11813_, _11809_);
  or _43031_ (_11815_, _11814_, _05535_);
  and _43032_ (_11816_, _11815_, _09805_);
  and _43033_ (_11817_, _11816_, _11805_);
  or _43034_ (_11818_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _43035_ (_11819_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and _43036_ (_11820_, _11819_, _11818_);
  and _43037_ (_11821_, _11820_, _09792_);
  or _43038_ (_11822_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _43039_ (_11823_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and _43040_ (_11824_, _11823_, _11822_);
  and _43041_ (_11825_, _11824_, _05549_);
  or _43042_ (_11826_, _11825_, _11821_);
  or _43043_ (_11827_, _11826_, _09791_);
  or _43044_ (_11828_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _43045_ (_11829_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and _43046_ (_11830_, _11829_, _11828_);
  and _43047_ (_11831_, _11830_, _09792_);
  or _43048_ (_11832_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _43049_ (_11833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and _43050_ (_11834_, _11833_, _11832_);
  and _43051_ (_11835_, _11834_, _05549_);
  or _43052_ (_11836_, _11835_, _11831_);
  or _43053_ (_11837_, _11836_, _05535_);
  and _43054_ (_11838_, _11837_, _05542_);
  and _43055_ (_11839_, _11838_, _11827_);
  or _43056_ (_11840_, _11839_, _11817_);
  and _43057_ (_11841_, _11840_, _05518_);
  or _43058_ (_11842_, _11841_, _11794_);
  and _43059_ (_11843_, _11842_, _09790_);
  or _43060_ (_11844_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _43061_ (_11845_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and _43062_ (_11846_, _11845_, _11844_);
  and _43063_ (_11847_, _11846_, _09792_);
  or _43064_ (_11848_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _43065_ (_11849_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and _43066_ (_11850_, _11849_, _11848_);
  and _43067_ (_11851_, _11850_, _05549_);
  or _43068_ (_11852_, _11851_, _11847_);
  and _43069_ (_11853_, _11852_, _09791_);
  or _43070_ (_11854_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _43071_ (_11855_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and _43072_ (_11856_, _11855_, _11854_);
  and _43073_ (_11857_, _11856_, _09792_);
  or _43074_ (_11858_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _43075_ (_11859_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and _43076_ (_11860_, _11859_, _11858_);
  and _43077_ (_11861_, _11860_, _05549_);
  or _43078_ (_11862_, _11861_, _11857_);
  and _43079_ (_11863_, _11862_, _05535_);
  or _43080_ (_11864_, _11863_, _11853_);
  and _43081_ (_11865_, _11864_, _05542_);
  and _43082_ (_11866_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and _43083_ (_11867_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _43084_ (_11868_, _11867_, _11866_);
  and _43085_ (_11869_, _11868_, _09792_);
  and _43086_ (_11870_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and _43087_ (_11871_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _43088_ (_11872_, _11871_, _11870_);
  and _43089_ (_11873_, _11872_, _05549_);
  or _43090_ (_11874_, _11873_, _11869_);
  and _43091_ (_11875_, _11874_, _09791_);
  and _43092_ (_11876_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and _43093_ (_11877_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _43094_ (_11878_, _11877_, _11876_);
  and _43095_ (_11879_, _11878_, _09792_);
  and _43096_ (_11880_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and _43097_ (_11881_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _43098_ (_11882_, _11881_, _11880_);
  and _43099_ (_11883_, _11882_, _05549_);
  or _43100_ (_11884_, _11883_, _11879_);
  and _43101_ (_11885_, _11884_, _05535_);
  or _43102_ (_11886_, _11885_, _11875_);
  and _43103_ (_11887_, _11886_, _09805_);
  or _43104_ (_11888_, _11887_, _11865_);
  and _43105_ (_11889_, _11888_, _05518_);
  or _43106_ (_11890_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or _43107_ (_11892_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and _43108_ (_11893_, _11892_, _05549_);
  and _43109_ (_11894_, _11893_, _11890_);
  or _43110_ (_11895_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _43111_ (_11896_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and _43112_ (_11897_, _11896_, _09792_);
  and _43113_ (_11898_, _11897_, _11895_);
  or _43114_ (_11899_, _11898_, _11894_);
  and _43115_ (_11900_, _11899_, _09791_);
  or _43116_ (_11901_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or _43117_ (_11903_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and _43118_ (_11904_, _11903_, _05549_);
  and _43119_ (_11905_, _11904_, _11901_);
  or _43120_ (_11907_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _43121_ (_11908_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and _43122_ (_11910_, _11908_, _09792_);
  and _43123_ (_11911_, _11910_, _11907_);
  or _43124_ (_11912_, _11911_, _11905_);
  and _43125_ (_11913_, _11912_, _05535_);
  or _43126_ (_11915_, _11913_, _11900_);
  and _43127_ (_11917_, _11915_, _05542_);
  and _43128_ (_11918_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and _43129_ (_11919_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _43130_ (_11921_, _11919_, _11918_);
  and _43131_ (_11922_, _11921_, _09792_);
  and _43132_ (_11923_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and _43133_ (_11924_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _43134_ (_11926_, _11924_, _11923_);
  and _43135_ (_11928_, _11926_, _05549_);
  or _43136_ (_11929_, _11928_, _11922_);
  and _43137_ (_11930_, _11929_, _09791_);
  and _43138_ (_11931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and _43139_ (_11933_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _43140_ (_11935_, _11933_, _11931_);
  and _43141_ (_11936_, _11935_, _09792_);
  and _43142_ (_11938_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and _43143_ (_11939_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _43144_ (_11940_, _11939_, _11938_);
  and _43145_ (_11941_, _11940_, _05549_);
  or _43146_ (_11942_, _11941_, _11936_);
  and _43147_ (_11943_, _11942_, _05535_);
  or _43148_ (_11944_, _11943_, _11930_);
  and _43149_ (_11945_, _11944_, _09805_);
  or _43150_ (_11946_, _11945_, _11917_);
  and _43151_ (_11947_, _11946_, _09850_);
  or _43152_ (_11948_, _11947_, _11889_);
  and _43153_ (_11949_, _11948_, _05520_);
  or _43154_ (_11950_, _11949_, _11843_);
  or _43155_ (_11951_, _11950_, _10033_);
  and _43156_ (_11952_, _11951_, _11733_);
  or _43157_ (_11953_, _11952_, _00143_);
  and _43158_ (_11954_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and _43159_ (_11955_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _43160_ (_11956_, _11955_, _11954_);
  and _43161_ (_11957_, _11956_, _09792_);
  and _43162_ (_11958_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and _43163_ (_11959_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _43164_ (_11960_, _11959_, _11958_);
  and _43165_ (_11961_, _11960_, _05549_);
  or _43166_ (_11962_, _11961_, _11957_);
  or _43167_ (_11963_, _11962_, _09791_);
  and _43168_ (_11964_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and _43169_ (_11965_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _43170_ (_11966_, _11965_, _11964_);
  and _43171_ (_11967_, _11966_, _09792_);
  and _43172_ (_11968_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and _43173_ (_11969_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _43174_ (_11970_, _11969_, _11968_);
  and _43175_ (_11971_, _11970_, _05549_);
  or _43176_ (_11972_, _11971_, _11967_);
  or _43177_ (_11974_, _11972_, _05535_);
  and _43178_ (_11975_, _11974_, _09805_);
  and _43179_ (_11976_, _11975_, _11963_);
  or _43180_ (_11977_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _43181_ (_11978_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and _43182_ (_11979_, _11978_, _11977_);
  and _43183_ (_11980_, _11979_, _09792_);
  or _43184_ (_11981_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _43185_ (_11982_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and _43186_ (_11983_, _11982_, _11981_);
  and _43187_ (_11984_, _11983_, _05549_);
  or _43188_ (_11985_, _11984_, _11980_);
  or _43189_ (_11986_, _11985_, _09791_);
  or _43190_ (_11987_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _43191_ (_11988_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and _43192_ (_11989_, _11988_, _11987_);
  and _43193_ (_11990_, _11989_, _09792_);
  or _43194_ (_11991_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _43195_ (_11992_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and _43196_ (_11993_, _11992_, _11991_);
  and _43197_ (_11995_, _11993_, _05549_);
  or _43198_ (_11996_, _11995_, _11990_);
  or _43199_ (_11997_, _11996_, _05535_);
  and _43200_ (_11998_, _11997_, _05542_);
  and _43201_ (_11999_, _11998_, _11986_);
  or _43202_ (_12000_, _11999_, _11976_);
  and _43203_ (_12001_, _12000_, _05518_);
  and _43204_ (_12002_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _43205_ (_12003_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _43206_ (_12004_, _12003_, _12002_);
  and _43207_ (_12005_, _12004_, _09792_);
  and _43208_ (_12006_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _43209_ (_12007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or _43210_ (_12008_, _12007_, _12006_);
  and _43211_ (_12009_, _12008_, _05549_);
  or _43212_ (_12010_, _12009_, _12005_);
  or _43213_ (_12011_, _12010_, _09791_);
  and _43214_ (_12012_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _43215_ (_12013_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _43216_ (_12014_, _12013_, _12012_);
  and _43217_ (_12015_, _12014_, _09792_);
  and _43218_ (_12016_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _43219_ (_12017_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _43220_ (_12018_, _12017_, _12016_);
  and _43221_ (_12019_, _12018_, _05549_);
  or _43222_ (_12020_, _12019_, _12015_);
  or _43223_ (_12021_, _12020_, _05535_);
  and _43224_ (_12022_, _12021_, _09805_);
  and _43225_ (_12023_, _12022_, _12011_);
  or _43226_ (_12024_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _43227_ (_12025_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _43228_ (_12026_, _12025_, _05549_);
  and _43229_ (_12027_, _12026_, _12024_);
  or _43230_ (_12028_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or _43231_ (_12029_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _43232_ (_12030_, _12029_, _09792_);
  and _43233_ (_12031_, _12030_, _12028_);
  or _43234_ (_12032_, _12031_, _12027_);
  or _43235_ (_12033_, _12032_, _09791_);
  or _43236_ (_12034_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _43237_ (_12035_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _43238_ (_12036_, _12035_, _05549_);
  and _43239_ (_12037_, _12036_, _12034_);
  or _43240_ (_12038_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or _43241_ (_12039_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _43242_ (_12040_, _12039_, _09792_);
  and _43243_ (_12041_, _12040_, _12038_);
  or _43244_ (_12042_, _12041_, _12037_);
  or _43245_ (_12043_, _12042_, _05535_);
  and _43246_ (_12044_, _12043_, _05542_);
  and _43247_ (_12045_, _12044_, _12033_);
  or _43248_ (_12046_, _12045_, _12023_);
  and _43249_ (_12047_, _12046_, _09850_);
  or _43250_ (_12048_, _12047_, _12001_);
  and _43251_ (_12049_, _12048_, _09790_);
  and _43252_ (_12050_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _43253_ (_12051_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or _43254_ (_12052_, _12051_, _12050_);
  and _43255_ (_12053_, _12052_, _09792_);
  and _43256_ (_12054_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _43257_ (_12055_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _43258_ (_12056_, _12055_, _12054_);
  and _43259_ (_12057_, _12056_, _05549_);
  or _43260_ (_12058_, _12057_, _12053_);
  and _43261_ (_12059_, _12058_, _05535_);
  and _43262_ (_12060_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _43263_ (_12061_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or _43264_ (_12062_, _12061_, _12060_);
  and _43265_ (_12063_, _12062_, _09792_);
  and _43266_ (_12064_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _43267_ (_12066_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or _43268_ (_12067_, _12066_, _12064_);
  and _43269_ (_12068_, _12067_, _05549_);
  or _43270_ (_12069_, _12068_, _12063_);
  and _43271_ (_12070_, _12069_, _09791_);
  or _43272_ (_12071_, _12070_, _12059_);
  and _43273_ (_12072_, _12071_, _09805_);
  or _43274_ (_12073_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _43275_ (_12074_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _43276_ (_12075_, _12074_, _05549_);
  and _43277_ (_12076_, _12075_, _12073_);
  or _43278_ (_12077_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _43279_ (_12078_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and _43280_ (_12079_, _12078_, _09792_);
  and _43281_ (_12080_, _12079_, _12077_);
  or _43282_ (_12081_, _12080_, _12076_);
  and _43283_ (_12082_, _12081_, _05535_);
  or _43284_ (_12083_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _43285_ (_12084_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _43286_ (_12085_, _12084_, _05549_);
  and _43287_ (_12086_, _12085_, _12083_);
  or _43288_ (_12087_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or _43289_ (_12088_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _43290_ (_12089_, _12088_, _09792_);
  and _43291_ (_12090_, _12089_, _12087_);
  or _43292_ (_12091_, _12090_, _12086_);
  and _43293_ (_12093_, _12091_, _09791_);
  or _43294_ (_12094_, _12093_, _12082_);
  and _43295_ (_12095_, _12094_, _05542_);
  or _43296_ (_12096_, _12095_, _12072_);
  and _43297_ (_12097_, _12096_, _09850_);
  and _43298_ (_12098_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and _43299_ (_12099_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _43300_ (_12100_, _12099_, _12098_);
  and _43301_ (_12101_, _12100_, _09792_);
  and _43302_ (_12102_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and _43303_ (_12103_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _43304_ (_12104_, _12103_, _12102_);
  and _43305_ (_12105_, _12104_, _05549_);
  or _43306_ (_12106_, _12105_, _12101_);
  and _43307_ (_12107_, _12106_, _05535_);
  and _43308_ (_12108_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and _43309_ (_12109_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _43310_ (_12110_, _12109_, _12108_);
  and _43311_ (_12111_, _12110_, _09792_);
  and _43312_ (_12112_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _43313_ (_12113_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _43314_ (_12114_, _12113_, _12112_);
  and _43315_ (_12115_, _12114_, _05549_);
  or _43316_ (_12116_, _12115_, _12111_);
  and _43317_ (_12117_, _12116_, _09791_);
  or _43318_ (_12118_, _12117_, _12107_);
  and _43319_ (_12119_, _12118_, _09805_);
  or _43320_ (_12120_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _43321_ (_12121_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _43322_ (_12122_, _12121_, _12120_);
  and _43323_ (_12123_, _12122_, _09792_);
  or _43324_ (_12124_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _43325_ (_12125_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and _43326_ (_12126_, _12125_, _12124_);
  and _43327_ (_12127_, _12126_, _05549_);
  or _43328_ (_12128_, _12127_, _12123_);
  and _43329_ (_12129_, _12128_, _05535_);
  or _43330_ (_12130_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _43331_ (_12131_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _43332_ (_12132_, _12131_, _12130_);
  and _43333_ (_12133_, _12132_, _09792_);
  or _43334_ (_12134_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _43335_ (_12135_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and _43336_ (_12136_, _12135_, _12134_);
  and _43337_ (_12137_, _12136_, _05549_);
  or _43338_ (_12138_, _12137_, _12133_);
  and _43339_ (_12139_, _12138_, _09791_);
  or _43340_ (_12141_, _12139_, _12129_);
  and _43341_ (_12143_, _12141_, _05542_);
  or _43342_ (_12144_, _12143_, _12119_);
  and _43343_ (_12145_, _12144_, _05518_);
  or _43344_ (_12146_, _12145_, _12097_);
  and _43345_ (_12147_, _12146_, _05520_);
  or _43346_ (_12149_, _12147_, _12049_);
  or _43347_ (_12150_, _12149_, _05526_);
  and _43348_ (_12151_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and _43349_ (_12152_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _43350_ (_12153_, _12152_, _12151_);
  and _43351_ (_12155_, _12153_, _09792_);
  and _43352_ (_12156_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and _43353_ (_12157_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _43354_ (_12158_, _12157_, _12156_);
  and _43355_ (_12159_, _12158_, _05549_);
  or _43356_ (_12160_, _12159_, _12155_);
  or _43357_ (_12161_, _12160_, _09791_);
  and _43358_ (_12162_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and _43359_ (_12163_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _43360_ (_12164_, _12163_, _12162_);
  and _43361_ (_12165_, _12164_, _09792_);
  and _43362_ (_12166_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and _43363_ (_12167_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _43364_ (_12168_, _12167_, _12166_);
  and _43365_ (_12169_, _12168_, _05549_);
  or _43366_ (_12170_, _12169_, _12165_);
  or _43367_ (_12171_, _12170_, _05535_);
  and _43368_ (_12172_, _12171_, _09805_);
  and _43369_ (_12173_, _12172_, _12161_);
  or _43370_ (_12174_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _43371_ (_12175_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and _43372_ (_12176_, _12175_, _05549_);
  and _43373_ (_12177_, _12176_, _12174_);
  or _43374_ (_12178_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _43375_ (_12179_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and _43376_ (_12180_, _12179_, _09792_);
  and _43377_ (_12181_, _12180_, _12178_);
  or _43378_ (_12182_, _12181_, _12177_);
  or _43379_ (_12183_, _12182_, _09791_);
  or _43380_ (_12184_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _43381_ (_12185_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and _43382_ (_12186_, _12185_, _05549_);
  and _43383_ (_12187_, _12186_, _12184_);
  or _43384_ (_12188_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _43385_ (_12189_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and _43386_ (_12190_, _12189_, _09792_);
  and _43387_ (_12191_, _12190_, _12188_);
  or _43388_ (_12192_, _12191_, _12187_);
  or _43389_ (_12193_, _12192_, _05535_);
  and _43390_ (_12194_, _12193_, _05542_);
  and _43391_ (_12195_, _12194_, _12183_);
  or _43392_ (_12196_, _12195_, _12173_);
  and _43393_ (_12197_, _12196_, _09850_);
  and _43394_ (_12198_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _43395_ (_12199_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _43396_ (_12200_, _12199_, _12198_);
  and _43397_ (_12201_, _12200_, _09792_);
  and _43398_ (_12203_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _43399_ (_12204_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or _43400_ (_12205_, _12204_, _12203_);
  and _43401_ (_12206_, _12205_, _05549_);
  or _43402_ (_12207_, _12206_, _12201_);
  or _43403_ (_12208_, _12207_, _09791_);
  and _43404_ (_12209_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and _43405_ (_12210_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or _43406_ (_12211_, _12210_, _12209_);
  and _43407_ (_12212_, _12211_, _09792_);
  and _43408_ (_12213_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _43409_ (_12214_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _43410_ (_12215_, _12214_, _12213_);
  and _43411_ (_12216_, _12215_, _05549_);
  or _43412_ (_12217_, _12216_, _12212_);
  or _43413_ (_12218_, _12217_, _05535_);
  and _43414_ (_12219_, _12218_, _09805_);
  and _43415_ (_12220_, _12219_, _12208_);
  or _43416_ (_12221_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _43417_ (_12222_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _43418_ (_12223_, _12222_, _12221_);
  and _43419_ (_12225_, _12223_, _09792_);
  or _43420_ (_12226_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _43421_ (_12227_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _43422_ (_12228_, _12227_, _12226_);
  and _43423_ (_12229_, _12228_, _05549_);
  or _43424_ (_12230_, _12229_, _12225_);
  or _43425_ (_12231_, _12230_, _09791_);
  or _43426_ (_12232_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or _43427_ (_12233_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _43428_ (_12234_, _12233_, _12232_);
  and _43429_ (_12235_, _12234_, _09792_);
  or _43430_ (_12236_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _43431_ (_12237_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _43432_ (_12238_, _12237_, _12236_);
  and _43433_ (_12239_, _12238_, _05549_);
  or _43434_ (_12240_, _12239_, _12235_);
  or _43435_ (_12241_, _12240_, _05535_);
  and _43436_ (_12242_, _12241_, _05542_);
  and _43437_ (_12244_, _12242_, _12231_);
  or _43438_ (_12245_, _12244_, _12220_);
  and _43439_ (_12246_, _12245_, _05518_);
  or _43440_ (_12247_, _12246_, _12197_);
  and _43441_ (_12248_, _12247_, _09790_);
  or _43442_ (_12249_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or _43443_ (_12250_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and _43444_ (_12252_, _12250_, _12249_);
  and _43445_ (_12253_, _12252_, _09792_);
  or _43446_ (_12254_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _43447_ (_12255_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _43448_ (_12256_, _12255_, _12254_);
  and _43449_ (_12257_, _12256_, _05549_);
  or _43450_ (_12258_, _12257_, _12253_);
  and _43451_ (_12259_, _12258_, _09791_);
  or _43452_ (_12260_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _43453_ (_12262_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and _43454_ (_12263_, _12262_, _12260_);
  and _43455_ (_12264_, _12263_, _09792_);
  or _43456_ (_12265_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _43457_ (_12267_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _43458_ (_12269_, _12267_, _12265_);
  and _43459_ (_12270_, _12269_, _05549_);
  or _43460_ (_12271_, _12270_, _12264_);
  and _43461_ (_12272_, _12271_, _05535_);
  or _43462_ (_12273_, _12272_, _12259_);
  and _43463_ (_12275_, _12273_, _05542_);
  and _43464_ (_12276_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and _43465_ (_12277_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _43466_ (_12278_, _12277_, _12276_);
  and _43467_ (_12279_, _12278_, _09792_);
  and _43468_ (_12281_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _43469_ (_12282_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _43470_ (_12283_, _12282_, _12281_);
  and _43471_ (_12284_, _12283_, _05549_);
  or _43472_ (_12285_, _12284_, _12279_);
  and _43473_ (_12286_, _12285_, _09791_);
  and _43474_ (_12287_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _43475_ (_12288_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _43476_ (_12289_, _12288_, _12287_);
  and _43477_ (_12290_, _12289_, _09792_);
  and _43478_ (_12291_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _43479_ (_12292_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or _43480_ (_12294_, _12292_, _12291_);
  and _43481_ (_12295_, _12294_, _05549_);
  or _43482_ (_12296_, _12295_, _12290_);
  and _43483_ (_12297_, _12296_, _05535_);
  or _43484_ (_12298_, _12297_, _12286_);
  and _43485_ (_12299_, _12298_, _09805_);
  or _43486_ (_12300_, _12299_, _12275_);
  and _43487_ (_12302_, _12300_, _05518_);
  or _43488_ (_12303_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _43489_ (_12304_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and _43490_ (_12305_, _12304_, _05549_);
  and _43491_ (_12306_, _12305_, _12303_);
  or _43492_ (_12307_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _43493_ (_12308_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and _43494_ (_12309_, _12308_, _09792_);
  and _43495_ (_12310_, _12309_, _12307_);
  or _43496_ (_12311_, _12310_, _12306_);
  and _43497_ (_12312_, _12311_, _09791_);
  or _43498_ (_12313_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _43499_ (_12314_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and _43500_ (_12315_, _12314_, _05549_);
  and _43501_ (_12317_, _12315_, _12313_);
  or _43502_ (_12318_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or _43503_ (_12319_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and _43504_ (_12320_, _12319_, _09792_);
  and _43505_ (_12321_, _12320_, _12318_);
  or _43506_ (_12322_, _12321_, _12317_);
  and _43507_ (_12323_, _12322_, _05535_);
  or _43508_ (_12324_, _12323_, _12312_);
  and _43509_ (_12326_, _12324_, _05542_);
  and _43510_ (_12327_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and _43511_ (_12328_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _43512_ (_12329_, _12328_, _12327_);
  and _43513_ (_12330_, _12329_, _09792_);
  and _43514_ (_12331_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and _43515_ (_12333_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _43516_ (_12335_, _12333_, _12331_);
  and _43517_ (_12336_, _12335_, _05549_);
  or _43518_ (_12337_, _12336_, _12330_);
  and _43519_ (_12338_, _12337_, _09791_);
  and _43520_ (_12339_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and _43521_ (_12341_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _43522_ (_12343_, _12341_, _12339_);
  and _43523_ (_12345_, _12343_, _09792_);
  and _43524_ (_12346_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and _43525_ (_12347_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _43526_ (_12349_, _12347_, _12346_);
  and _43527_ (_12350_, _12349_, _05549_);
  or _43528_ (_12352_, _12350_, _12345_);
  and _43529_ (_12354_, _12352_, _05535_);
  or _43530_ (_12356_, _12354_, _12338_);
  and _43531_ (_12358_, _12356_, _09805_);
  or _43532_ (_12359_, _12358_, _12326_);
  and _43533_ (_12360_, _12359_, _09850_);
  or _43534_ (_12361_, _12360_, _12302_);
  and _43535_ (_12362_, _12361_, _05520_);
  or _43536_ (_12363_, _12362_, _12248_);
  or _43537_ (_12364_, _12363_, _10033_);
  and _43538_ (_12365_, _12364_, _12150_);
  or _43539_ (_12366_, _12365_, _04413_);
  and _43540_ (_12367_, _12366_, _11953_);
  or _43541_ (_12368_, _12367_, _05563_);
  or _43542_ (_12370_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _43543_ (_12371_, _12370_, _22731_);
  and _43544_ (_04460_, _12371_, _12368_);
  and _43545_ (_12372_, _09779_, _23941_);
  and _43546_ (_12373_, _12372_, _23887_);
  not _43547_ (_12374_, _12372_);
  and _43548_ (_12375_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or _43549_ (_04471_, _12375_, _12373_);
  and _43550_ (_12376_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and _43551_ (_12377_, _02513_, _23583_);
  or _43552_ (_04473_, _12377_, _12376_);
  and _43553_ (_12378_, _10746_, _23548_);
  and _43554_ (_12379_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or _43555_ (_04487_, _12379_, _12378_);
  and _43556_ (_12380_, _06763_, _24089_);
  and _43557_ (_12381_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _43558_ (_04490_, _12381_, _12380_);
  and _43559_ (_12382_, _12372_, _23548_);
  and _43560_ (_12383_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or _43561_ (_04492_, _12383_, _12382_);
  and _43562_ (_12385_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and _43563_ (_12386_, _02513_, _24134_);
  or _43564_ (_27089_, _12386_, _12385_);
  and _43565_ (_12388_, _07038_, _23548_);
  and _43566_ (_12389_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _43567_ (_04504_, _12389_, _12388_);
  and _43568_ (_12392_, _07038_, _23583_);
  and _43569_ (_12394_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _43570_ (_04506_, _12394_, _12392_);
  and _43571_ (_12395_, _05438_, _24089_);
  and _43572_ (_12396_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _43573_ (_04509_, _12396_, _12395_);
  and _43574_ (_12398_, _05438_, _24134_);
  and _43575_ (_12400_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _43576_ (_04511_, _12400_, _12398_);
  and _43577_ (_12401_, _07013_, _24051_);
  and _43578_ (_12402_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _43579_ (_04515_, _12402_, _12401_);
  and _43580_ (_12403_, _07038_, _23887_);
  and _43581_ (_12405_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _43582_ (_04525_, _12405_, _12403_);
  and _43583_ (_12406_, _05438_, _24051_);
  and _43584_ (_12407_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _43585_ (_04546_, _12407_, _12406_);
  and _43586_ (_12408_, _24409_, _24089_);
  and _43587_ (_12409_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or _43588_ (_04562_, _12409_, _12408_);
  and _43589_ (_12410_, _12372_, _23583_);
  and _43590_ (_12411_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or _43591_ (_26996_, _12411_, _12410_);
  and _43592_ (_12414_, _12372_, _24051_);
  and _43593_ (_12415_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or _43594_ (_04571_, _12415_, _12414_);
  and _43595_ (_12418_, _12372_, _24089_);
  and _43596_ (_12419_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  or _43597_ (_04576_, _12419_, _12418_);
  and _43598_ (_12421_, _05442_, _24051_);
  and _43599_ (_12423_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _43600_ (_04588_, _12423_, _12421_);
  and _43601_ (_12425_, _05442_, _23996_);
  and _43602_ (_12426_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _43603_ (_04591_, _12426_, _12425_);
  and _43604_ (_12427_, _07013_, _23996_);
  and _43605_ (_12428_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _43606_ (_04600_, _12428_, _12427_);
  and _43607_ (_12429_, _24476_, _23941_);
  and _43608_ (_12430_, _12429_, _23996_);
  not _43609_ (_12431_, _12429_);
  and _43610_ (_12433_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or _43611_ (_04618_, _12433_, _12430_);
  and _43612_ (_12434_, _24510_, _23887_);
  and _43613_ (_12435_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _43614_ (_04621_, _12435_, _12434_);
  and _43615_ (_12436_, _24510_, _23548_);
  and _43616_ (_12437_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _43617_ (_04624_, _12437_, _12436_);
  and _43618_ (_12438_, _24476_, _24297_);
  and _43619_ (_12439_, _12438_, _23887_);
  not _43620_ (_12440_, _12438_);
  and _43621_ (_12441_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or _43622_ (_04655_, _12441_, _12439_);
  and _43623_ (_12442_, _09779_, _24899_);
  and _43624_ (_12443_, _12442_, _24089_);
  not _43625_ (_12444_, _12442_);
  and _43626_ (_12445_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or _43627_ (_04664_, _12445_, _12443_);
  and _43628_ (_12446_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _43629_ (_12447_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _43630_ (_12448_, _12447_, _12446_);
  and _43631_ (_12449_, _12448_, _09792_);
  and _43632_ (_12450_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and _43633_ (_12451_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _43634_ (_12452_, _12451_, _12450_);
  and _43635_ (_12453_, _12452_, _05549_);
  or _43636_ (_12454_, _12453_, _12449_);
  or _43637_ (_12455_, _12454_, _09791_);
  and _43638_ (_12456_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and _43639_ (_12457_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _43640_ (_12458_, _12457_, _12456_);
  and _43641_ (_12459_, _12458_, _09792_);
  and _43642_ (_12460_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and _43643_ (_12461_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _43644_ (_12462_, _12461_, _12460_);
  and _43645_ (_12463_, _12462_, _05549_);
  or _43646_ (_12464_, _12463_, _12459_);
  or _43647_ (_12465_, _12464_, _05535_);
  and _43648_ (_12466_, _12465_, _09805_);
  and _43649_ (_12467_, _12466_, _12455_);
  or _43650_ (_12468_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _43651_ (_12469_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and _43652_ (_12470_, _12469_, _12468_);
  and _43653_ (_12471_, _12470_, _09792_);
  or _43654_ (_12472_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _43655_ (_12473_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and _43656_ (_12474_, _12473_, _12472_);
  and _43657_ (_12475_, _12474_, _05549_);
  or _43658_ (_12476_, _12475_, _12471_);
  or _43659_ (_12477_, _12476_, _09791_);
  or _43660_ (_12478_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _43661_ (_12479_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and _43662_ (_12480_, _12479_, _12478_);
  and _43663_ (_12481_, _12480_, _09792_);
  or _43664_ (_12482_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _43665_ (_12483_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and _43666_ (_12484_, _12483_, _12482_);
  and _43667_ (_12485_, _12484_, _05549_);
  or _43668_ (_12486_, _12485_, _12481_);
  or _43669_ (_12487_, _12486_, _05535_);
  and _43670_ (_12488_, _12487_, _05542_);
  and _43671_ (_12489_, _12488_, _12477_);
  or _43672_ (_12490_, _12489_, _12467_);
  and _43673_ (_12491_, _12490_, _05518_);
  and _43674_ (_12492_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and _43675_ (_12493_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _43676_ (_12494_, _12493_, _12492_);
  and _43677_ (_12495_, _12494_, _09792_);
  and _43678_ (_12496_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and _43679_ (_12497_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _43680_ (_12498_, _12497_, _12496_);
  and _43681_ (_12499_, _12498_, _05549_);
  or _43682_ (_12500_, _12499_, _12495_);
  or _43683_ (_12501_, _12500_, _09791_);
  and _43684_ (_12502_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and _43685_ (_12503_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _43686_ (_12504_, _12503_, _12502_);
  and _43687_ (_12505_, _12504_, _09792_);
  and _43688_ (_12506_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and _43689_ (_12507_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _43690_ (_12508_, _12507_, _12506_);
  and _43691_ (_12509_, _12508_, _05549_);
  or _43692_ (_12510_, _12509_, _12505_);
  or _43693_ (_12511_, _12510_, _05535_);
  and _43694_ (_12512_, _12511_, _09805_);
  and _43695_ (_12513_, _12512_, _12501_);
  or _43696_ (_12514_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _43697_ (_12516_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and _43698_ (_12517_, _12516_, _05549_);
  and _43699_ (_12518_, _12517_, _12514_);
  or _43700_ (_12519_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _43701_ (_12520_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and _43702_ (_12521_, _12520_, _09792_);
  and _43703_ (_12522_, _12521_, _12519_);
  or _43704_ (_12523_, _12522_, _12518_);
  or _43705_ (_12524_, _12523_, _09791_);
  or _43706_ (_12525_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _43707_ (_12526_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and _43708_ (_12527_, _12526_, _05549_);
  and _43709_ (_12528_, _12527_, _12525_);
  or _43710_ (_12529_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _43711_ (_12530_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and _43712_ (_12531_, _12530_, _09792_);
  and _43713_ (_12532_, _12531_, _12529_);
  or _43714_ (_12533_, _12532_, _12528_);
  or _43715_ (_12534_, _12533_, _05535_);
  and _43716_ (_12535_, _12534_, _05542_);
  and _43717_ (_12536_, _12535_, _12524_);
  or _43718_ (_12537_, _12536_, _12513_);
  and _43719_ (_12538_, _12537_, _09850_);
  or _43720_ (_12539_, _12538_, _12491_);
  and _43721_ (_12540_, _12539_, _09790_);
  and _43722_ (_12541_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _43723_ (_12542_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or _43724_ (_12543_, _12542_, _12541_);
  and _43725_ (_12544_, _12543_, _09792_);
  and _43726_ (_12545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and _43727_ (_12546_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _43728_ (_12547_, _12546_, _12545_);
  and _43729_ (_12548_, _12547_, _05549_);
  or _43730_ (_12549_, _12548_, _12544_);
  and _43731_ (_12550_, _12549_, _05535_);
  and _43732_ (_12551_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _43733_ (_12552_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _43734_ (_12553_, _12552_, _12551_);
  and _43735_ (_12554_, _12553_, _09792_);
  and _43736_ (_12555_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and _43737_ (_12556_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _43738_ (_12557_, _12556_, _12555_);
  and _43739_ (_12558_, _12557_, _05549_);
  or _43740_ (_12559_, _12558_, _12554_);
  and _43741_ (_12560_, _12559_, _09791_);
  or _43742_ (_12561_, _12560_, _12550_);
  and _43743_ (_12562_, _12561_, _09805_);
  or _43744_ (_12563_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _43745_ (_12564_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and _43746_ (_12565_, _12564_, _05549_);
  and _43747_ (_12566_, _12565_, _12563_);
  or _43748_ (_12567_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _43749_ (_12568_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and _43750_ (_12569_, _12568_, _09792_);
  and _43751_ (_12570_, _12569_, _12567_);
  or _43752_ (_12571_, _12570_, _12566_);
  and _43753_ (_12572_, _12571_, _05535_);
  or _43754_ (_12573_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _43755_ (_12574_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _43756_ (_12575_, _12574_, _05549_);
  and _43757_ (_12576_, _12575_, _12573_);
  or _43758_ (_12577_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _43759_ (_12578_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and _43760_ (_12579_, _12578_, _09792_);
  and _43761_ (_12580_, _12579_, _12577_);
  or _43762_ (_12581_, _12580_, _12576_);
  and _43763_ (_12582_, _12581_, _09791_);
  or _43764_ (_12583_, _12582_, _12572_);
  and _43765_ (_12584_, _12583_, _05542_);
  or _43766_ (_12585_, _12584_, _12562_);
  and _43767_ (_12586_, _12585_, _09850_);
  and _43768_ (_12587_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and _43769_ (_12588_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _43770_ (_12589_, _12588_, _12587_);
  and _43771_ (_12590_, _12589_, _09792_);
  and _43772_ (_12591_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and _43773_ (_12592_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _43774_ (_12593_, _12592_, _12591_);
  and _43775_ (_12594_, _12593_, _05549_);
  or _43776_ (_12595_, _12594_, _12590_);
  and _43777_ (_12596_, _12595_, _05535_);
  and _43778_ (_12597_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and _43779_ (_12598_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _43780_ (_12599_, _12598_, _12597_);
  and _43781_ (_12600_, _12599_, _09792_);
  and _43782_ (_12601_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and _43783_ (_12602_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _43784_ (_12603_, _12602_, _12601_);
  and _43785_ (_12604_, _12603_, _05549_);
  or _43786_ (_12605_, _12604_, _12600_);
  and _43787_ (_12606_, _12605_, _09791_);
  or _43788_ (_12607_, _12606_, _12596_);
  and _43789_ (_12608_, _12607_, _09805_);
  or _43790_ (_12609_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _43791_ (_12610_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and _43792_ (_12611_, _12610_, _12609_);
  and _43793_ (_12612_, _12611_, _09792_);
  or _43794_ (_12613_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _43795_ (_12614_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and _43796_ (_12615_, _12614_, _12613_);
  and _43797_ (_12617_, _12615_, _05549_);
  or _43798_ (_12618_, _12617_, _12612_);
  and _43799_ (_12619_, _12618_, _05535_);
  or _43800_ (_12620_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _43801_ (_12621_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and _43802_ (_12622_, _12621_, _12620_);
  and _43803_ (_12623_, _12622_, _09792_);
  or _43804_ (_12624_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _43805_ (_12625_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and _43806_ (_12626_, _12625_, _12624_);
  and _43807_ (_12627_, _12626_, _05549_);
  or _43808_ (_12628_, _12627_, _12623_);
  and _43809_ (_12629_, _12628_, _09791_);
  or _43810_ (_12630_, _12629_, _12619_);
  and _43811_ (_12631_, _12630_, _05542_);
  or _43812_ (_12632_, _12631_, _12608_);
  and _43813_ (_12633_, _12632_, _05518_);
  or _43814_ (_12634_, _12633_, _12586_);
  and _43815_ (_12635_, _12634_, _05520_);
  or _43816_ (_12636_, _12635_, _12540_);
  or _43817_ (_12638_, _12636_, _05526_);
  and _43818_ (_12639_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and _43819_ (_12640_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _43820_ (_12641_, _12640_, _12639_);
  and _43821_ (_12642_, _12641_, _09792_);
  and _43822_ (_12643_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and _43823_ (_12644_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _43824_ (_12645_, _12644_, _12643_);
  and _43825_ (_12646_, _12645_, _05549_);
  or _43826_ (_12647_, _12646_, _12642_);
  or _43827_ (_12648_, _12647_, _09791_);
  and _43828_ (_12649_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and _43829_ (_12650_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _43830_ (_12651_, _12650_, _12649_);
  and _43831_ (_12652_, _12651_, _09792_);
  and _43832_ (_12653_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and _43833_ (_12654_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _43834_ (_12655_, _12654_, _12653_);
  and _43835_ (_12656_, _12655_, _05549_);
  or _43836_ (_12657_, _12656_, _12652_);
  or _43837_ (_12658_, _12657_, _05535_);
  and _43838_ (_12659_, _12658_, _09805_);
  and _43839_ (_12660_, _12659_, _12648_);
  or _43840_ (_12661_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _43841_ (_12662_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and _43842_ (_12663_, _12662_, _05549_);
  and _43843_ (_12664_, _12663_, _12661_);
  or _43844_ (_12665_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _43845_ (_12666_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and _43846_ (_12667_, _12666_, _09792_);
  and _43847_ (_12668_, _12667_, _12665_);
  or _43848_ (_12669_, _12668_, _12664_);
  or _43849_ (_12670_, _12669_, _09791_);
  or _43850_ (_12671_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _43851_ (_12672_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and _43852_ (_12673_, _12672_, _05549_);
  and _43853_ (_12674_, _12673_, _12671_);
  or _43854_ (_12675_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _43855_ (_12676_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and _43856_ (_12677_, _12676_, _09792_);
  and _43857_ (_12678_, _12677_, _12675_);
  or _43858_ (_12679_, _12678_, _12674_);
  or _43859_ (_12680_, _12679_, _05535_);
  and _43860_ (_12681_, _12680_, _05542_);
  and _43861_ (_12682_, _12681_, _12670_);
  or _43862_ (_12683_, _12682_, _12660_);
  and _43863_ (_12684_, _12683_, _09850_);
  and _43864_ (_12685_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and _43865_ (_12686_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _43866_ (_12687_, _12686_, _12685_);
  and _43867_ (_12688_, _12687_, _09792_);
  and _43868_ (_12689_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and _43869_ (_12690_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _43870_ (_12691_, _12690_, _12689_);
  and _43871_ (_12692_, _12691_, _05549_);
  or _43872_ (_12693_, _12692_, _12688_);
  or _43873_ (_12694_, _12693_, _09791_);
  and _43874_ (_12695_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and _43875_ (_12696_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _43876_ (_12697_, _12696_, _12695_);
  and _43877_ (_12698_, _12697_, _09792_);
  and _43878_ (_12699_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and _43879_ (_12700_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _43880_ (_12701_, _12700_, _12699_);
  and _43881_ (_12702_, _12701_, _05549_);
  or _43882_ (_12703_, _12702_, _12698_);
  or _43883_ (_12704_, _12703_, _05535_);
  and _43884_ (_12705_, _12704_, _09805_);
  and _43885_ (_12706_, _12705_, _12694_);
  or _43886_ (_12707_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _43887_ (_12708_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and _43888_ (_12709_, _12708_, _12707_);
  and _43889_ (_12710_, _12709_, _09792_);
  or _43890_ (_12711_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _43891_ (_12712_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and _43892_ (_12713_, _12712_, _12711_);
  and _43893_ (_12714_, _12713_, _05549_);
  or _43894_ (_12715_, _12714_, _12710_);
  or _43895_ (_12716_, _12715_, _09791_);
  or _43896_ (_12717_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _43897_ (_12718_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and _43898_ (_12719_, _12718_, _12717_);
  and _43899_ (_12720_, _12719_, _09792_);
  or _43900_ (_12721_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _43901_ (_12722_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and _43902_ (_12723_, _12722_, _12721_);
  and _43903_ (_12724_, _12723_, _05549_);
  or _43904_ (_12725_, _12724_, _12720_);
  or _43905_ (_12726_, _12725_, _05535_);
  and _43906_ (_12727_, _12726_, _05542_);
  and _43907_ (_12728_, _12727_, _12716_);
  or _43908_ (_12729_, _12728_, _12706_);
  and _43909_ (_12730_, _12729_, _05518_);
  or _43910_ (_12731_, _12730_, _12684_);
  and _43911_ (_12732_, _12731_, _09790_);
  or _43912_ (_12733_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _43913_ (_12734_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and _43914_ (_12735_, _12734_, _12733_);
  and _43915_ (_12736_, _12735_, _09792_);
  or _43916_ (_12737_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _43917_ (_12738_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and _43918_ (_12739_, _12738_, _12737_);
  and _43919_ (_12740_, _12739_, _05549_);
  or _43920_ (_12741_, _12740_, _12736_);
  and _43921_ (_12742_, _12741_, _09791_);
  or _43922_ (_12743_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _43923_ (_12744_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and _43924_ (_12745_, _12744_, _12743_);
  and _43925_ (_12746_, _12745_, _09792_);
  or _43926_ (_12747_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _43927_ (_12749_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and _43928_ (_12750_, _12749_, _12747_);
  and _43929_ (_12751_, _12750_, _05549_);
  or _43930_ (_12752_, _12751_, _12746_);
  and _43931_ (_12753_, _12752_, _05535_);
  or _43932_ (_12754_, _12753_, _12742_);
  and _43933_ (_12755_, _12754_, _05542_);
  and _43934_ (_12756_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and _43935_ (_12757_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _43936_ (_12758_, _12757_, _12756_);
  and _43937_ (_12759_, _12758_, _09792_);
  and _43938_ (_12760_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and _43939_ (_12761_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _43940_ (_12762_, _12761_, _12760_);
  and _43941_ (_12763_, _12762_, _05549_);
  or _43942_ (_12764_, _12763_, _12759_);
  and _43943_ (_12765_, _12764_, _09791_);
  and _43944_ (_12766_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and _43945_ (_12767_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _43946_ (_12768_, _12767_, _12766_);
  and _43947_ (_12769_, _12768_, _09792_);
  and _43948_ (_12770_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and _43949_ (_12771_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _43950_ (_12772_, _12771_, _12770_);
  and _43951_ (_12773_, _12772_, _05549_);
  or _43952_ (_12774_, _12773_, _12769_);
  and _43953_ (_12775_, _12774_, _05535_);
  or _43954_ (_12776_, _12775_, _12765_);
  and _43955_ (_12777_, _12776_, _09805_);
  or _43956_ (_12778_, _12777_, _12755_);
  and _43957_ (_12779_, _12778_, _05518_);
  or _43958_ (_12780_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or _43959_ (_12781_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and _43960_ (_12782_, _12781_, _05549_);
  and _43961_ (_12783_, _12782_, _12780_);
  or _43962_ (_12784_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or _43963_ (_12785_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and _43964_ (_12786_, _12785_, _09792_);
  and _43965_ (_12787_, _12786_, _12784_);
  or _43966_ (_12788_, _12787_, _12783_);
  and _43967_ (_12789_, _12788_, _09791_);
  or _43968_ (_12790_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or _43969_ (_12791_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and _43970_ (_12792_, _12791_, _05549_);
  and _43971_ (_12793_, _12792_, _12790_);
  or _43972_ (_12794_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or _43973_ (_12795_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and _43974_ (_12796_, _12795_, _09792_);
  and _43975_ (_12797_, _12796_, _12794_);
  or _43976_ (_12798_, _12797_, _12793_);
  and _43977_ (_12799_, _12798_, _05535_);
  or _43978_ (_12800_, _12799_, _12789_);
  and _43979_ (_12801_, _12800_, _05542_);
  and _43980_ (_12802_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and _43981_ (_12803_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or _43982_ (_12804_, _12803_, _12802_);
  and _43983_ (_12805_, _12804_, _09792_);
  and _43984_ (_12806_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and _43985_ (_12807_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or _43986_ (_12808_, _12807_, _12806_);
  and _43987_ (_12809_, _12808_, _05549_);
  or _43988_ (_12810_, _12809_, _12805_);
  and _43989_ (_12811_, _12810_, _09791_);
  and _43990_ (_12812_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and _43991_ (_12813_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or _43992_ (_12814_, _12813_, _12812_);
  and _43993_ (_12815_, _12814_, _09792_);
  and _43994_ (_12816_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and _43995_ (_12817_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or _43996_ (_12818_, _12817_, _12816_);
  and _43997_ (_12819_, _12818_, _05549_);
  or _43998_ (_12820_, _12819_, _12815_);
  and _43999_ (_12821_, _12820_, _05535_);
  or _44000_ (_12822_, _12821_, _12811_);
  and _44001_ (_12823_, _12822_, _09805_);
  or _44002_ (_12824_, _12823_, _12801_);
  and _44003_ (_12825_, _12824_, _09850_);
  or _44004_ (_12826_, _12825_, _12779_);
  and _44005_ (_12827_, _12826_, _05520_);
  or _44006_ (_12828_, _12827_, _12732_);
  or _44007_ (_12829_, _12828_, _10033_);
  and _44008_ (_12830_, _12829_, _12638_);
  or _44009_ (_12831_, _12830_, _00143_);
  and _44010_ (_12832_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and _44011_ (_12833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _44012_ (_12834_, _12833_, _12832_);
  and _44013_ (_12835_, _12834_, _09792_);
  and _44014_ (_12836_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and _44015_ (_12837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _44016_ (_12838_, _12837_, _12836_);
  and _44017_ (_12839_, _12838_, _05549_);
  or _44018_ (_12840_, _12839_, _12835_);
  or _44019_ (_12841_, _12840_, _09791_);
  and _44020_ (_12842_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and _44021_ (_12843_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _44022_ (_12844_, _12843_, _12842_);
  and _44023_ (_12845_, _12844_, _09792_);
  and _44024_ (_12846_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and _44025_ (_12847_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _44026_ (_12848_, _12847_, _12846_);
  and _44027_ (_12849_, _12848_, _05549_);
  or _44028_ (_12850_, _12849_, _12845_);
  or _44029_ (_12851_, _12850_, _05535_);
  and _44030_ (_12852_, _12851_, _09805_);
  and _44031_ (_12853_, _12852_, _12841_);
  or _44032_ (_12854_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _44033_ (_12855_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and _44034_ (_12856_, _12855_, _12854_);
  and _44035_ (_12857_, _12856_, _09792_);
  or _44036_ (_12858_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _44037_ (_12859_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and _44038_ (_12860_, _12859_, _12858_);
  and _44039_ (_12861_, _12860_, _05549_);
  or _44040_ (_12862_, _12861_, _12857_);
  or _44041_ (_12863_, _12862_, _09791_);
  or _44042_ (_12864_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _44043_ (_12865_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and _44044_ (_12866_, _12865_, _12864_);
  and _44045_ (_12867_, _12866_, _09792_);
  or _44046_ (_12868_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _44047_ (_12869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and _44048_ (_12870_, _12869_, _12868_);
  and _44049_ (_12871_, _12870_, _05549_);
  or _44050_ (_12872_, _12871_, _12867_);
  or _44051_ (_12873_, _12872_, _05535_);
  and _44052_ (_12874_, _12873_, _05542_);
  and _44053_ (_12875_, _12874_, _12863_);
  or _44054_ (_12876_, _12875_, _12853_);
  and _44055_ (_12877_, _12876_, _05518_);
  and _44056_ (_12878_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and _44057_ (_12879_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or _44058_ (_12880_, _12879_, _12878_);
  and _44059_ (_12881_, _12880_, _09792_);
  and _44060_ (_12882_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _44061_ (_12883_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or _44062_ (_12884_, _12883_, _12882_);
  and _44063_ (_12885_, _12884_, _05549_);
  or _44064_ (_12886_, _12885_, _12881_);
  or _44065_ (_12887_, _12886_, _09791_);
  and _44066_ (_12888_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _44067_ (_12889_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _44068_ (_12890_, _12889_, _12888_);
  and _44069_ (_12891_, _12890_, _09792_);
  and _44070_ (_12892_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _44071_ (_12893_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _44072_ (_12894_, _12893_, _12892_);
  and _44073_ (_12895_, _12894_, _05549_);
  or _44074_ (_12896_, _12895_, _12891_);
  or _44075_ (_12897_, _12896_, _05535_);
  and _44076_ (_12898_, _12897_, _09805_);
  and _44077_ (_12899_, _12898_, _12887_);
  or _44078_ (_12900_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or _44079_ (_12901_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _44080_ (_12902_, _12901_, _05549_);
  and _44081_ (_12903_, _12902_, _12900_);
  or _44082_ (_12904_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _44083_ (_12905_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _44084_ (_12906_, _12905_, _09792_);
  and _44085_ (_12907_, _12906_, _12904_);
  or _44086_ (_12908_, _12907_, _12903_);
  or _44087_ (_12909_, _12908_, _09791_);
  or _44088_ (_12910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or _44089_ (_12911_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and _44090_ (_12912_, _12911_, _05549_);
  and _44091_ (_12913_, _12912_, _12910_);
  or _44092_ (_12914_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _44093_ (_12915_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _44094_ (_12916_, _12915_, _09792_);
  and _44095_ (_12917_, _12916_, _12914_);
  or _44096_ (_12918_, _12917_, _12913_);
  or _44097_ (_12919_, _12918_, _05535_);
  and _44098_ (_12920_, _12919_, _05542_);
  and _44099_ (_12921_, _12920_, _12909_);
  or _44100_ (_12922_, _12921_, _12899_);
  and _44101_ (_12923_, _12922_, _09850_);
  or _44102_ (_12924_, _12923_, _12877_);
  and _44103_ (_12925_, _12924_, _09790_);
  and _44104_ (_12926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and _44105_ (_12927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or _44106_ (_12928_, _12927_, _12926_);
  and _44107_ (_12929_, _12928_, _09792_);
  and _44108_ (_12930_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _44109_ (_12931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or _44110_ (_12932_, _12931_, _12930_);
  and _44111_ (_12933_, _12932_, _05549_);
  or _44112_ (_12934_, _12933_, _12929_);
  and _44113_ (_12935_, _12934_, _05535_);
  and _44114_ (_12936_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and _44115_ (_12937_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or _44116_ (_12938_, _12937_, _12936_);
  and _44117_ (_12939_, _12938_, _09792_);
  and _44118_ (_12940_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and _44119_ (_12941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or _44120_ (_12942_, _12941_, _12940_);
  and _44121_ (_12943_, _12942_, _05549_);
  or _44122_ (_12944_, _12943_, _12939_);
  and _44123_ (_12945_, _12944_, _09791_);
  or _44124_ (_12946_, _12945_, _12935_);
  and _44125_ (_12947_, _12946_, _09805_);
  or _44126_ (_12948_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or _44127_ (_12949_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and _44128_ (_12950_, _12949_, _05549_);
  and _44129_ (_12951_, _12950_, _12948_);
  or _44130_ (_12952_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or _44131_ (_12953_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and _44132_ (_12954_, _12953_, _09792_);
  and _44133_ (_12955_, _12954_, _12952_);
  or _44134_ (_12956_, _12955_, _12951_);
  and _44135_ (_12957_, _12956_, _05535_);
  or _44136_ (_12958_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or _44137_ (_12959_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and _44138_ (_12960_, _12959_, _05549_);
  and _44139_ (_12961_, _12960_, _12958_);
  or _44140_ (_12962_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or _44141_ (_12963_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and _44142_ (_12964_, _12963_, _09792_);
  and _44143_ (_12965_, _12964_, _12962_);
  or _44144_ (_12966_, _12965_, _12961_);
  and _44145_ (_12967_, _12966_, _09791_);
  or _44146_ (_12968_, _12967_, _12957_);
  and _44147_ (_12969_, _12968_, _05542_);
  or _44148_ (_12970_, _12969_, _12947_);
  and _44149_ (_12971_, _12970_, _09850_);
  and _44150_ (_12972_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _44151_ (_12973_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _44152_ (_12974_, _12973_, _12972_);
  and _44153_ (_12975_, _12974_, _09792_);
  and _44154_ (_12976_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and _44155_ (_12977_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _44156_ (_12978_, _12977_, _12976_);
  and _44157_ (_12979_, _12978_, _05549_);
  or _44158_ (_12980_, _12979_, _12975_);
  and _44159_ (_12981_, _12980_, _05535_);
  and _44160_ (_12982_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and _44161_ (_12983_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _44162_ (_12984_, _12983_, _12982_);
  and _44163_ (_12985_, _12984_, _09792_);
  and _44164_ (_12986_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and _44165_ (_12987_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _44166_ (_12988_, _12987_, _12986_);
  and _44167_ (_12989_, _12988_, _05549_);
  or _44168_ (_12990_, _12989_, _12985_);
  and _44169_ (_12991_, _12990_, _09791_);
  or _44170_ (_12992_, _12991_, _12981_);
  and _44171_ (_12993_, _12992_, _09805_);
  or _44172_ (_12994_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _44173_ (_12995_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and _44174_ (_12996_, _12995_, _12994_);
  and _44175_ (_12997_, _12996_, _09792_);
  or _44176_ (_12998_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _44177_ (_12999_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and _44178_ (_13000_, _12999_, _12998_);
  and _44179_ (_13001_, _13000_, _05549_);
  or _44180_ (_13002_, _13001_, _12997_);
  and _44181_ (_13003_, _13002_, _05535_);
  or _44182_ (_13004_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _44183_ (_13005_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _44184_ (_13006_, _13005_, _13004_);
  and _44185_ (_13007_, _13006_, _09792_);
  or _44186_ (_13008_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _44187_ (_13009_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and _44188_ (_13010_, _13009_, _13008_);
  and _44189_ (_13011_, _13010_, _05549_);
  or _44190_ (_13012_, _13011_, _13007_);
  and _44191_ (_13013_, _13012_, _09791_);
  or _44192_ (_13014_, _13013_, _13003_);
  and _44193_ (_13015_, _13014_, _05542_);
  or _44194_ (_13016_, _13015_, _12993_);
  and _44195_ (_13017_, _13016_, _05518_);
  or _44196_ (_13018_, _13017_, _12971_);
  and _44197_ (_13019_, _13018_, _05520_);
  or _44198_ (_13020_, _13019_, _12925_);
  or _44199_ (_13021_, _13020_, _05526_);
  and _44200_ (_13022_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and _44201_ (_13023_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _44202_ (_13024_, _13023_, _13022_);
  and _44203_ (_13025_, _13024_, _09792_);
  and _44204_ (_13026_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and _44205_ (_13027_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _44206_ (_13028_, _13027_, _13026_);
  and _44207_ (_13029_, _13028_, _05549_);
  or _44208_ (_13030_, _13029_, _13025_);
  or _44209_ (_13031_, _13030_, _09791_);
  and _44210_ (_13032_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and _44211_ (_13033_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _44212_ (_13034_, _13033_, _13032_);
  and _44213_ (_13035_, _13034_, _09792_);
  and _44214_ (_13036_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and _44215_ (_13037_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _44216_ (_13038_, _13037_, _13036_);
  and _44217_ (_13039_, _13038_, _05549_);
  or _44218_ (_13040_, _13039_, _13035_);
  or _44219_ (_13041_, _13040_, _05535_);
  and _44220_ (_13042_, _13041_, _09805_);
  and _44221_ (_13043_, _13042_, _13031_);
  or _44222_ (_13044_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _44223_ (_13045_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and _44224_ (_13046_, _13045_, _05549_);
  and _44225_ (_13047_, _13046_, _13044_);
  or _44226_ (_13048_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _44227_ (_13049_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and _44228_ (_13050_, _13049_, _09792_);
  and _44229_ (_13051_, _13050_, _13048_);
  or _44230_ (_13052_, _13051_, _13047_);
  or _44231_ (_13053_, _13052_, _09791_);
  or _44232_ (_13054_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _44233_ (_13055_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and _44234_ (_13056_, _13055_, _05549_);
  and _44235_ (_13057_, _13056_, _13054_);
  or _44236_ (_13058_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _44237_ (_13059_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and _44238_ (_13060_, _13059_, _09792_);
  and _44239_ (_13061_, _13060_, _13058_);
  or _44240_ (_13062_, _13061_, _13057_);
  or _44241_ (_13063_, _13062_, _05535_);
  and _44242_ (_13064_, _13063_, _05542_);
  and _44243_ (_13065_, _13064_, _13053_);
  or _44244_ (_13066_, _13065_, _13043_);
  and _44245_ (_13067_, _13066_, _09850_);
  and _44246_ (_13068_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and _44247_ (_13069_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or _44248_ (_13070_, _13069_, _13068_);
  and _44249_ (_13071_, _13070_, _09792_);
  and _44250_ (_13072_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _44251_ (_13073_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _44252_ (_13074_, _13073_, _13072_);
  and _44253_ (_13075_, _13074_, _05549_);
  or _44254_ (_13076_, _13075_, _13071_);
  or _44255_ (_13077_, _13076_, _09791_);
  and _44256_ (_13078_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _44257_ (_13079_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or _44258_ (_13080_, _13079_, _13078_);
  and _44259_ (_13081_, _13080_, _09792_);
  and _44260_ (_13082_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _44261_ (_13083_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _44262_ (_13084_, _13083_, _13082_);
  and _44263_ (_13085_, _13084_, _05549_);
  or _44264_ (_13086_, _13085_, _13081_);
  or _44265_ (_13087_, _13086_, _05535_);
  and _44266_ (_13088_, _13087_, _09805_);
  and _44267_ (_13089_, _13088_, _13077_);
  or _44268_ (_13090_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _44269_ (_13091_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _44270_ (_13092_, _13091_, _13090_);
  and _44271_ (_13093_, _13092_, _09792_);
  or _44272_ (_13094_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _44273_ (_13095_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and _44274_ (_13096_, _13095_, _13094_);
  and _44275_ (_13097_, _13096_, _05549_);
  or _44276_ (_13098_, _13097_, _13093_);
  or _44277_ (_13099_, _13098_, _09791_);
  or _44278_ (_13100_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or _44279_ (_13101_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _44280_ (_13102_, _13101_, _13100_);
  and _44281_ (_13103_, _13102_, _09792_);
  or _44282_ (_13104_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _44283_ (_13105_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _44284_ (_13106_, _13105_, _13104_);
  and _44285_ (_13107_, _13106_, _05549_);
  or _44286_ (_13108_, _13107_, _13103_);
  or _44287_ (_13110_, _13108_, _05535_);
  and _44288_ (_13111_, _13110_, _05542_);
  and _44289_ (_13112_, _13111_, _13099_);
  or _44290_ (_13113_, _13112_, _13089_);
  and _44291_ (_13114_, _13113_, _05518_);
  or _44292_ (_13115_, _13114_, _13067_);
  and _44293_ (_13116_, _13115_, _09790_);
  or _44294_ (_13117_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _44295_ (_13118_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and _44296_ (_13119_, _13118_, _13117_);
  and _44297_ (_13120_, _13119_, _09792_);
  or _44298_ (_13121_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _44299_ (_13122_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _44300_ (_13123_, _13122_, _13121_);
  and _44301_ (_13124_, _13123_, _05549_);
  or _44302_ (_13125_, _13124_, _13120_);
  and _44303_ (_13126_, _13125_, _09791_);
  or _44304_ (_13127_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _44305_ (_13128_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _44306_ (_13129_, _13128_, _13127_);
  and _44307_ (_13130_, _13129_, _09792_);
  or _44308_ (_13131_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or _44309_ (_13132_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _44310_ (_13133_, _13132_, _13131_);
  and _44311_ (_13134_, _13133_, _05549_);
  or _44312_ (_13135_, _13134_, _13130_);
  and _44313_ (_13136_, _13135_, _05535_);
  or _44314_ (_13137_, _13136_, _13126_);
  and _44315_ (_13138_, _13137_, _05542_);
  and _44316_ (_13139_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _44317_ (_13140_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or _44318_ (_13141_, _13140_, _13139_);
  and _44319_ (_13142_, _13141_, _09792_);
  and _44320_ (_13143_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _44321_ (_13144_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _44322_ (_13145_, _13144_, _13143_);
  and _44323_ (_13146_, _13145_, _05549_);
  or _44324_ (_13147_, _13146_, _13142_);
  and _44325_ (_13148_, _13147_, _09791_);
  and _44326_ (_13149_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _44327_ (_13150_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _44328_ (_13151_, _13150_, _13149_);
  and _44329_ (_13152_, _13151_, _09792_);
  and _44330_ (_13153_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _44331_ (_13154_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or _44332_ (_13155_, _13154_, _13153_);
  and _44333_ (_13156_, _13155_, _05549_);
  or _44334_ (_13157_, _13156_, _13152_);
  and _44335_ (_13158_, _13157_, _05535_);
  or _44336_ (_13159_, _13158_, _13148_);
  and _44337_ (_13160_, _13159_, _09805_);
  or _44338_ (_13161_, _13160_, _13138_);
  and _44339_ (_13162_, _13161_, _05518_);
  or _44340_ (_13163_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _44341_ (_13164_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and _44342_ (_13165_, _13164_, _05549_);
  and _44343_ (_13166_, _13165_, _13163_);
  or _44344_ (_13167_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _44345_ (_13168_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and _44346_ (_13169_, _13168_, _09792_);
  and _44347_ (_13170_, _13169_, _13167_);
  or _44348_ (_13171_, _13170_, _13166_);
  and _44349_ (_13172_, _13171_, _09791_);
  or _44350_ (_13173_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _44351_ (_13174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and _44352_ (_13175_, _13174_, _05549_);
  and _44353_ (_13176_, _13175_, _13173_);
  or _44354_ (_13177_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _44355_ (_13178_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and _44356_ (_13179_, _13178_, _09792_);
  and _44357_ (_13180_, _13179_, _13177_);
  or _44358_ (_13181_, _13180_, _13176_);
  and _44359_ (_13182_, _13181_, _05535_);
  or _44360_ (_13183_, _13182_, _13172_);
  and _44361_ (_13184_, _13183_, _05542_);
  and _44362_ (_13185_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and _44363_ (_13186_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _44364_ (_13187_, _13186_, _13185_);
  and _44365_ (_13188_, _13187_, _09792_);
  and _44366_ (_13189_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and _44367_ (_13190_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _44368_ (_13191_, _13190_, _13189_);
  and _44369_ (_13192_, _13191_, _05549_);
  or _44370_ (_13193_, _13192_, _13188_);
  and _44371_ (_13194_, _13193_, _09791_);
  and _44372_ (_13195_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and _44373_ (_13196_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _44374_ (_13197_, _13196_, _13195_);
  and _44375_ (_13198_, _13197_, _09792_);
  and _44376_ (_13199_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _44377_ (_13200_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _44378_ (_13201_, _13200_, _13199_);
  and _44379_ (_13202_, _13201_, _05549_);
  or _44380_ (_13203_, _13202_, _13198_);
  and _44381_ (_13204_, _13203_, _05535_);
  or _44382_ (_13205_, _13204_, _13194_);
  and _44383_ (_13206_, _13205_, _09805_);
  or _44384_ (_13207_, _13206_, _13184_);
  and _44385_ (_13208_, _13207_, _09850_);
  or _44386_ (_13209_, _13208_, _13162_);
  and _44387_ (_13210_, _13209_, _05520_);
  or _44388_ (_13211_, _13210_, _13116_);
  or _44389_ (_13212_, _13211_, _10033_);
  and _44390_ (_13213_, _13212_, _13021_);
  or _44391_ (_13214_, _13213_, _04413_);
  and _44392_ (_13215_, _13214_, _12831_);
  or _44393_ (_13216_, _13215_, _05563_);
  or _44394_ (_13217_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _44395_ (_13218_, _13217_, _22731_);
  and _44396_ (_04666_, _13218_, _13216_);
  and _44397_ (_13219_, _12438_, _23548_);
  and _44398_ (_13220_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or _44399_ (_27191_, _13220_, _13219_);
  and _44400_ (_13221_, _12442_, _23583_);
  and _44401_ (_13222_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  or _44402_ (_04679_, _13222_, _13221_);
  and _44403_ (_13223_, _05465_, _24089_);
  and _44404_ (_13224_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or _44405_ (_27069_, _13224_, _13223_);
  and _44406_ (_13225_, _12442_, _23887_);
  and _44407_ (_13226_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  or _44408_ (_26994_, _13226_, _13225_);
  and _44409_ (_13227_, _12438_, _24134_);
  and _44410_ (_13228_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or _44411_ (_04713_, _13228_, _13227_);
  and _44412_ (_13229_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and _44413_ (_13230_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _44414_ (_13231_, _13230_, _13229_);
  and _44415_ (_13232_, _13231_, _09792_);
  and _44416_ (_13233_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and _44417_ (_13234_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _44418_ (_13235_, _13234_, _13233_);
  and _44419_ (_13236_, _13235_, _05549_);
  or _44420_ (_13237_, _13236_, _13232_);
  or _44421_ (_13238_, _13237_, _09791_);
  and _44422_ (_13239_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and _44423_ (_13240_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _44424_ (_13241_, _13240_, _13239_);
  and _44425_ (_13242_, _13241_, _09792_);
  and _44426_ (_13243_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and _44427_ (_13244_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _44428_ (_13245_, _13244_, _13243_);
  and _44429_ (_13246_, _13245_, _05549_);
  or _44430_ (_13247_, _13246_, _13242_);
  or _44431_ (_13248_, _13247_, _05535_);
  and _44432_ (_13249_, _13248_, _09805_);
  and _44433_ (_13250_, _13249_, _13238_);
  or _44434_ (_13251_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _44435_ (_13252_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and _44436_ (_13253_, _13252_, _13251_);
  and _44437_ (_13254_, _13253_, _09792_);
  or _44438_ (_13255_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _44439_ (_13256_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and _44440_ (_13257_, _13256_, _13255_);
  and _44441_ (_13258_, _13257_, _05549_);
  or _44442_ (_13259_, _13258_, _13254_);
  or _44443_ (_13260_, _13259_, _09791_);
  or _44444_ (_13261_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _44445_ (_13262_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and _44446_ (_13263_, _13262_, _13261_);
  and _44447_ (_13264_, _13263_, _09792_);
  or _44448_ (_13265_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _44449_ (_13266_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and _44450_ (_13267_, _13266_, _13265_);
  and _44451_ (_13268_, _13267_, _05549_);
  or _44452_ (_13269_, _13268_, _13264_);
  or _44453_ (_13270_, _13269_, _05535_);
  and _44454_ (_13271_, _13270_, _05542_);
  and _44455_ (_13272_, _13271_, _13260_);
  or _44456_ (_13273_, _13272_, _13250_);
  and _44457_ (_13274_, _13273_, _05518_);
  and _44458_ (_13275_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and _44459_ (_13276_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _44460_ (_13277_, _13276_, _13275_);
  and _44461_ (_13278_, _13277_, _09792_);
  and _44462_ (_13279_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and _44463_ (_13280_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _44464_ (_13281_, _13280_, _13279_);
  and _44465_ (_13282_, _13281_, _05549_);
  or _44466_ (_13283_, _13282_, _13278_);
  or _44467_ (_13284_, _13283_, _09791_);
  and _44468_ (_13285_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and _44469_ (_13286_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _44470_ (_13287_, _13286_, _13285_);
  and _44471_ (_13288_, _13287_, _09792_);
  and _44472_ (_13289_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and _44473_ (_13290_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _44474_ (_13291_, _13290_, _13289_);
  and _44475_ (_13292_, _13291_, _05549_);
  or _44476_ (_13293_, _13292_, _13288_);
  or _44477_ (_13294_, _13293_, _05535_);
  and _44478_ (_13295_, _13294_, _09805_);
  and _44479_ (_13296_, _13295_, _13284_);
  or _44480_ (_13297_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _44481_ (_13298_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and _44482_ (_13299_, _13298_, _05549_);
  and _44483_ (_13300_, _13299_, _13297_);
  or _44484_ (_13301_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _44485_ (_13302_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and _44486_ (_13303_, _13302_, _09792_);
  and _44487_ (_13304_, _13303_, _13301_);
  or _44488_ (_13305_, _13304_, _13300_);
  or _44489_ (_13306_, _13305_, _09791_);
  or _44490_ (_13307_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _44491_ (_13308_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and _44492_ (_13309_, _13308_, _05549_);
  and _44493_ (_13310_, _13309_, _13307_);
  or _44494_ (_13311_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _44495_ (_13312_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and _44496_ (_13313_, _13312_, _09792_);
  and _44497_ (_13314_, _13313_, _13311_);
  or _44498_ (_13315_, _13314_, _13310_);
  or _44499_ (_13316_, _13315_, _05535_);
  and _44500_ (_13317_, _13316_, _05542_);
  and _44501_ (_13318_, _13317_, _13306_);
  or _44502_ (_13319_, _13318_, _13296_);
  and _44503_ (_13320_, _13319_, _09850_);
  or _44504_ (_13321_, _13320_, _13274_);
  and _44505_ (_13322_, _13321_, _09790_);
  and _44506_ (_13323_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _44507_ (_13324_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _44508_ (_13325_, _13324_, _13323_);
  and _44509_ (_13326_, _13325_, _09792_);
  and _44510_ (_13327_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _44511_ (_13328_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _44512_ (_13329_, _13328_, _13327_);
  and _44513_ (_13330_, _13329_, _05549_);
  or _44514_ (_13331_, _13330_, _13326_);
  and _44515_ (_13332_, _13331_, _05535_);
  and _44516_ (_13333_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _44517_ (_13334_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _44518_ (_13335_, _13334_, _13333_);
  and _44519_ (_13336_, _13335_, _09792_);
  and _44520_ (_13337_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _44521_ (_13338_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _44522_ (_13339_, _13338_, _13337_);
  and _44523_ (_13340_, _13339_, _05549_);
  or _44524_ (_13341_, _13340_, _13336_);
  and _44525_ (_13342_, _13341_, _09791_);
  or _44526_ (_13343_, _13342_, _13332_);
  and _44527_ (_13344_, _13343_, _09805_);
  or _44528_ (_13345_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _44529_ (_13346_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _44530_ (_13347_, _13346_, _05549_);
  and _44531_ (_13348_, _13347_, _13345_);
  or _44532_ (_13349_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _44533_ (_13350_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _44534_ (_13351_, _13350_, _09792_);
  and _44535_ (_13352_, _13351_, _13349_);
  or _44536_ (_13353_, _13352_, _13348_);
  and _44537_ (_13354_, _13353_, _05535_);
  or _44538_ (_13355_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _44539_ (_13356_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _44540_ (_13357_, _13356_, _05549_);
  and _44541_ (_13358_, _13357_, _13355_);
  or _44542_ (_13359_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _44543_ (_13360_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _44544_ (_13361_, _13360_, _09792_);
  and _44545_ (_13362_, _13361_, _13359_);
  or _44546_ (_13363_, _13362_, _13358_);
  and _44547_ (_13364_, _13363_, _09791_);
  or _44548_ (_13365_, _13364_, _13354_);
  and _44549_ (_13366_, _13365_, _05542_);
  or _44550_ (_13367_, _13366_, _13344_);
  and _44551_ (_13368_, _13367_, _09850_);
  and _44552_ (_13369_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and _44553_ (_13370_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _44554_ (_13371_, _13370_, _13369_);
  and _44555_ (_13372_, _13371_, _09792_);
  and _44556_ (_13373_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and _44557_ (_13374_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _44558_ (_13375_, _13374_, _13373_);
  and _44559_ (_13376_, _13375_, _05549_);
  or _44560_ (_13377_, _13376_, _13372_);
  and _44561_ (_13378_, _13377_, _05535_);
  and _44562_ (_13379_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and _44563_ (_13380_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _44564_ (_13381_, _13380_, _13379_);
  and _44565_ (_13382_, _13381_, _09792_);
  and _44566_ (_13383_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and _44567_ (_13384_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _44568_ (_13385_, _13384_, _13383_);
  and _44569_ (_13386_, _13385_, _05549_);
  or _44570_ (_13387_, _13386_, _13382_);
  and _44571_ (_13388_, _13387_, _09791_);
  or _44572_ (_13389_, _13388_, _13378_);
  and _44573_ (_13390_, _13389_, _09805_);
  or _44574_ (_13391_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _44575_ (_13392_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and _44576_ (_13393_, _13392_, _13391_);
  and _44577_ (_13394_, _13393_, _09792_);
  or _44578_ (_13395_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _44579_ (_13396_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and _44580_ (_13397_, _13396_, _13395_);
  and _44581_ (_13398_, _13397_, _05549_);
  or _44582_ (_13399_, _13398_, _13394_);
  and _44583_ (_13400_, _13399_, _05535_);
  or _44584_ (_13401_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _44585_ (_13402_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and _44586_ (_13403_, _13402_, _13401_);
  and _44587_ (_13404_, _13403_, _09792_);
  or _44588_ (_13405_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _44589_ (_13406_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and _44590_ (_13407_, _13406_, _13405_);
  and _44591_ (_13408_, _13407_, _05549_);
  or _44592_ (_13409_, _13408_, _13404_);
  and _44593_ (_13410_, _13409_, _09791_);
  or _44594_ (_13411_, _13410_, _13400_);
  and _44595_ (_13412_, _13411_, _05542_);
  or _44596_ (_13413_, _13412_, _13390_);
  and _44597_ (_13414_, _13413_, _05518_);
  or _44598_ (_13415_, _13414_, _13368_);
  and _44599_ (_13416_, _13415_, _05520_);
  or _44600_ (_13417_, _13416_, _13322_);
  or _44601_ (_13418_, _13417_, _05526_);
  and _44602_ (_13419_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and _44603_ (_13420_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _44604_ (_13421_, _13420_, _13419_);
  and _44605_ (_13422_, _13421_, _09792_);
  and _44606_ (_13423_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and _44607_ (_13424_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _44608_ (_13425_, _13424_, _13423_);
  and _44609_ (_13426_, _13425_, _05549_);
  or _44610_ (_13427_, _13426_, _13422_);
  or _44611_ (_13428_, _13427_, _09791_);
  and _44612_ (_13429_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and _44613_ (_13430_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _44614_ (_13431_, _13430_, _13429_);
  and _44615_ (_13432_, _13431_, _09792_);
  and _44616_ (_13433_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and _44617_ (_13434_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _44618_ (_13435_, _13434_, _13433_);
  and _44619_ (_13436_, _13435_, _05549_);
  or _44620_ (_13437_, _13436_, _13432_);
  or _44621_ (_13438_, _13437_, _05535_);
  and _44622_ (_13439_, _13438_, _09805_);
  and _44623_ (_13440_, _13439_, _13428_);
  or _44624_ (_13441_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _44625_ (_13442_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and _44626_ (_13443_, _13442_, _05549_);
  and _44627_ (_13444_, _13443_, _13441_);
  or _44628_ (_13445_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _44629_ (_13446_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and _44630_ (_13447_, _13446_, _09792_);
  and _44631_ (_13448_, _13447_, _13445_);
  or _44632_ (_13449_, _13448_, _13444_);
  or _44633_ (_13450_, _13449_, _09791_);
  or _44634_ (_13451_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _44635_ (_13452_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and _44636_ (_13453_, _13452_, _05549_);
  and _44637_ (_13454_, _13453_, _13451_);
  or _44638_ (_13455_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _44639_ (_13456_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and _44640_ (_13457_, _13456_, _09792_);
  and _44641_ (_13458_, _13457_, _13455_);
  or _44642_ (_13459_, _13458_, _13454_);
  or _44643_ (_13460_, _13459_, _05535_);
  and _44644_ (_13461_, _13460_, _05542_);
  and _44645_ (_13462_, _13461_, _13450_);
  or _44646_ (_13463_, _13462_, _13440_);
  and _44647_ (_13464_, _13463_, _09850_);
  and _44648_ (_13465_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and _44649_ (_13466_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _44650_ (_13467_, _13466_, _13465_);
  and _44651_ (_13468_, _13467_, _09792_);
  and _44652_ (_13469_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and _44653_ (_13470_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _44654_ (_13471_, _13470_, _13469_);
  and _44655_ (_13472_, _13471_, _05549_);
  or _44656_ (_13473_, _13472_, _13468_);
  or _44657_ (_13474_, _13473_, _09791_);
  and _44658_ (_13475_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _44659_ (_13476_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _44660_ (_13477_, _13476_, _13475_);
  and _44661_ (_13478_, _13477_, _09792_);
  and _44662_ (_13479_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _44663_ (_13480_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _44664_ (_13481_, _13480_, _13479_);
  and _44665_ (_13482_, _13481_, _05549_);
  or _44666_ (_13483_, _13482_, _13478_);
  or _44667_ (_13484_, _13483_, _05535_);
  and _44668_ (_13485_, _13484_, _09805_);
  and _44669_ (_13486_, _13485_, _13474_);
  or _44670_ (_13487_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _44671_ (_13488_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and _44672_ (_13489_, _13488_, _13487_);
  and _44673_ (_13490_, _13489_, _09792_);
  or _44674_ (_13491_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _44675_ (_13492_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and _44676_ (_13493_, _13492_, _13491_);
  and _44677_ (_13494_, _13493_, _05549_);
  or _44678_ (_13495_, _13494_, _13490_);
  or _44679_ (_13496_, _13495_, _09791_);
  or _44680_ (_13497_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _44681_ (_13498_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and _44682_ (_13499_, _13498_, _13497_);
  and _44683_ (_13500_, _13499_, _09792_);
  or _44684_ (_13501_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _44685_ (_13502_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and _44686_ (_13503_, _13502_, _13501_);
  and _44687_ (_13504_, _13503_, _05549_);
  or _44688_ (_13505_, _13504_, _13500_);
  or _44689_ (_13506_, _13505_, _05535_);
  and _44690_ (_13507_, _13506_, _05542_);
  and _44691_ (_13508_, _13507_, _13496_);
  or _44692_ (_13509_, _13508_, _13486_);
  and _44693_ (_13510_, _13509_, _05518_);
  or _44694_ (_13511_, _13510_, _13464_);
  and _44695_ (_13512_, _13511_, _09790_);
  or _44696_ (_13513_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _44697_ (_13514_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and _44698_ (_13515_, _13514_, _13513_);
  and _44699_ (_13516_, _13515_, _09792_);
  or _44700_ (_13517_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _44701_ (_13518_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and _44702_ (_13519_, _13518_, _13517_);
  and _44703_ (_13520_, _13519_, _05549_);
  or _44704_ (_13521_, _13520_, _13516_);
  and _44705_ (_13522_, _13521_, _09791_);
  or _44706_ (_13523_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _44707_ (_13524_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and _44708_ (_13525_, _13524_, _13523_);
  and _44709_ (_13526_, _13525_, _09792_);
  or _44710_ (_13527_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _44711_ (_13528_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and _44712_ (_13529_, _13528_, _13527_);
  and _44713_ (_13530_, _13529_, _05549_);
  or _44714_ (_13531_, _13530_, _13526_);
  and _44715_ (_13532_, _13531_, _05535_);
  or _44716_ (_13533_, _13532_, _13522_);
  and _44717_ (_13534_, _13533_, _05542_);
  and _44718_ (_13535_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and _44719_ (_13536_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _44720_ (_13537_, _13536_, _13535_);
  and _44721_ (_13538_, _13537_, _09792_);
  and _44722_ (_13539_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and _44723_ (_13540_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _44724_ (_13541_, _13540_, _13539_);
  and _44725_ (_13542_, _13541_, _05549_);
  or _44726_ (_13543_, _13542_, _13538_);
  and _44727_ (_13544_, _13543_, _09791_);
  and _44728_ (_13545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and _44729_ (_13546_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _44730_ (_13547_, _13546_, _13545_);
  and _44731_ (_13548_, _13547_, _09792_);
  and _44732_ (_13549_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and _44733_ (_13550_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _44734_ (_13551_, _13550_, _13549_);
  and _44735_ (_13552_, _13551_, _05549_);
  or _44736_ (_13553_, _13552_, _13548_);
  and _44737_ (_13554_, _13553_, _05535_);
  or _44738_ (_13555_, _13554_, _13544_);
  and _44739_ (_13556_, _13555_, _09805_);
  or _44740_ (_13557_, _13556_, _13534_);
  and _44741_ (_13558_, _13557_, _05518_);
  or _44742_ (_13559_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _44743_ (_13560_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and _44744_ (_13561_, _13560_, _05549_);
  and _44745_ (_13562_, _13561_, _13559_);
  or _44746_ (_13563_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or _44747_ (_13564_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and _44748_ (_13565_, _13564_, _09792_);
  and _44749_ (_13566_, _13565_, _13563_);
  or _44750_ (_13567_, _13566_, _13562_);
  and _44751_ (_13568_, _13567_, _09791_);
  or _44752_ (_13569_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _44753_ (_13570_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and _44754_ (_13571_, _13570_, _05549_);
  and _44755_ (_13572_, _13571_, _13569_);
  or _44756_ (_13573_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or _44757_ (_13574_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and _44758_ (_13575_, _13574_, _09792_);
  and _44759_ (_13576_, _13575_, _13573_);
  or _44760_ (_13577_, _13576_, _13572_);
  and _44761_ (_13578_, _13577_, _05535_);
  or _44762_ (_13579_, _13578_, _13568_);
  and _44763_ (_13580_, _13579_, _05542_);
  and _44764_ (_13581_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and _44765_ (_13582_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or _44766_ (_13583_, _13582_, _13581_);
  and _44767_ (_13584_, _13583_, _09792_);
  and _44768_ (_13585_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and _44769_ (_13586_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or _44770_ (_13587_, _13586_, _13585_);
  and _44771_ (_13588_, _13587_, _05549_);
  or _44772_ (_13589_, _13588_, _13584_);
  and _44773_ (_13590_, _13589_, _09791_);
  and _44774_ (_13591_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and _44775_ (_13592_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or _44776_ (_13593_, _13592_, _13591_);
  and _44777_ (_13594_, _13593_, _09792_);
  and _44778_ (_13595_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and _44779_ (_13596_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _44780_ (_13597_, _13596_, _13595_);
  and _44781_ (_13598_, _13597_, _05549_);
  or _44782_ (_13599_, _13598_, _13594_);
  and _44783_ (_13600_, _13599_, _05535_);
  or _44784_ (_13601_, _13600_, _13590_);
  and _44785_ (_13602_, _13601_, _09805_);
  or _44786_ (_13603_, _13602_, _13580_);
  and _44787_ (_13604_, _13603_, _09850_);
  or _44788_ (_13605_, _13604_, _13558_);
  and _44789_ (_13606_, _13605_, _05520_);
  or _44790_ (_13607_, _13606_, _13512_);
  or _44791_ (_13608_, _13607_, _10033_);
  and _44792_ (_13609_, _13608_, _13418_);
  or _44793_ (_13610_, _13609_, _00143_);
  and _44794_ (_13611_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and _44795_ (_13612_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _44796_ (_13613_, _13612_, _13611_);
  and _44797_ (_13614_, _13613_, _09792_);
  and _44798_ (_13615_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and _44799_ (_13616_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _44800_ (_13617_, _13616_, _13615_);
  and _44801_ (_13618_, _13617_, _05549_);
  or _44802_ (_13619_, _13618_, _13614_);
  or _44803_ (_13620_, _13619_, _09791_);
  and _44804_ (_13621_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and _44805_ (_13622_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _44806_ (_13623_, _13622_, _13621_);
  and _44807_ (_13624_, _13623_, _09792_);
  and _44808_ (_13625_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and _44809_ (_13626_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _44810_ (_13627_, _13626_, _13625_);
  and _44811_ (_13628_, _13627_, _05549_);
  or _44812_ (_13629_, _13628_, _13624_);
  or _44813_ (_13630_, _13629_, _05535_);
  and _44814_ (_13631_, _13630_, _09805_);
  and _44815_ (_13632_, _13631_, _13620_);
  or _44816_ (_13633_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _44817_ (_13634_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and _44818_ (_13635_, _13634_, _13633_);
  and _44819_ (_13636_, _13635_, _09792_);
  or _44820_ (_13637_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _44821_ (_13638_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and _44822_ (_13639_, _13638_, _13637_);
  and _44823_ (_13640_, _13639_, _05549_);
  or _44824_ (_13641_, _13640_, _13636_);
  or _44825_ (_13642_, _13641_, _09791_);
  or _44826_ (_13643_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _44827_ (_13644_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and _44828_ (_13645_, _13644_, _13643_);
  and _44829_ (_13646_, _13645_, _09792_);
  or _44830_ (_13647_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _44831_ (_13648_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and _44832_ (_13649_, _13648_, _13647_);
  and _44833_ (_13650_, _13649_, _05549_);
  or _44834_ (_13651_, _13650_, _13646_);
  or _44835_ (_13652_, _13651_, _05535_);
  and _44836_ (_13653_, _13652_, _05542_);
  and _44837_ (_13654_, _13653_, _13642_);
  or _44838_ (_13655_, _13654_, _13632_);
  and _44839_ (_13656_, _13655_, _05518_);
  and _44840_ (_13657_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _44841_ (_13658_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or _44842_ (_13659_, _13658_, _13657_);
  and _44843_ (_13660_, _13659_, _09792_);
  and _44844_ (_13661_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _44845_ (_13662_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or _44846_ (_13663_, _13662_, _13661_);
  and _44847_ (_13664_, _13663_, _05549_);
  or _44848_ (_13665_, _13664_, _13660_);
  or _44849_ (_13666_, _13665_, _09791_);
  and _44850_ (_13667_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _44851_ (_13668_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _44852_ (_13669_, _13668_, _13667_);
  and _44853_ (_13670_, _13669_, _09792_);
  and _44854_ (_13671_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _44855_ (_13672_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or _44856_ (_13673_, _13672_, _13671_);
  and _44857_ (_13674_, _13673_, _05549_);
  or _44858_ (_13675_, _13674_, _13670_);
  or _44859_ (_13676_, _13675_, _05535_);
  and _44860_ (_13677_, _13676_, _09805_);
  and _44861_ (_13678_, _13677_, _13666_);
  or _44862_ (_13679_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or _44863_ (_13680_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _44864_ (_13681_, _13680_, _05549_);
  and _44865_ (_13682_, _13681_, _13679_);
  or _44866_ (_13683_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _44867_ (_13684_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and _44868_ (_13685_, _13684_, _09792_);
  and _44869_ (_13686_, _13685_, _13683_);
  or _44870_ (_13687_, _13686_, _13682_);
  or _44871_ (_13688_, _13687_, _09791_);
  or _44872_ (_13689_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or _44873_ (_13690_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _44874_ (_13691_, _13690_, _05549_);
  and _44875_ (_13692_, _13691_, _13689_);
  or _44876_ (_13693_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _44877_ (_13694_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _44878_ (_13695_, _13694_, _09792_);
  and _44879_ (_13696_, _13695_, _13693_);
  or _44880_ (_13697_, _13696_, _13692_);
  or _44881_ (_13698_, _13697_, _05535_);
  and _44882_ (_13699_, _13698_, _05542_);
  and _44883_ (_13700_, _13699_, _13688_);
  or _44884_ (_13701_, _13700_, _13678_);
  and _44885_ (_13702_, _13701_, _09850_);
  or _44886_ (_13703_, _13702_, _13656_);
  and _44887_ (_13704_, _13703_, _09790_);
  and _44888_ (_13705_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and _44889_ (_13706_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or _44890_ (_13707_, _13706_, _13705_);
  and _44891_ (_13708_, _13707_, _09792_);
  and _44892_ (_13709_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and _44893_ (_13710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or _44894_ (_13711_, _13710_, _13709_);
  and _44895_ (_13712_, _13711_, _05549_);
  or _44896_ (_13713_, _13712_, _13708_);
  and _44897_ (_13714_, _13713_, _05535_);
  and _44898_ (_13715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and _44899_ (_13716_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or _44900_ (_13717_, _13716_, _13715_);
  and _44901_ (_13718_, _13717_, _09792_);
  and _44902_ (_13719_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _44903_ (_13720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or _44904_ (_13721_, _13720_, _13719_);
  and _44905_ (_13722_, _13721_, _05549_);
  or _44906_ (_13723_, _13722_, _13718_);
  and _44907_ (_13724_, _13723_, _09791_);
  or _44908_ (_13725_, _13724_, _13714_);
  and _44909_ (_13726_, _13725_, _09805_);
  or _44910_ (_13727_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or _44911_ (_13728_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and _44912_ (_13729_, _13728_, _05549_);
  and _44913_ (_13730_, _13729_, _13727_);
  or _44914_ (_13731_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or _44915_ (_13732_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and _44916_ (_13733_, _13732_, _09792_);
  and _44917_ (_13734_, _13733_, _13731_);
  or _44918_ (_13735_, _13734_, _13730_);
  and _44919_ (_13736_, _13735_, _05535_);
  or _44920_ (_13737_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or _44921_ (_13738_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and _44922_ (_13739_, _13738_, _05549_);
  and _44923_ (_13740_, _13739_, _13737_);
  or _44924_ (_13741_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or _44925_ (_13742_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and _44926_ (_13743_, _13742_, _09792_);
  and _44927_ (_13744_, _13743_, _13741_);
  or _44928_ (_13745_, _13744_, _13740_);
  and _44929_ (_13746_, _13745_, _09791_);
  or _44930_ (_13747_, _13746_, _13736_);
  and _44931_ (_13748_, _13747_, _05542_);
  or _44932_ (_13749_, _13748_, _13726_);
  and _44933_ (_13750_, _13749_, _09850_);
  and _44934_ (_13751_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _44935_ (_13752_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _44936_ (_13753_, _13752_, _13751_);
  and _44937_ (_13754_, _13753_, _09792_);
  and _44938_ (_13755_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and _44939_ (_13756_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _44940_ (_13757_, _13756_, _13755_);
  and _44941_ (_13758_, _13757_, _05549_);
  or _44942_ (_13759_, _13758_, _13754_);
  and _44943_ (_13760_, _13759_, _05535_);
  and _44944_ (_13761_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _44945_ (_13762_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _44946_ (_13763_, _13762_, _13761_);
  and _44947_ (_13764_, _13763_, _09792_);
  and _44948_ (_13765_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and _44949_ (_13766_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _44950_ (_13767_, _13766_, _13765_);
  and _44951_ (_13768_, _13767_, _05549_);
  or _44952_ (_13769_, _13768_, _13764_);
  and _44953_ (_13770_, _13769_, _09791_);
  or _44954_ (_13771_, _13770_, _13760_);
  and _44955_ (_13772_, _13771_, _09805_);
  or _44956_ (_13773_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _44957_ (_13774_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and _44958_ (_13775_, _13774_, _13773_);
  and _44959_ (_13776_, _13775_, _09792_);
  or _44960_ (_13777_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _44961_ (_13778_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _44962_ (_13779_, _13778_, _13777_);
  and _44963_ (_13780_, _13779_, _05549_);
  or _44964_ (_13781_, _13780_, _13776_);
  and _44965_ (_13782_, _13781_, _05535_);
  or _44966_ (_13783_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _44967_ (_13784_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and _44968_ (_13785_, _13784_, _13783_);
  and _44969_ (_13786_, _13785_, _09792_);
  or _44970_ (_13787_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _44971_ (_13788_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _44972_ (_13789_, _13788_, _13787_);
  and _44973_ (_13790_, _13789_, _05549_);
  or _44974_ (_13791_, _13790_, _13786_);
  and _44975_ (_13792_, _13791_, _09791_);
  or _44976_ (_13793_, _13792_, _13782_);
  and _44977_ (_13794_, _13793_, _05542_);
  or _44978_ (_13795_, _13794_, _13772_);
  and _44979_ (_13796_, _13795_, _05518_);
  or _44980_ (_13797_, _13796_, _13750_);
  and _44981_ (_13798_, _13797_, _05520_);
  or _44982_ (_13799_, _13798_, _13704_);
  or _44983_ (_13800_, _13799_, _05526_);
  and _44984_ (_13801_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and _44985_ (_13802_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _44986_ (_13803_, _13802_, _13801_);
  and _44987_ (_13804_, _13803_, _09792_);
  and _44988_ (_13805_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and _44989_ (_13806_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _44990_ (_13807_, _13806_, _13805_);
  and _44991_ (_13808_, _13807_, _05549_);
  or _44992_ (_13809_, _13808_, _13804_);
  or _44993_ (_13810_, _13809_, _09791_);
  and _44994_ (_13811_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and _44995_ (_13812_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _44996_ (_13813_, _13812_, _13811_);
  and _44997_ (_13814_, _13813_, _09792_);
  and _44998_ (_13815_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and _44999_ (_13816_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _45000_ (_13817_, _13816_, _13815_);
  and _45001_ (_13818_, _13817_, _05549_);
  or _45002_ (_13819_, _13818_, _13814_);
  or _45003_ (_13820_, _13819_, _05535_);
  and _45004_ (_13821_, _13820_, _09805_);
  and _45005_ (_13822_, _13821_, _13810_);
  or _45006_ (_13823_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _45007_ (_13824_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and _45008_ (_13825_, _13824_, _05549_);
  and _45009_ (_13826_, _13825_, _13823_);
  or _45010_ (_13827_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _45011_ (_13828_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and _45012_ (_13829_, _13828_, _09792_);
  and _45013_ (_13830_, _13829_, _13827_);
  or _45014_ (_13831_, _13830_, _13826_);
  or _45015_ (_13832_, _13831_, _09791_);
  or _45016_ (_13833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _45017_ (_13834_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and _45018_ (_13835_, _13834_, _05549_);
  and _45019_ (_13836_, _13835_, _13833_);
  or _45020_ (_13837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _45021_ (_13838_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and _45022_ (_13839_, _13838_, _09792_);
  and _45023_ (_13840_, _13839_, _13837_);
  or _45024_ (_13841_, _13840_, _13836_);
  or _45025_ (_13842_, _13841_, _05535_);
  and _45026_ (_13843_, _13842_, _05542_);
  and _45027_ (_13844_, _13843_, _13832_);
  or _45028_ (_13845_, _13844_, _13822_);
  and _45029_ (_13846_, _13845_, _09850_);
  and _45030_ (_13847_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _45031_ (_13848_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _45032_ (_13849_, _13848_, _13847_);
  and _45033_ (_13850_, _13849_, _09792_);
  and _45034_ (_13851_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _45035_ (_13852_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or _45036_ (_13853_, _13852_, _13851_);
  and _45037_ (_13854_, _13853_, _05549_);
  or _45038_ (_13855_, _13854_, _13850_);
  or _45039_ (_13856_, _13855_, _09791_);
  and _45040_ (_13857_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _45041_ (_13858_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or _45042_ (_13859_, _13858_, _13857_);
  and _45043_ (_13860_, _13859_, _09792_);
  and _45044_ (_13861_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _45045_ (_13862_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _45046_ (_13863_, _13862_, _13861_);
  and _45047_ (_13864_, _13863_, _05549_);
  or _45048_ (_13865_, _13864_, _13860_);
  or _45049_ (_13866_, _13865_, _05535_);
  and _45050_ (_13867_, _13866_, _09805_);
  and _45051_ (_13868_, _13867_, _13856_);
  or _45052_ (_13869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or _45053_ (_13870_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _45054_ (_13871_, _13870_, _13869_);
  and _45055_ (_13872_, _13871_, _09792_);
  or _45056_ (_13873_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or _45057_ (_13874_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and _45058_ (_13875_, _13874_, _13873_);
  and _45059_ (_13876_, _13875_, _05549_);
  or _45060_ (_13877_, _13876_, _13872_);
  or _45061_ (_13878_, _13877_, _09791_);
  or _45062_ (_13879_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _45063_ (_13880_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _45064_ (_13881_, _13880_, _13879_);
  and _45065_ (_13882_, _13881_, _09792_);
  or _45066_ (_13883_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _45067_ (_13884_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and _45068_ (_13885_, _13884_, _13883_);
  and _45069_ (_13886_, _13885_, _05549_);
  or _45070_ (_13887_, _13886_, _13882_);
  or _45071_ (_13888_, _13887_, _05535_);
  and _45072_ (_13889_, _13888_, _05542_);
  and _45073_ (_13890_, _13889_, _13878_);
  or _45074_ (_13891_, _13890_, _13868_);
  and _45075_ (_13892_, _13891_, _05518_);
  or _45076_ (_13893_, _13892_, _13846_);
  and _45077_ (_13894_, _13893_, _09790_);
  or _45078_ (_13895_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _45079_ (_13896_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _45080_ (_13897_, _13896_, _13895_);
  and _45081_ (_13898_, _13897_, _09792_);
  or _45082_ (_13899_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _45083_ (_13900_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and _45084_ (_13901_, _13900_, _13899_);
  and _45085_ (_13902_, _13901_, _05549_);
  or _45086_ (_13903_, _13902_, _13898_);
  and _45087_ (_13904_, _13903_, _09791_);
  or _45088_ (_13905_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or _45089_ (_13906_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and _45090_ (_13907_, _13906_, _13905_);
  and _45091_ (_13908_, _13907_, _09792_);
  or _45092_ (_13909_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or _45093_ (_13910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _45094_ (_13911_, _13910_, _13909_);
  and _45095_ (_13912_, _13911_, _05549_);
  or _45096_ (_13913_, _13912_, _13908_);
  and _45097_ (_13914_, _13913_, _05535_);
  or _45098_ (_13915_, _13914_, _13904_);
  and _45099_ (_13916_, _13915_, _05542_);
  and _45100_ (_13917_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _45101_ (_13918_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or _45102_ (_13919_, _13918_, _13917_);
  and _45103_ (_13920_, _13919_, _09792_);
  and _45104_ (_13921_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _45105_ (_13922_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _45106_ (_13923_, _13922_, _13921_);
  and _45107_ (_13924_, _13923_, _05549_);
  or _45108_ (_13925_, _13924_, _13920_);
  and _45109_ (_13926_, _13925_, _09791_);
  and _45110_ (_13927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _45111_ (_13928_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or _45112_ (_13929_, _13928_, _13927_);
  and _45113_ (_13930_, _13929_, _09792_);
  and _45114_ (_13931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and _45115_ (_13932_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _45116_ (_13933_, _13932_, _13931_);
  and _45117_ (_13934_, _13933_, _05549_);
  or _45118_ (_13935_, _13934_, _13930_);
  and _45119_ (_13936_, _13935_, _05535_);
  or _45120_ (_13937_, _13936_, _13926_);
  and _45121_ (_13938_, _13937_, _09805_);
  or _45122_ (_13939_, _13938_, _13916_);
  and _45123_ (_13940_, _13939_, _05518_);
  or _45124_ (_13941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _45125_ (_13942_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and _45126_ (_13943_, _13942_, _05549_);
  and _45127_ (_13944_, _13943_, _13941_);
  or _45128_ (_13945_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _45129_ (_13946_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and _45130_ (_13947_, _13946_, _09792_);
  and _45131_ (_13948_, _13947_, _13945_);
  or _45132_ (_13949_, _13948_, _13944_);
  and _45133_ (_13950_, _13949_, _09791_);
  or _45134_ (_13951_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _45135_ (_13952_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _45136_ (_13953_, _13952_, _05549_);
  and _45137_ (_13954_, _13953_, _13951_);
  or _45138_ (_13955_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _45139_ (_13956_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and _45140_ (_13957_, _13956_, _09792_);
  and _45141_ (_13958_, _13957_, _13955_);
  or _45142_ (_13959_, _13958_, _13954_);
  and _45143_ (_13960_, _13959_, _05535_);
  or _45144_ (_13961_, _13960_, _13950_);
  and _45145_ (_13962_, _13961_, _05542_);
  and _45146_ (_13963_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _45147_ (_13964_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _45148_ (_13965_, _13964_, _13963_);
  and _45149_ (_13966_, _13965_, _09792_);
  and _45150_ (_13967_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and _45151_ (_13968_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _45152_ (_13969_, _13968_, _13967_);
  and _45153_ (_13970_, _13969_, _05549_);
  or _45154_ (_13971_, _13970_, _13966_);
  and _45155_ (_13972_, _13971_, _09791_);
  and _45156_ (_13973_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and _45157_ (_13974_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _45158_ (_13975_, _13974_, _13973_);
  and _45159_ (_13976_, _13975_, _09792_);
  and _45160_ (_13977_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and _45161_ (_13978_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _45162_ (_13979_, _13978_, _13977_);
  and _45163_ (_13980_, _13979_, _05549_);
  or _45164_ (_13981_, _13980_, _13976_);
  and _45165_ (_13982_, _13981_, _05535_);
  or _45166_ (_13983_, _13982_, _13972_);
  and _45167_ (_13984_, _13983_, _09805_);
  or _45168_ (_13985_, _13984_, _13962_);
  and _45169_ (_13986_, _13985_, _09850_);
  or _45170_ (_13987_, _13986_, _13940_);
  and _45171_ (_13988_, _13987_, _05520_);
  or _45172_ (_13989_, _13988_, _13894_);
  or _45173_ (_13990_, _13989_, _10033_);
  and _45174_ (_13991_, _13990_, _13800_);
  or _45175_ (_13992_, _13991_, _04413_);
  and _45176_ (_13993_, _13992_, _13610_);
  or _45177_ (_13994_, _13993_, _05563_);
  or _45178_ (_13995_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and _45179_ (_13996_, _13995_, _22731_);
  and _45180_ (_04717_, _13996_, _13994_);
  and _45181_ (_13997_, _12438_, _24051_);
  and _45182_ (_13998_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or _45183_ (_04720_, _13998_, _13997_);
  and _45184_ (_13999_, _12438_, _24089_);
  and _45185_ (_14000_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or _45186_ (_04728_, _14000_, _13999_);
  and _45187_ (_14001_, _07013_, _24134_);
  and _45188_ (_14002_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _45189_ (_04731_, _14002_, _14001_);
  and _45190_ (_14003_, _12442_, _24051_);
  and _45191_ (_14004_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  or _45192_ (_04734_, _14004_, _14003_);
  and _45193_ (_14005_, _12442_, _23996_);
  and _45194_ (_14006_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or _45195_ (_04740_, _14006_, _14005_);
  and _45196_ (_14007_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and _45197_ (_14008_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _45198_ (_14009_, _14008_, _14007_);
  and _45199_ (_14010_, _14009_, _09792_);
  and _45200_ (_14011_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and _45201_ (_14012_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _45202_ (_14013_, _14012_, _14011_);
  and _45203_ (_14014_, _14013_, _05549_);
  or _45204_ (_14015_, _14014_, _14010_);
  or _45205_ (_14016_, _14015_, _09791_);
  and _45206_ (_14017_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and _45207_ (_14018_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _45208_ (_14019_, _14018_, _14017_);
  and _45209_ (_14020_, _14019_, _09792_);
  and _45210_ (_14021_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and _45211_ (_14022_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _45212_ (_14023_, _14022_, _14021_);
  and _45213_ (_14024_, _14023_, _05549_);
  or _45214_ (_14025_, _14024_, _14020_);
  or _45215_ (_14026_, _14025_, _05535_);
  and _45216_ (_14027_, _14026_, _09805_);
  and _45217_ (_14028_, _14027_, _14016_);
  or _45218_ (_14029_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _45219_ (_14030_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and _45220_ (_14031_, _14030_, _14029_);
  and _45221_ (_14032_, _14031_, _09792_);
  or _45222_ (_14033_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _45223_ (_14034_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and _45224_ (_14035_, _14034_, _14033_);
  and _45225_ (_14036_, _14035_, _05549_);
  or _45226_ (_14037_, _14036_, _14032_);
  or _45227_ (_14038_, _14037_, _09791_);
  or _45228_ (_14039_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _45229_ (_14040_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and _45230_ (_14041_, _14040_, _14039_);
  and _45231_ (_14042_, _14041_, _09792_);
  or _45232_ (_14043_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _45233_ (_14044_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and _45234_ (_14045_, _14044_, _14043_);
  and _45235_ (_14046_, _14045_, _05549_);
  or _45236_ (_14047_, _14046_, _14042_);
  or _45237_ (_14048_, _14047_, _05535_);
  and _45238_ (_14049_, _14048_, _05542_);
  and _45239_ (_14050_, _14049_, _14038_);
  or _45240_ (_14051_, _14050_, _14028_);
  or _45241_ (_14052_, _14051_, _09850_);
  and _45242_ (_14053_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and _45243_ (_14054_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _45244_ (_14055_, _14054_, _14053_);
  and _45245_ (_14056_, _14055_, _09792_);
  and _45246_ (_14057_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and _45247_ (_14058_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _45248_ (_14059_, _14058_, _14057_);
  and _45249_ (_14060_, _14059_, _05549_);
  or _45250_ (_14061_, _14060_, _14056_);
  or _45251_ (_14062_, _14061_, _09791_);
  and _45252_ (_14063_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and _45253_ (_14064_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _45254_ (_14065_, _14064_, _14063_);
  and _45255_ (_14066_, _14065_, _09792_);
  and _45256_ (_14067_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and _45257_ (_14068_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _45258_ (_14069_, _14068_, _14067_);
  and _45259_ (_14070_, _14069_, _05549_);
  or _45260_ (_14071_, _14070_, _14066_);
  or _45261_ (_14072_, _14071_, _05535_);
  and _45262_ (_14073_, _14072_, _09805_);
  and _45263_ (_14074_, _14073_, _14062_);
  or _45264_ (_14075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _45265_ (_14076_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and _45266_ (_14077_, _14076_, _05549_);
  and _45267_ (_14078_, _14077_, _14075_);
  or _45268_ (_14079_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _45269_ (_14080_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and _45270_ (_14081_, _14080_, _09792_);
  and _45271_ (_14082_, _14081_, _14079_);
  or _45272_ (_14083_, _14082_, _14078_);
  or _45273_ (_14084_, _14083_, _09791_);
  or _45274_ (_14085_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _45275_ (_14086_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and _45276_ (_14087_, _14086_, _05549_);
  and _45277_ (_14088_, _14087_, _14085_);
  or _45278_ (_14089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _45279_ (_14090_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and _45280_ (_14091_, _14090_, _09792_);
  and _45281_ (_14092_, _14091_, _14089_);
  or _45282_ (_14093_, _14092_, _14088_);
  or _45283_ (_14094_, _14093_, _05535_);
  and _45284_ (_14095_, _14094_, _05542_);
  and _45285_ (_14096_, _14095_, _14084_);
  or _45286_ (_14097_, _14096_, _14074_);
  or _45287_ (_14098_, _14097_, _05518_);
  and _45288_ (_14099_, _14098_, _09790_);
  and _45289_ (_14100_, _14099_, _14052_);
  and _45290_ (_14101_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _45291_ (_14102_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or _45292_ (_14103_, _14102_, _14101_);
  and _45293_ (_14104_, _14103_, _09792_);
  and _45294_ (_14105_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _45295_ (_14106_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _45296_ (_14107_, _14106_, _14105_);
  and _45297_ (_14108_, _14107_, _05549_);
  or _45298_ (_14109_, _14108_, _14104_);
  and _45299_ (_14110_, _14109_, _05535_);
  and _45300_ (_14111_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _45301_ (_14112_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _45302_ (_14113_, _14112_, _14111_);
  and _45303_ (_14114_, _14113_, _09792_);
  and _45304_ (_14115_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and _45305_ (_14116_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _45306_ (_14117_, _14116_, _14115_);
  and _45307_ (_14118_, _14117_, _05549_);
  or _45308_ (_14119_, _14118_, _14114_);
  and _45309_ (_14120_, _14119_, _09791_);
  or _45310_ (_14121_, _14120_, _05542_);
  or _45311_ (_14122_, _14121_, _14110_);
  or _45312_ (_14123_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _45313_ (_14124_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and _45314_ (_14125_, _14124_, _05549_);
  and _45315_ (_14126_, _14125_, _14123_);
  or _45316_ (_14127_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _45317_ (_14128_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _45318_ (_14129_, _14128_, _09792_);
  and _45319_ (_14130_, _14129_, _14127_);
  or _45320_ (_14131_, _14130_, _14126_);
  and _45321_ (_14132_, _14131_, _05535_);
  or _45322_ (_14133_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _45323_ (_14134_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _45324_ (_14135_, _14134_, _05549_);
  and _45325_ (_14136_, _14135_, _14133_);
  or _45326_ (_14137_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _45327_ (_14138_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _45328_ (_14139_, _14138_, _09792_);
  and _45329_ (_14140_, _14139_, _14137_);
  or _45330_ (_14141_, _14140_, _14136_);
  and _45331_ (_14142_, _14141_, _09791_);
  or _45332_ (_14143_, _14142_, _09805_);
  or _45333_ (_14144_, _14143_, _14132_);
  and _45334_ (_14145_, _14144_, _14122_);
  or _45335_ (_14146_, _14145_, _05518_);
  and _45336_ (_14147_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and _45337_ (_14148_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _45338_ (_14149_, _14148_, _14147_);
  and _45339_ (_14150_, _14149_, _09792_);
  and _45340_ (_14151_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and _45341_ (_14152_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _45342_ (_14153_, _14152_, _14151_);
  and _45343_ (_14154_, _14153_, _05549_);
  or _45344_ (_14155_, _14154_, _14150_);
  and _45345_ (_14156_, _14155_, _05535_);
  and _45346_ (_14157_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and _45347_ (_14158_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _45348_ (_14159_, _14158_, _14157_);
  and _45349_ (_14160_, _14159_, _09792_);
  and _45350_ (_14161_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and _45351_ (_14162_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _45352_ (_14163_, _14162_, _14161_);
  and _45353_ (_14164_, _14163_, _05549_);
  or _45354_ (_14165_, _14164_, _14160_);
  and _45355_ (_14166_, _14165_, _09791_);
  or _45356_ (_14167_, _14166_, _05542_);
  or _45357_ (_14168_, _14167_, _14156_);
  or _45358_ (_14169_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _45359_ (_14170_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and _45360_ (_14171_, _14170_, _14169_);
  and _45361_ (_14172_, _14171_, _09792_);
  or _45362_ (_14173_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _45363_ (_14174_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and _45364_ (_14175_, _14174_, _14173_);
  and _45365_ (_14176_, _14175_, _05549_);
  or _45366_ (_14177_, _14176_, _14172_);
  and _45367_ (_14178_, _14177_, _05535_);
  or _45368_ (_14179_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _45369_ (_14180_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and _45370_ (_14181_, _14180_, _14179_);
  and _45371_ (_14182_, _14181_, _09792_);
  or _45372_ (_14183_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _45373_ (_14184_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and _45374_ (_14185_, _14184_, _14183_);
  and _45375_ (_14186_, _14185_, _05549_);
  or _45376_ (_14187_, _14186_, _14182_);
  and _45377_ (_14188_, _14187_, _09791_);
  or _45378_ (_14189_, _14188_, _09805_);
  or _45379_ (_14190_, _14189_, _14178_);
  and _45380_ (_14191_, _14190_, _14168_);
  or _45381_ (_14192_, _14191_, _09850_);
  and _45382_ (_14193_, _14192_, _05520_);
  and _45383_ (_14194_, _14193_, _14146_);
  or _45384_ (_14195_, _14194_, _14100_);
  or _45385_ (_14196_, _14195_, _05526_);
  and _45386_ (_14197_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and _45387_ (_14198_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or _45388_ (_14199_, _14198_, _14197_);
  and _45389_ (_14200_, _14199_, _09792_);
  and _45390_ (_14201_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and _45391_ (_14202_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or _45392_ (_14203_, _14202_, _14201_);
  and _45393_ (_14204_, _14203_, _05549_);
  or _45394_ (_14205_, _14204_, _14200_);
  and _45395_ (_14206_, _14205_, _05535_);
  and _45396_ (_14207_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and _45397_ (_14208_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or _45398_ (_14209_, _14208_, _14207_);
  and _45399_ (_14210_, _14209_, _09792_);
  and _45400_ (_14211_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  and _45401_ (_14212_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or _45402_ (_14213_, _14212_, _14211_);
  and _45403_ (_14214_, _14213_, _05549_);
  or _45404_ (_14215_, _14214_, _14210_);
  and _45405_ (_14216_, _14215_, _09791_);
  or _45406_ (_14217_, _14216_, _05542_);
  or _45407_ (_14218_, _14217_, _14206_);
  or _45408_ (_14219_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or _45409_ (_14220_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and _45410_ (_14221_, _14220_, _14219_);
  and _45411_ (_14222_, _14221_, _09792_);
  or _45412_ (_14223_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or _45413_ (_14224_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  and _45414_ (_14225_, _14224_, _14223_);
  and _45415_ (_14226_, _14225_, _05549_);
  or _45416_ (_14227_, _14226_, _14222_);
  and _45417_ (_14228_, _14227_, _05535_);
  or _45418_ (_14229_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or _45419_ (_14230_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and _45420_ (_14231_, _14230_, _14229_);
  and _45421_ (_14232_, _14231_, _09792_);
  or _45422_ (_14233_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or _45423_ (_14234_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and _45424_ (_14235_, _14234_, _14233_);
  and _45425_ (_14236_, _14235_, _05549_);
  or _45426_ (_14237_, _14236_, _14232_);
  and _45427_ (_14238_, _14237_, _09791_);
  or _45428_ (_14239_, _14238_, _09805_);
  or _45429_ (_14240_, _14239_, _14228_);
  and _45430_ (_14241_, _14240_, _14218_);
  or _45431_ (_14242_, _14241_, _05518_);
  and _45432_ (_14243_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and _45433_ (_14244_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _45434_ (_14245_, _14244_, _14243_);
  and _45435_ (_14246_, _14245_, _09792_);
  and _45436_ (_14247_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and _45437_ (_14248_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _45438_ (_14249_, _14248_, _14247_);
  and _45439_ (_14250_, _14249_, _05549_);
  or _45440_ (_14251_, _14250_, _14246_);
  and _45441_ (_14252_, _14251_, _05535_);
  and _45442_ (_14253_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and _45443_ (_14254_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _45444_ (_14255_, _14254_, _14253_);
  and _45445_ (_14256_, _14255_, _09792_);
  and _45446_ (_14257_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and _45447_ (_14258_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _45448_ (_14259_, _14258_, _14257_);
  and _45449_ (_14260_, _14259_, _05549_);
  or _45450_ (_14261_, _14260_, _14256_);
  and _45451_ (_14262_, _14261_, _09791_);
  or _45452_ (_14263_, _14262_, _05542_);
  or _45453_ (_14264_, _14263_, _14252_);
  or _45454_ (_14265_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _45455_ (_14266_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and _45456_ (_14267_, _14266_, _14265_);
  and _45457_ (_14269_, _14267_, _09792_);
  or _45458_ (_14270_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _45459_ (_14271_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and _45460_ (_14272_, _14271_, _14270_);
  and _45461_ (_14273_, _14272_, _05549_);
  or _45462_ (_14274_, _14273_, _14269_);
  and _45463_ (_14275_, _14274_, _05535_);
  or _45464_ (_14276_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _45465_ (_14277_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and _45466_ (_14278_, _14277_, _14276_);
  and _45467_ (_14279_, _14278_, _09792_);
  or _45468_ (_14280_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _45469_ (_14281_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and _45470_ (_14282_, _14281_, _14280_);
  and _45471_ (_14283_, _14282_, _05549_);
  or _45472_ (_14284_, _14283_, _14279_);
  and _45473_ (_14285_, _14284_, _09791_);
  or _45474_ (_14286_, _14285_, _09805_);
  or _45475_ (_14287_, _14286_, _14275_);
  and _45476_ (_14288_, _14287_, _14264_);
  or _45477_ (_14289_, _14288_, _09850_);
  and _45478_ (_14290_, _14289_, _05520_);
  and _45479_ (_14291_, _14290_, _14242_);
  and _45480_ (_14292_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and _45481_ (_14293_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _45482_ (_14294_, _14293_, _14292_);
  and _45483_ (_14295_, _14294_, _05549_);
  and _45484_ (_14296_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and _45485_ (_14297_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _45486_ (_14298_, _14297_, _14296_);
  and _45487_ (_14299_, _14298_, _09792_);
  or _45488_ (_14300_, _14299_, _14295_);
  or _45489_ (_14301_, _14300_, _09791_);
  and _45490_ (_14302_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and _45491_ (_14303_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _45492_ (_14304_, _14303_, _14302_);
  and _45493_ (_14305_, _14304_, _05549_);
  and _45494_ (_14306_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and _45495_ (_14307_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _45496_ (_14308_, _14307_, _14306_);
  and _45497_ (_14309_, _14308_, _09792_);
  or _45498_ (_14310_, _14309_, _14305_);
  or _45499_ (_14311_, _14310_, _05535_);
  and _45500_ (_14312_, _14311_, _09805_);
  and _45501_ (_14313_, _14312_, _14301_);
  or _45502_ (_14314_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _45503_ (_14315_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and _45504_ (_14316_, _14315_, _09792_);
  and _45505_ (_14317_, _14316_, _14314_);
  or _45506_ (_14318_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _45507_ (_14319_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and _45508_ (_14320_, _14319_, _05549_);
  and _45509_ (_14321_, _14320_, _14318_);
  or _45510_ (_14322_, _14321_, _14317_);
  or _45511_ (_14323_, _14322_, _09791_);
  or _45512_ (_14324_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _45513_ (_14325_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and _45514_ (_14326_, _14325_, _09792_);
  and _45515_ (_14327_, _14326_, _14324_);
  or _45516_ (_14328_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _45517_ (_14329_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and _45518_ (_14330_, _14329_, _05549_);
  and _45519_ (_14331_, _14330_, _14328_);
  or _45520_ (_14332_, _14331_, _14327_);
  or _45521_ (_14333_, _14332_, _05535_);
  and _45522_ (_14334_, _14333_, _05542_);
  and _45523_ (_14335_, _14334_, _14323_);
  or _45524_ (_14336_, _14335_, _14313_);
  and _45525_ (_14337_, _14336_, _09850_);
  and _45526_ (_14338_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _45527_ (_14339_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _45528_ (_14340_, _14339_, _09792_);
  or _45529_ (_14341_, _14340_, _14338_);
  and _45530_ (_14342_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and _45531_ (_14343_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _45532_ (_14344_, _14343_, _05549_);
  or _45533_ (_14345_, _14344_, _14342_);
  and _45534_ (_14346_, _14345_, _14341_);
  or _45535_ (_14347_, _14346_, _09791_);
  and _45536_ (_14348_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and _45537_ (_14349_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _45538_ (_14350_, _14349_, _09792_);
  or _45539_ (_14351_, _14350_, _14348_);
  and _45540_ (_14352_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and _45541_ (_14353_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _45542_ (_14354_, _14353_, _05549_);
  or _45543_ (_14355_, _14354_, _14352_);
  and _45544_ (_14356_, _14355_, _14351_);
  or _45545_ (_14357_, _14356_, _05535_);
  and _45546_ (_14358_, _14357_, _09805_);
  and _45547_ (_14359_, _14358_, _14347_);
  or _45548_ (_14360_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _45549_ (_14361_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and _45550_ (_14362_, _14361_, _14360_);
  or _45551_ (_14363_, _14362_, _05549_);
  or _45552_ (_14364_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _45553_ (_14365_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _45554_ (_14366_, _14365_, _14364_);
  or _45555_ (_14367_, _14366_, _09792_);
  and _45556_ (_14368_, _14367_, _14363_);
  or _45557_ (_14369_, _14368_, _09791_);
  or _45558_ (_14370_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _45559_ (_14371_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and _45560_ (_14372_, _14371_, _14370_);
  or _45561_ (_14373_, _14372_, _05549_);
  or _45562_ (_14374_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _45563_ (_14375_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _45564_ (_14376_, _14375_, _14374_);
  or _45565_ (_14377_, _14376_, _09792_);
  and _45566_ (_14378_, _14377_, _14373_);
  or _45567_ (_14379_, _14378_, _05535_);
  and _45568_ (_14380_, _14379_, _05542_);
  and _45569_ (_14381_, _14380_, _14369_);
  or _45570_ (_14382_, _14381_, _14359_);
  and _45571_ (_14383_, _14382_, _05518_);
  or _45572_ (_14384_, _14383_, _14337_);
  and _45573_ (_14385_, _14384_, _09790_);
  or _45574_ (_14386_, _14385_, _14291_);
  or _45575_ (_14387_, _14386_, _10033_);
  and _45576_ (_14388_, _14387_, _14196_);
  or _45577_ (_14389_, _14388_, _00143_);
  and _45578_ (_14390_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and _45579_ (_14391_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _45580_ (_14392_, _14391_, _14390_);
  and _45581_ (_14393_, _14392_, _09792_);
  and _45582_ (_14394_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and _45583_ (_14395_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _45584_ (_14396_, _14395_, _14394_);
  and _45585_ (_14397_, _14396_, _05549_);
  or _45586_ (_14398_, _14397_, _14393_);
  or _45587_ (_14399_, _14398_, _09791_);
  and _45588_ (_14400_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and _45589_ (_14401_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _45590_ (_14402_, _14401_, _14400_);
  and _45591_ (_14403_, _14402_, _09792_);
  and _45592_ (_14404_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and _45593_ (_14405_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _45594_ (_14406_, _14405_, _14404_);
  and _45595_ (_14407_, _14406_, _05549_);
  or _45596_ (_14408_, _14407_, _14403_);
  or _45597_ (_14409_, _14408_, _05535_);
  and _45598_ (_14410_, _14409_, _09805_);
  and _45599_ (_14411_, _14410_, _14399_);
  or _45600_ (_14412_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _45601_ (_14413_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and _45602_ (_14414_, _14413_, _14412_);
  and _45603_ (_14415_, _14414_, _09792_);
  or _45604_ (_14416_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _45605_ (_14417_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and _45606_ (_14418_, _14417_, _14416_);
  and _45607_ (_14419_, _14418_, _05549_);
  or _45608_ (_14420_, _14419_, _14415_);
  or _45609_ (_14421_, _14420_, _09791_);
  or _45610_ (_14422_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _45611_ (_14423_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and _45612_ (_14424_, _14423_, _14422_);
  and _45613_ (_14425_, _14424_, _09792_);
  or _45614_ (_14426_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _45615_ (_14427_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and _45616_ (_14428_, _14427_, _14426_);
  and _45617_ (_14429_, _14428_, _05549_);
  or _45618_ (_14430_, _14429_, _14425_);
  or _45619_ (_14431_, _14430_, _05535_);
  and _45620_ (_14432_, _14431_, _05542_);
  and _45621_ (_14433_, _14432_, _14421_);
  or _45622_ (_14434_, _14433_, _14411_);
  and _45623_ (_14435_, _14434_, _05518_);
  and _45624_ (_14436_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and _45625_ (_14437_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _45626_ (_14438_, _14437_, _14436_);
  and _45627_ (_14439_, _14438_, _09792_);
  and _45628_ (_14440_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _45629_ (_14441_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _45630_ (_14442_, _14441_, _14440_);
  and _45631_ (_14443_, _14442_, _05549_);
  or _45632_ (_14444_, _14443_, _14439_);
  or _45633_ (_14445_, _14444_, _09791_);
  and _45634_ (_14446_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and _45635_ (_14447_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or _45636_ (_14448_, _14447_, _14446_);
  and _45637_ (_14449_, _14448_, _09792_);
  and _45638_ (_14450_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _45639_ (_14451_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _45640_ (_14452_, _14451_, _14450_);
  and _45641_ (_14453_, _14452_, _05549_);
  or _45642_ (_14454_, _14453_, _14449_);
  or _45643_ (_14455_, _14454_, _05535_);
  and _45644_ (_14456_, _14455_, _09805_);
  and _45645_ (_14457_, _14456_, _14445_);
  or _45646_ (_14458_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or _45647_ (_14459_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _45648_ (_14460_, _14459_, _05549_);
  and _45649_ (_14461_, _14460_, _14458_);
  or _45650_ (_14462_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _45651_ (_14463_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _45652_ (_14464_, _14463_, _09792_);
  and _45653_ (_14465_, _14464_, _14462_);
  or _45654_ (_14466_, _14465_, _14461_);
  or _45655_ (_14467_, _14466_, _09791_);
  or _45656_ (_14468_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _45657_ (_14469_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _45658_ (_14470_, _14469_, _05549_);
  and _45659_ (_14471_, _14470_, _14468_);
  or _45660_ (_14472_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or _45661_ (_14473_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and _45662_ (_14474_, _14473_, _09792_);
  and _45663_ (_14475_, _14474_, _14472_);
  or _45664_ (_14476_, _14475_, _14471_);
  or _45665_ (_14477_, _14476_, _05535_);
  and _45666_ (_14478_, _14477_, _05542_);
  and _45667_ (_14479_, _14478_, _14467_);
  or _45668_ (_14480_, _14479_, _14457_);
  and _45669_ (_14481_, _14480_, _09850_);
  or _45670_ (_14482_, _14481_, _14435_);
  and _45671_ (_14483_, _14482_, _09790_);
  and _45672_ (_14484_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and _45673_ (_14485_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or _45674_ (_14486_, _14485_, _14484_);
  and _45675_ (_14487_, _14486_, _09792_);
  and _45676_ (_14488_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and _45677_ (_14489_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or _45678_ (_14490_, _14489_, _14488_);
  and _45679_ (_14491_, _14490_, _05549_);
  or _45680_ (_14492_, _14491_, _14487_);
  and _45681_ (_14493_, _14492_, _05535_);
  and _45682_ (_14494_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and _45683_ (_14495_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or _45684_ (_14496_, _14495_, _14494_);
  and _45685_ (_14497_, _14496_, _09792_);
  and _45686_ (_14498_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _45687_ (_14499_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or _45688_ (_14500_, _14499_, _14498_);
  and _45689_ (_14501_, _14500_, _05549_);
  or _45690_ (_14502_, _14501_, _14497_);
  and _45691_ (_14503_, _14502_, _09791_);
  or _45692_ (_14504_, _14503_, _14493_);
  and _45693_ (_14505_, _14504_, _09805_);
  or _45694_ (_14506_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or _45695_ (_14507_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and _45696_ (_14508_, _14507_, _05549_);
  and _45697_ (_14509_, _14508_, _14506_);
  or _45698_ (_14510_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or _45699_ (_14511_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and _45700_ (_14512_, _14511_, _09792_);
  and _45701_ (_14513_, _14512_, _14510_);
  or _45702_ (_14514_, _14513_, _14509_);
  and _45703_ (_14515_, _14514_, _05535_);
  or _45704_ (_14516_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or _45705_ (_14517_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and _45706_ (_14518_, _14517_, _05549_);
  and _45707_ (_14519_, _14518_, _14516_);
  or _45708_ (_14520_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or _45709_ (_14521_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _45710_ (_14522_, _14521_, _09792_);
  and _45711_ (_14523_, _14522_, _14520_);
  or _45712_ (_14524_, _14523_, _14519_);
  and _45713_ (_14525_, _14524_, _09791_);
  or _45714_ (_14526_, _14525_, _14515_);
  and _45715_ (_14527_, _14526_, _05542_);
  or _45716_ (_14528_, _14527_, _14505_);
  and _45717_ (_14529_, _14528_, _09850_);
  and _45718_ (_14530_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _45719_ (_14531_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _45720_ (_14532_, _14531_, _14530_);
  and _45721_ (_14533_, _14532_, _09792_);
  and _45722_ (_14534_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _45723_ (_14535_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _45724_ (_14536_, _14535_, _14534_);
  and _45725_ (_14537_, _14536_, _05549_);
  or _45726_ (_14538_, _14537_, _14533_);
  and _45727_ (_14539_, _14538_, _05535_);
  and _45728_ (_14540_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and _45729_ (_14541_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _45730_ (_14542_, _14541_, _14540_);
  and _45731_ (_14543_, _14542_, _09792_);
  and _45732_ (_14544_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and _45733_ (_14545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _45734_ (_14546_, _14545_, _14544_);
  and _45735_ (_14547_, _14546_, _05549_);
  or _45736_ (_14548_, _14547_, _14543_);
  and _45737_ (_14549_, _14548_, _09791_);
  or _45738_ (_14550_, _14549_, _14539_);
  and _45739_ (_14551_, _14550_, _09805_);
  or _45740_ (_14552_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _45741_ (_14553_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and _45742_ (_14554_, _14553_, _14552_);
  and _45743_ (_14555_, _14554_, _09792_);
  or _45744_ (_14556_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _45745_ (_14557_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and _45746_ (_14558_, _14557_, _14556_);
  and _45747_ (_14559_, _14558_, _05549_);
  or _45748_ (_14560_, _14559_, _14555_);
  and _45749_ (_14561_, _14560_, _05535_);
  or _45750_ (_14562_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _45751_ (_14563_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and _45752_ (_14564_, _14563_, _14562_);
  and _45753_ (_14565_, _14564_, _09792_);
  or _45754_ (_14566_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _45755_ (_14567_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _45756_ (_14568_, _14567_, _14566_);
  and _45757_ (_14569_, _14568_, _05549_);
  or _45758_ (_14570_, _14569_, _14565_);
  and _45759_ (_14571_, _14570_, _09791_);
  or _45760_ (_14572_, _14571_, _14561_);
  and _45761_ (_14573_, _14572_, _05542_);
  or _45762_ (_14574_, _14573_, _14551_);
  and _45763_ (_14575_, _14574_, _05518_);
  or _45764_ (_14576_, _14575_, _14529_);
  and _45765_ (_14577_, _14576_, _05520_);
  or _45766_ (_14578_, _14577_, _14483_);
  or _45767_ (_14579_, _14578_, _05526_);
  and _45768_ (_14580_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and _45769_ (_14581_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _45770_ (_14582_, _14581_, _14580_);
  and _45771_ (_14583_, _14582_, _09792_);
  and _45772_ (_14584_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and _45773_ (_14585_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _45774_ (_14586_, _14585_, _14584_);
  and _45775_ (_14587_, _14586_, _05549_);
  or _45776_ (_14588_, _14587_, _14583_);
  or _45777_ (_14589_, _14588_, _09791_);
  and _45778_ (_14590_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and _45779_ (_14591_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _45780_ (_14592_, _14591_, _14590_);
  and _45781_ (_14593_, _14592_, _09792_);
  and _45782_ (_14594_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and _45783_ (_14595_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _45784_ (_14596_, _14595_, _14594_);
  and _45785_ (_14597_, _14596_, _05549_);
  or _45786_ (_14598_, _14597_, _14593_);
  or _45787_ (_14599_, _14598_, _05535_);
  and _45788_ (_14600_, _14599_, _09805_);
  and _45789_ (_14601_, _14600_, _14589_);
  or _45790_ (_14602_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _45791_ (_14603_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and _45792_ (_14604_, _14603_, _05549_);
  and _45793_ (_14605_, _14604_, _14602_);
  or _45794_ (_14606_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _45795_ (_14607_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and _45796_ (_14608_, _14607_, _09792_);
  and _45797_ (_14609_, _14608_, _14606_);
  or _45798_ (_14610_, _14609_, _14605_);
  or _45799_ (_14611_, _14610_, _09791_);
  or _45800_ (_14612_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _45801_ (_14613_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and _45802_ (_14614_, _14613_, _05549_);
  and _45803_ (_14615_, _14614_, _14612_);
  or _45804_ (_14616_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _45805_ (_14617_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and _45806_ (_14618_, _14617_, _09792_);
  and _45807_ (_14619_, _14618_, _14616_);
  or _45808_ (_14620_, _14619_, _14615_);
  or _45809_ (_14621_, _14620_, _05535_);
  and _45810_ (_14622_, _14621_, _05542_);
  and _45811_ (_14623_, _14622_, _14611_);
  or _45812_ (_14624_, _14623_, _14601_);
  and _45813_ (_14625_, _14624_, _09850_);
  and _45814_ (_14626_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _45815_ (_14627_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _45816_ (_14628_, _14627_, _14626_);
  and _45817_ (_14629_, _14628_, _09792_);
  and _45818_ (_14630_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _45819_ (_14631_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or _45820_ (_14632_, _14631_, _14630_);
  and _45821_ (_14633_, _14632_, _05549_);
  or _45822_ (_14634_, _14633_, _14629_);
  or _45823_ (_14635_, _14634_, _09791_);
  and _45824_ (_14636_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _45825_ (_14637_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _45826_ (_14638_, _14637_, _14636_);
  and _45827_ (_14639_, _14638_, _09792_);
  and _45828_ (_14640_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _45829_ (_14641_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or _45830_ (_14642_, _14641_, _14640_);
  and _45831_ (_14643_, _14642_, _05549_);
  or _45832_ (_14644_, _14643_, _14639_);
  or _45833_ (_14645_, _14644_, _05535_);
  and _45834_ (_14646_, _14645_, _09805_);
  and _45835_ (_14647_, _14646_, _14635_);
  or _45836_ (_14648_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _45837_ (_14649_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _45838_ (_14650_, _14649_, _14648_);
  and _45839_ (_14651_, _14650_, _09792_);
  or _45840_ (_14652_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _45841_ (_14653_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _45842_ (_14654_, _14653_, _14652_);
  and _45843_ (_14655_, _14654_, _05549_);
  or _45844_ (_14656_, _14655_, _14651_);
  or _45845_ (_14657_, _14656_, _09791_);
  or _45846_ (_14658_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or _45847_ (_14659_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _45848_ (_14660_, _14659_, _14658_);
  and _45849_ (_14661_, _14660_, _09792_);
  or _45850_ (_14662_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _45851_ (_14663_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _45852_ (_14664_, _14663_, _14662_);
  and _45853_ (_14665_, _14664_, _05549_);
  or _45854_ (_14666_, _14665_, _14661_);
  or _45855_ (_14667_, _14666_, _05535_);
  and _45856_ (_14668_, _14667_, _05542_);
  and _45857_ (_14669_, _14668_, _14657_);
  or _45858_ (_14670_, _14669_, _14647_);
  and _45859_ (_14671_, _14670_, _05518_);
  or _45860_ (_14672_, _14671_, _14625_);
  and _45861_ (_14673_, _14672_, _09790_);
  or _45862_ (_14674_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or _45863_ (_14675_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _45864_ (_14676_, _14675_, _14674_);
  and _45865_ (_14677_, _14676_, _09792_);
  or _45866_ (_14678_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or _45867_ (_14679_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _45868_ (_14680_, _14679_, _14678_);
  and _45869_ (_14681_, _14680_, _05549_);
  or _45870_ (_14682_, _14681_, _14677_);
  and _45871_ (_14683_, _14682_, _09791_);
  or _45872_ (_14684_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or _45873_ (_14685_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _45874_ (_14686_, _14685_, _14684_);
  and _45875_ (_14687_, _14686_, _09792_);
  or _45876_ (_14688_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _45877_ (_14689_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and _45878_ (_14690_, _14689_, _14688_);
  and _45879_ (_14691_, _14690_, _05549_);
  or _45880_ (_14692_, _14691_, _14687_);
  and _45881_ (_14693_, _14692_, _05535_);
  or _45882_ (_14694_, _14693_, _14683_);
  and _45883_ (_14695_, _14694_, _05542_);
  and _45884_ (_14696_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _45885_ (_14697_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _45886_ (_14698_, _14697_, _14696_);
  and _45887_ (_14699_, _14698_, _09792_);
  and _45888_ (_14700_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and _45889_ (_14701_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or _45890_ (_14702_, _14701_, _14700_);
  and _45891_ (_14703_, _14702_, _05549_);
  or _45892_ (_14704_, _14703_, _14699_);
  and _45893_ (_14705_, _14704_, _09791_);
  and _45894_ (_14706_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _45895_ (_14707_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _45896_ (_14708_, _14707_, _14706_);
  and _45897_ (_14709_, _14708_, _09792_);
  and _45898_ (_14710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and _45899_ (_14711_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or _45900_ (_14712_, _14711_, _14710_);
  and _45901_ (_14713_, _14712_, _05549_);
  or _45902_ (_14714_, _14713_, _14709_);
  and _45903_ (_14715_, _14714_, _05535_);
  or _45904_ (_14716_, _14715_, _14705_);
  and _45905_ (_14717_, _14716_, _09805_);
  or _45906_ (_14718_, _14717_, _14695_);
  and _45907_ (_14719_, _14718_, _05518_);
  or _45908_ (_14720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _45909_ (_14721_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and _45910_ (_14722_, _14721_, _05549_);
  and _45911_ (_14723_, _14722_, _14720_);
  or _45912_ (_14724_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _45913_ (_14725_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _45914_ (_14726_, _14725_, _09792_);
  and _45915_ (_14727_, _14726_, _14724_);
  or _45916_ (_14728_, _14727_, _14723_);
  and _45917_ (_14729_, _14728_, _09791_);
  or _45918_ (_14730_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _45919_ (_14731_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and _45920_ (_14732_, _14731_, _05549_);
  and _45921_ (_14733_, _14732_, _14730_);
  or _45922_ (_14734_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _45923_ (_14735_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and _45924_ (_14736_, _14735_, _09792_);
  and _45925_ (_14737_, _14736_, _14734_);
  or _45926_ (_14738_, _14737_, _14733_);
  and _45927_ (_14739_, _14738_, _05535_);
  or _45928_ (_14740_, _14739_, _14729_);
  and _45929_ (_14741_, _14740_, _05542_);
  and _45930_ (_14742_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and _45931_ (_14743_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _45932_ (_14744_, _14743_, _14742_);
  and _45933_ (_14745_, _14744_, _09792_);
  and _45934_ (_14746_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _45935_ (_14747_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _45936_ (_14748_, _14747_, _14746_);
  and _45937_ (_14749_, _14748_, _05549_);
  or _45938_ (_14750_, _14749_, _14745_);
  and _45939_ (_14751_, _14750_, _09791_);
  and _45940_ (_14752_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _45941_ (_14753_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _45942_ (_14754_, _14753_, _14752_);
  and _45943_ (_14755_, _14754_, _09792_);
  and _45944_ (_14756_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and _45945_ (_14757_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _45946_ (_14758_, _14757_, _14756_);
  and _45947_ (_14759_, _14758_, _05549_);
  or _45948_ (_14760_, _14759_, _14755_);
  and _45949_ (_14761_, _14760_, _05535_);
  or _45950_ (_14762_, _14761_, _14751_);
  and _45951_ (_14763_, _14762_, _09805_);
  or _45952_ (_14764_, _14763_, _14741_);
  and _45953_ (_14765_, _14764_, _09850_);
  or _45954_ (_14766_, _14765_, _14719_);
  and _45955_ (_14767_, _14766_, _05520_);
  or _45956_ (_14768_, _14767_, _14673_);
  or _45957_ (_14769_, _14768_, _10033_);
  and _45958_ (_14770_, _14769_, _14579_);
  or _45959_ (_14771_, _14770_, _04413_);
  and _45960_ (_14772_, _14771_, _14389_);
  or _45961_ (_14773_, _14772_, _05563_);
  or _45962_ (_14774_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _45963_ (_14775_, _14774_, _22731_);
  and _45964_ (_04746_, _14775_, _14773_);
  and _45965_ (_14776_, _12442_, _24134_);
  and _45966_ (_14777_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  or _45967_ (_04765_, _14777_, _14776_);
  and _45968_ (_14778_, _24476_, _24016_);
  and _45969_ (_14779_, _14778_, _24089_);
  not _45970_ (_14780_, _14778_);
  and _45971_ (_14781_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or _45972_ (_27188_, _14781_, _14779_);
  and _45973_ (_14782_, _14778_, _23583_);
  and _45974_ (_14783_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or _45975_ (_04771_, _14783_, _14782_);
  and _45976_ (_14784_, _08435_, _24134_);
  and _45977_ (_14785_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or _45978_ (_04776_, _14785_, _14784_);
  and _45979_ (_14786_, _14778_, _23887_);
  and _45980_ (_14787_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or _45981_ (_04784_, _14787_, _14786_);
  and _45982_ (_14788_, _14778_, _23548_);
  and _45983_ (_14789_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or _45984_ (_04788_, _14789_, _14788_);
  and _45985_ (_14790_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _45986_ (_14791_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _45987_ (_14792_, _14791_, _14790_);
  and _45988_ (_14793_, _14792_, _09792_);
  and _45989_ (_14794_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and _45990_ (_14795_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _45991_ (_14796_, _14795_, _14794_);
  and _45992_ (_14797_, _14796_, _05549_);
  or _45993_ (_14798_, _14797_, _14793_);
  or _45994_ (_14799_, _14798_, _09791_);
  and _45995_ (_14800_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and _45996_ (_14801_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _45997_ (_14802_, _14801_, _14800_);
  and _45998_ (_14803_, _14802_, _09792_);
  and _45999_ (_14804_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and _46000_ (_14805_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _46001_ (_14806_, _14805_, _14804_);
  and _46002_ (_14807_, _14806_, _05549_);
  or _46003_ (_14808_, _14807_, _14803_);
  or _46004_ (_14809_, _14808_, _05535_);
  and _46005_ (_14810_, _14809_, _09805_);
  and _46006_ (_14811_, _14810_, _14799_);
  or _46007_ (_14812_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _46008_ (_14813_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and _46009_ (_14814_, _14813_, _14812_);
  and _46010_ (_14815_, _14814_, _09792_);
  or _46011_ (_14816_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _46012_ (_14817_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and _46013_ (_14818_, _14817_, _14816_);
  and _46014_ (_14819_, _14818_, _05549_);
  or _46015_ (_14820_, _14819_, _14815_);
  or _46016_ (_14821_, _14820_, _09791_);
  or _46017_ (_14822_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _46018_ (_14823_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and _46019_ (_14824_, _14823_, _14822_);
  and _46020_ (_14825_, _14824_, _09792_);
  or _46021_ (_14826_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _46022_ (_14827_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and _46023_ (_14828_, _14827_, _14826_);
  and _46024_ (_14829_, _14828_, _05549_);
  or _46025_ (_14830_, _14829_, _14825_);
  or _46026_ (_14831_, _14830_, _05535_);
  and _46027_ (_14832_, _14831_, _05542_);
  and _46028_ (_14833_, _14832_, _14821_);
  or _46029_ (_14834_, _14833_, _14811_);
  or _46030_ (_14835_, _14834_, _09850_);
  and _46031_ (_14836_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and _46032_ (_14837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _46033_ (_14838_, _14837_, _14836_);
  and _46034_ (_14839_, _14838_, _09792_);
  and _46035_ (_14840_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and _46036_ (_14841_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _46037_ (_14842_, _14841_, _14840_);
  and _46038_ (_14843_, _14842_, _05549_);
  or _46039_ (_14844_, _14843_, _14839_);
  or _46040_ (_14845_, _14844_, _09791_);
  and _46041_ (_14846_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and _46042_ (_14847_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _46043_ (_14848_, _14847_, _14846_);
  and _46044_ (_14849_, _14848_, _09792_);
  and _46045_ (_14850_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and _46046_ (_14851_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _46047_ (_14852_, _14851_, _14850_);
  and _46048_ (_14853_, _14852_, _05549_);
  or _46049_ (_14854_, _14853_, _14849_);
  or _46050_ (_14855_, _14854_, _05535_);
  and _46051_ (_14856_, _14855_, _09805_);
  and _46052_ (_14857_, _14856_, _14845_);
  or _46053_ (_14858_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _46054_ (_14859_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and _46055_ (_14860_, _14859_, _05549_);
  and _46056_ (_14861_, _14860_, _14858_);
  or _46057_ (_14862_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _46058_ (_14863_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and _46059_ (_14864_, _14863_, _09792_);
  and _46060_ (_14865_, _14864_, _14862_);
  or _46061_ (_14866_, _14865_, _14861_);
  or _46062_ (_14867_, _14866_, _09791_);
  or _46063_ (_14868_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _46064_ (_14869_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and _46065_ (_14870_, _14869_, _05549_);
  and _46066_ (_14871_, _14870_, _14868_);
  or _46067_ (_14872_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _46068_ (_14873_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and _46069_ (_14874_, _14873_, _09792_);
  and _46070_ (_14875_, _14874_, _14872_);
  or _46071_ (_14876_, _14875_, _14871_);
  or _46072_ (_14877_, _14876_, _05535_);
  and _46073_ (_14878_, _14877_, _05542_);
  and _46074_ (_14879_, _14878_, _14867_);
  or _46075_ (_14880_, _14879_, _14857_);
  or _46076_ (_14881_, _14880_, _05518_);
  and _46077_ (_14882_, _14881_, _09790_);
  and _46078_ (_14883_, _14882_, _14835_);
  and _46079_ (_14884_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and _46080_ (_14885_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _46081_ (_14886_, _14885_, _14884_);
  and _46082_ (_14887_, _14886_, _09792_);
  and _46083_ (_14888_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and _46084_ (_14889_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _46085_ (_14890_, _14889_, _14888_);
  and _46086_ (_14891_, _14890_, _05549_);
  or _46087_ (_14892_, _14891_, _14887_);
  and _46088_ (_14893_, _14892_, _05535_);
  and _46089_ (_14894_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and _46090_ (_14895_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _46091_ (_14896_, _14895_, _14894_);
  and _46092_ (_14897_, _14896_, _09792_);
  and _46093_ (_14898_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _46094_ (_14899_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _46095_ (_14900_, _14899_, _14898_);
  and _46096_ (_14901_, _14900_, _05549_);
  or _46097_ (_14902_, _14901_, _14897_);
  and _46098_ (_14903_, _14902_, _09791_);
  or _46099_ (_14904_, _14903_, _05542_);
  or _46100_ (_14905_, _14904_, _14893_);
  or _46101_ (_14906_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _46102_ (_14907_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _46103_ (_14908_, _14907_, _05549_);
  and _46104_ (_14909_, _14908_, _14906_);
  or _46105_ (_14910_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _46106_ (_14911_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _46107_ (_14912_, _14911_, _09792_);
  and _46108_ (_14913_, _14912_, _14910_);
  or _46109_ (_14914_, _14913_, _14909_);
  and _46110_ (_14915_, _14914_, _05535_);
  or _46111_ (_14916_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _46112_ (_14917_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _46113_ (_14918_, _14917_, _05549_);
  and _46114_ (_14919_, _14918_, _14916_);
  or _46115_ (_14920_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _46116_ (_14921_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _46117_ (_14922_, _14921_, _09792_);
  and _46118_ (_14923_, _14922_, _14920_);
  or _46119_ (_14924_, _14923_, _14919_);
  and _46120_ (_14925_, _14924_, _09791_);
  or _46121_ (_14926_, _14925_, _09805_);
  or _46122_ (_14927_, _14926_, _14915_);
  and _46123_ (_14928_, _14927_, _14905_);
  or _46124_ (_14929_, _14928_, _05518_);
  and _46125_ (_14930_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and _46126_ (_14931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _46127_ (_14932_, _14931_, _14930_);
  and _46128_ (_14933_, _14932_, _09792_);
  and _46129_ (_14934_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and _46130_ (_14935_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _46131_ (_14936_, _14935_, _14934_);
  and _46132_ (_14937_, _14936_, _05549_);
  or _46133_ (_14938_, _14937_, _14933_);
  and _46134_ (_14939_, _14938_, _05535_);
  and _46135_ (_14940_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and _46136_ (_14941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _46137_ (_14942_, _14941_, _14940_);
  and _46138_ (_14943_, _14942_, _09792_);
  and _46139_ (_14944_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and _46140_ (_14945_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _46141_ (_14946_, _14945_, _14944_);
  and _46142_ (_14947_, _14946_, _05549_);
  or _46143_ (_14948_, _14947_, _14943_);
  and _46144_ (_14949_, _14948_, _09791_);
  or _46145_ (_14950_, _14949_, _05542_);
  or _46146_ (_14951_, _14950_, _14939_);
  or _46147_ (_14952_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _46148_ (_14953_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and _46149_ (_14954_, _14953_, _14952_);
  and _46150_ (_14955_, _14954_, _09792_);
  or _46151_ (_14956_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _46152_ (_14957_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and _46153_ (_14958_, _14957_, _14956_);
  and _46154_ (_14959_, _14958_, _05549_);
  or _46155_ (_14960_, _14959_, _14955_);
  and _46156_ (_14961_, _14960_, _05535_);
  or _46157_ (_14962_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _46158_ (_14963_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and _46159_ (_14964_, _14963_, _14962_);
  and _46160_ (_14965_, _14964_, _09792_);
  or _46161_ (_14966_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _46162_ (_14967_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and _46163_ (_14968_, _14967_, _14966_);
  and _46164_ (_14969_, _14968_, _05549_);
  or _46165_ (_14970_, _14969_, _14965_);
  and _46166_ (_14971_, _14970_, _09791_);
  or _46167_ (_14972_, _14971_, _09805_);
  or _46168_ (_14973_, _14972_, _14961_);
  and _46169_ (_14974_, _14973_, _14951_);
  or _46170_ (_14975_, _14974_, _09850_);
  and _46171_ (_14976_, _14975_, _05520_);
  and _46172_ (_14977_, _14976_, _14929_);
  or _46173_ (_14978_, _14977_, _14883_);
  or _46174_ (_14979_, _14978_, _05526_);
  and _46175_ (_14980_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and _46176_ (_14981_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or _46177_ (_14982_, _14981_, _14980_);
  and _46178_ (_14983_, _14982_, _09792_);
  and _46179_ (_14984_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and _46180_ (_14985_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or _46181_ (_14986_, _14985_, _14984_);
  and _46182_ (_14987_, _14986_, _05549_);
  or _46183_ (_14988_, _14987_, _14983_);
  and _46184_ (_14989_, _14988_, _05535_);
  and _46185_ (_14990_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and _46186_ (_14991_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or _46187_ (_14992_, _14991_, _14990_);
  and _46188_ (_14993_, _14992_, _09792_);
  and _46189_ (_14994_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and _46190_ (_14995_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or _46191_ (_14996_, _14995_, _14994_);
  and _46192_ (_14997_, _14996_, _05549_);
  or _46193_ (_14998_, _14997_, _14993_);
  and _46194_ (_14999_, _14998_, _09791_);
  or _46195_ (_15000_, _14999_, _05542_);
  or _46196_ (_15001_, _15000_, _14989_);
  or _46197_ (_15002_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or _46198_ (_15003_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  and _46199_ (_15004_, _15003_, _15002_);
  and _46200_ (_15005_, _15004_, _09792_);
  or _46201_ (_15006_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or _46202_ (_15007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and _46203_ (_15008_, _15007_, _15006_);
  and _46204_ (_15009_, _15008_, _05549_);
  or _46205_ (_15010_, _15009_, _15005_);
  and _46206_ (_15011_, _15010_, _05535_);
  or _46207_ (_15012_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or _46208_ (_15013_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  and _46209_ (_15014_, _15013_, _15012_);
  and _46210_ (_15015_, _15014_, _09792_);
  or _46211_ (_15016_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or _46212_ (_15017_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and _46213_ (_15018_, _15017_, _15016_);
  and _46214_ (_15019_, _15018_, _05549_);
  or _46215_ (_15020_, _15019_, _15015_);
  and _46216_ (_15021_, _15020_, _09791_);
  or _46217_ (_15022_, _15021_, _09805_);
  or _46218_ (_15023_, _15022_, _15011_);
  and _46219_ (_15024_, _15023_, _15001_);
  or _46220_ (_15025_, _15024_, _05518_);
  and _46221_ (_15026_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and _46222_ (_15027_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _46223_ (_15028_, _15027_, _15026_);
  and _46224_ (_15029_, _15028_, _09792_);
  and _46225_ (_15030_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and _46226_ (_15031_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _46227_ (_15032_, _15031_, _15030_);
  and _46228_ (_15033_, _15032_, _05549_);
  or _46229_ (_15034_, _15033_, _15029_);
  and _46230_ (_15035_, _15034_, _05535_);
  and _46231_ (_15036_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and _46232_ (_15037_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _46233_ (_15038_, _15037_, _15036_);
  and _46234_ (_15039_, _15038_, _09792_);
  and _46235_ (_15040_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and _46236_ (_15041_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _46237_ (_15042_, _15041_, _15040_);
  and _46238_ (_15043_, _15042_, _05549_);
  or _46239_ (_15044_, _15043_, _15039_);
  and _46240_ (_15045_, _15044_, _09791_);
  or _46241_ (_15046_, _15045_, _05542_);
  or _46242_ (_15047_, _15046_, _15035_);
  or _46243_ (_15048_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _46244_ (_15049_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and _46245_ (_15050_, _15049_, _15048_);
  and _46246_ (_15051_, _15050_, _09792_);
  or _46247_ (_15052_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _46248_ (_15053_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and _46249_ (_15054_, _15053_, _15052_);
  and _46250_ (_15055_, _15054_, _05549_);
  or _46251_ (_15056_, _15055_, _15051_);
  and _46252_ (_15057_, _15056_, _05535_);
  or _46253_ (_15058_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _46254_ (_15059_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and _46255_ (_15060_, _15059_, _15058_);
  and _46256_ (_15061_, _15060_, _09792_);
  or _46257_ (_15062_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _46258_ (_15063_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and _46259_ (_15064_, _15063_, _15062_);
  and _46260_ (_15065_, _15064_, _05549_);
  or _46261_ (_15066_, _15065_, _15061_);
  and _46262_ (_15067_, _15066_, _09791_);
  or _46263_ (_15068_, _15067_, _09805_);
  or _46264_ (_15069_, _15068_, _15057_);
  and _46265_ (_15070_, _15069_, _15047_);
  or _46266_ (_15071_, _15070_, _09850_);
  and _46267_ (_15072_, _15071_, _05520_);
  and _46268_ (_15073_, _15072_, _15025_);
  and _46269_ (_15074_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and _46270_ (_15075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _46271_ (_15076_, _15075_, _15074_);
  and _46272_ (_15077_, _15076_, _05549_);
  and _46273_ (_15078_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and _46274_ (_15079_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _46275_ (_15080_, _15079_, _15078_);
  and _46276_ (_15081_, _15080_, _09792_);
  or _46277_ (_15082_, _15081_, _15077_);
  or _46278_ (_15083_, _15082_, _09791_);
  and _46279_ (_15084_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and _46280_ (_15085_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _46281_ (_15086_, _15085_, _15084_);
  and _46282_ (_15087_, _15086_, _05549_);
  and _46283_ (_15088_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and _46284_ (_15089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _46285_ (_15090_, _15089_, _15088_);
  and _46286_ (_15091_, _15090_, _09792_);
  or _46287_ (_15092_, _15091_, _15087_);
  or _46288_ (_15093_, _15092_, _05535_);
  and _46289_ (_15094_, _15093_, _09805_);
  and _46290_ (_15095_, _15094_, _15083_);
  or _46291_ (_15096_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _46292_ (_15097_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and _46293_ (_15098_, _15097_, _09792_);
  and _46294_ (_15099_, _15098_, _15096_);
  or _46295_ (_15100_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _46296_ (_15101_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and _46297_ (_15102_, _15101_, _05549_);
  and _46298_ (_15103_, _15102_, _15100_);
  or _46299_ (_15104_, _15103_, _15099_);
  or _46300_ (_15105_, _15104_, _09791_);
  or _46301_ (_15106_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _46302_ (_15107_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and _46303_ (_15108_, _15107_, _09792_);
  and _46304_ (_15109_, _15108_, _15106_);
  or _46305_ (_15110_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _46306_ (_15111_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and _46307_ (_15112_, _15111_, _05549_);
  and _46308_ (_15113_, _15112_, _15110_);
  or _46309_ (_15114_, _15113_, _15109_);
  or _46310_ (_15115_, _15114_, _05535_);
  and _46311_ (_15116_, _15115_, _05542_);
  and _46312_ (_15117_, _15116_, _15105_);
  or _46313_ (_15118_, _15117_, _15095_);
  and _46314_ (_15119_, _15118_, _09850_);
  and _46315_ (_15120_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and _46316_ (_15121_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _46317_ (_15122_, _15121_, _09792_);
  or _46318_ (_15123_, _15122_, _15120_);
  and _46319_ (_15124_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _46320_ (_15125_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _46321_ (_15126_, _15125_, _05549_);
  or _46322_ (_15127_, _15126_, _15124_);
  and _46323_ (_15128_, _15127_, _15123_);
  or _46324_ (_15129_, _15128_, _09791_);
  and _46325_ (_15130_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _46326_ (_15131_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _46327_ (_15132_, _15131_, _09792_);
  or _46328_ (_15133_, _15132_, _15130_);
  and _46329_ (_15134_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and _46330_ (_15135_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _46331_ (_15136_, _15135_, _05549_);
  or _46332_ (_15137_, _15136_, _15134_);
  and _46333_ (_15138_, _15137_, _15133_);
  or _46334_ (_15139_, _15138_, _05535_);
  and _46335_ (_15140_, _15139_, _09805_);
  and _46336_ (_15141_, _15140_, _15129_);
  or _46337_ (_15142_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _46338_ (_15143_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _46339_ (_15144_, _15143_, _15142_);
  or _46340_ (_15145_, _15144_, _05549_);
  or _46341_ (_15146_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _46342_ (_15147_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and _46343_ (_15148_, _15147_, _15146_);
  or _46344_ (_15149_, _15148_, _09792_);
  and _46345_ (_15150_, _15149_, _15145_);
  or _46346_ (_15151_, _15150_, _09791_);
  or _46347_ (_15152_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _46348_ (_15153_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and _46349_ (_15154_, _15153_, _15152_);
  or _46350_ (_15155_, _15154_, _05549_);
  or _46351_ (_15156_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _46352_ (_15157_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and _46353_ (_15158_, _15157_, _15156_);
  or _46354_ (_15159_, _15158_, _09792_);
  and _46355_ (_15160_, _15159_, _15155_);
  or _46356_ (_15161_, _15160_, _05535_);
  and _46357_ (_15163_, _15161_, _05542_);
  and _46358_ (_15164_, _15163_, _15151_);
  or _46359_ (_15165_, _15164_, _15141_);
  and _46360_ (_15166_, _15165_, _05518_);
  or _46361_ (_15167_, _15166_, _15119_);
  and _46362_ (_15168_, _15167_, _09790_);
  or _46363_ (_15169_, _15168_, _15073_);
  or _46364_ (_15170_, _15169_, _10033_);
  and _46365_ (_15171_, _15170_, _14979_);
  or _46366_ (_15172_, _15171_, _00143_);
  and _46367_ (_15173_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and _46368_ (_15174_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _46369_ (_15175_, _15174_, _15173_);
  and _46370_ (_15176_, _15175_, _09792_);
  and _46371_ (_15177_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and _46372_ (_15178_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _46373_ (_15179_, _15178_, _15177_);
  and _46374_ (_15180_, _15179_, _05549_);
  or _46375_ (_15181_, _15180_, _15176_);
  or _46376_ (_15182_, _15181_, _09791_);
  and _46377_ (_15183_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and _46378_ (_15184_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _46379_ (_15185_, _15184_, _15183_);
  and _46380_ (_15186_, _15185_, _09792_);
  and _46381_ (_15187_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and _46382_ (_15188_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _46383_ (_15189_, _15188_, _15187_);
  and _46384_ (_15190_, _15189_, _05549_);
  or _46385_ (_15191_, _15190_, _15186_);
  or _46386_ (_15192_, _15191_, _05535_);
  and _46387_ (_15193_, _15192_, _09805_);
  and _46388_ (_15194_, _15193_, _15182_);
  or _46389_ (_15195_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _46390_ (_15196_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and _46391_ (_15197_, _15196_, _15195_);
  and _46392_ (_15198_, _15197_, _09792_);
  or _46393_ (_15199_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _46394_ (_15200_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and _46395_ (_15201_, _15200_, _15199_);
  and _46396_ (_15202_, _15201_, _05549_);
  or _46397_ (_15203_, _15202_, _15198_);
  or _46398_ (_15204_, _15203_, _09791_);
  or _46399_ (_15205_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _46400_ (_15206_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and _46401_ (_15207_, _15206_, _15205_);
  and _46402_ (_15208_, _15207_, _09792_);
  or _46403_ (_15209_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _46404_ (_15210_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and _46405_ (_15211_, _15210_, _15209_);
  and _46406_ (_15212_, _15211_, _05549_);
  or _46407_ (_15214_, _15212_, _15208_);
  or _46408_ (_15215_, _15214_, _05535_);
  and _46409_ (_15216_, _15215_, _05542_);
  and _46410_ (_15217_, _15216_, _15204_);
  or _46411_ (_15218_, _15217_, _15194_);
  and _46412_ (_15219_, _15218_, _05518_);
  and _46413_ (_15220_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _46414_ (_15221_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _46415_ (_15222_, _15221_, _15220_);
  and _46416_ (_15223_, _15222_, _09792_);
  and _46417_ (_15224_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and _46418_ (_15225_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or _46419_ (_15226_, _15225_, _15224_);
  and _46420_ (_15227_, _15226_, _05549_);
  or _46421_ (_15228_, _15227_, _15223_);
  or _46422_ (_15229_, _15228_, _09791_);
  and _46423_ (_15230_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and _46424_ (_15231_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _46425_ (_15232_, _15231_, _15230_);
  and _46426_ (_15233_, _15232_, _09792_);
  and _46427_ (_15235_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _46428_ (_15236_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _46429_ (_15237_, _15236_, _15235_);
  and _46430_ (_15238_, _15237_, _05549_);
  or _46431_ (_15239_, _15238_, _15233_);
  or _46432_ (_15240_, _15239_, _05535_);
  and _46433_ (_15241_, _15240_, _09805_);
  and _46434_ (_15242_, _15241_, _15229_);
  or _46435_ (_15243_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or _46436_ (_15244_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _46437_ (_15245_, _15244_, _05549_);
  and _46438_ (_15246_, _15245_, _15243_);
  or _46439_ (_15247_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _46440_ (_15248_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _46441_ (_15249_, _15248_, _09792_);
  and _46442_ (_15250_, _15249_, _15247_);
  or _46443_ (_15251_, _15250_, _15246_);
  or _46444_ (_15252_, _15251_, _09791_);
  or _46445_ (_15253_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _46446_ (_15254_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and _46447_ (_15255_, _15254_, _05549_);
  and _46448_ (_15256_, _15255_, _15253_);
  or _46449_ (_15257_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or _46450_ (_15258_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _46451_ (_15259_, _15258_, _09792_);
  and _46452_ (_15260_, _15259_, _15257_);
  or _46453_ (_15261_, _15260_, _15256_);
  or _46454_ (_15262_, _15261_, _05535_);
  and _46455_ (_15263_, _15262_, _05542_);
  and _46456_ (_15264_, _15263_, _15252_);
  or _46457_ (_15265_, _15264_, _15242_);
  and _46458_ (_15266_, _15265_, _09850_);
  or _46459_ (_15267_, _15266_, _15219_);
  and _46460_ (_15268_, _15267_, _09790_);
  and _46461_ (_15269_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _46462_ (_15270_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or _46463_ (_15271_, _15270_, _15269_);
  and _46464_ (_15272_, _15271_, _09792_);
  and _46465_ (_15273_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _46466_ (_15274_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _46467_ (_15275_, _15274_, _15273_);
  and _46468_ (_15276_, _15275_, _05549_);
  or _46469_ (_15277_, _15276_, _15272_);
  and _46470_ (_15278_, _15277_, _05535_);
  and _46471_ (_15279_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _46472_ (_15280_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or _46473_ (_15281_, _15280_, _15279_);
  and _46474_ (_15282_, _15281_, _09792_);
  and _46475_ (_15283_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _46476_ (_15284_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _46477_ (_15285_, _15284_, _15283_);
  and _46478_ (_15286_, _15285_, _05549_);
  or _46479_ (_15287_, _15286_, _15282_);
  and _46480_ (_15288_, _15287_, _09791_);
  or _46481_ (_15289_, _15288_, _15278_);
  and _46482_ (_15290_, _15289_, _09805_);
  or _46483_ (_15291_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or _46484_ (_15292_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _46485_ (_15293_, _15292_, _05549_);
  and _46486_ (_15294_, _15293_, _15291_);
  or _46487_ (_15295_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _46488_ (_15296_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _46489_ (_15297_, _15296_, _09792_);
  and _46490_ (_15298_, _15297_, _15295_);
  or _46491_ (_15299_, _15298_, _15294_);
  and _46492_ (_15300_, _15299_, _05535_);
  or _46493_ (_15301_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or _46494_ (_15302_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _46495_ (_15303_, _15302_, _05549_);
  and _46496_ (_15304_, _15303_, _15301_);
  or _46497_ (_15305_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _46498_ (_15306_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and _46499_ (_15307_, _15306_, _09792_);
  and _46500_ (_15308_, _15307_, _15305_);
  or _46501_ (_15309_, _15308_, _15304_);
  and _46502_ (_15310_, _15309_, _09791_);
  or _46503_ (_15311_, _15310_, _15300_);
  and _46504_ (_15312_, _15311_, _05542_);
  or _46505_ (_15313_, _15312_, _15290_);
  and _46506_ (_15314_, _15313_, _09850_);
  and _46507_ (_15315_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and _46508_ (_15316_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _46509_ (_15317_, _15316_, _15315_);
  and _46510_ (_15318_, _15317_, _09792_);
  and _46511_ (_15319_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and _46512_ (_15320_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _46513_ (_15321_, _15320_, _15319_);
  and _46514_ (_15322_, _15321_, _05549_);
  or _46515_ (_15323_, _15322_, _15318_);
  and _46516_ (_15324_, _15323_, _05535_);
  and _46517_ (_15325_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and _46518_ (_15326_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _46519_ (_15327_, _15326_, _15325_);
  and _46520_ (_15328_, _15327_, _09792_);
  and _46521_ (_15329_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and _46522_ (_15330_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _46523_ (_15331_, _15330_, _15329_);
  and _46524_ (_15332_, _15331_, _05549_);
  or _46525_ (_15333_, _15332_, _15328_);
  and _46526_ (_15334_, _15333_, _09791_);
  or _46527_ (_15335_, _15334_, _15324_);
  and _46528_ (_15336_, _15335_, _09805_);
  or _46529_ (_15337_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _46530_ (_15338_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _46531_ (_15339_, _15338_, _15337_);
  and _46532_ (_15340_, _15339_, _09792_);
  or _46533_ (_15341_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _46534_ (_15342_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and _46535_ (_15343_, _15342_, _15341_);
  and _46536_ (_15344_, _15343_, _05549_);
  or _46537_ (_15345_, _15344_, _15340_);
  and _46538_ (_15346_, _15345_, _05535_);
  or _46539_ (_15347_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _46540_ (_15348_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and _46541_ (_15349_, _15348_, _15347_);
  and _46542_ (_15350_, _15349_, _09792_);
  or _46543_ (_15351_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _46544_ (_15352_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and _46545_ (_15353_, _15352_, _15351_);
  and _46546_ (_15354_, _15353_, _05549_);
  or _46547_ (_15355_, _15354_, _15350_);
  and _46548_ (_15356_, _15355_, _09791_);
  or _46549_ (_15357_, _15356_, _15346_);
  and _46550_ (_15358_, _15357_, _05542_);
  or _46551_ (_15359_, _15358_, _15336_);
  and _46552_ (_15360_, _15359_, _05518_);
  or _46553_ (_15361_, _15360_, _15314_);
  and _46554_ (_15362_, _15361_, _05520_);
  or _46555_ (_15363_, _15362_, _15268_);
  or _46556_ (_15364_, _15363_, _05526_);
  and _46557_ (_15365_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and _46558_ (_15366_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _46559_ (_15367_, _15366_, _15365_);
  and _46560_ (_15368_, _15367_, _09792_);
  and _46561_ (_15369_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and _46562_ (_15370_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _46563_ (_15371_, _15370_, _15369_);
  and _46564_ (_15372_, _15371_, _05549_);
  or _46565_ (_15373_, _15372_, _15368_);
  or _46566_ (_15374_, _15373_, _09791_);
  and _46567_ (_15375_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and _46568_ (_15376_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _46569_ (_15377_, _15376_, _15375_);
  and _46570_ (_15378_, _15377_, _09792_);
  and _46571_ (_15379_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and _46572_ (_15380_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _46573_ (_15381_, _15380_, _15379_);
  and _46574_ (_15382_, _15381_, _05549_);
  or _46575_ (_15383_, _15382_, _15378_);
  or _46576_ (_15384_, _15383_, _05535_);
  and _46577_ (_15385_, _15384_, _09805_);
  and _46578_ (_15386_, _15385_, _15374_);
  or _46579_ (_15387_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _46580_ (_15388_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and _46581_ (_15389_, _15388_, _05549_);
  and _46582_ (_15390_, _15389_, _15387_);
  or _46583_ (_15391_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _46584_ (_15392_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and _46585_ (_15393_, _15392_, _09792_);
  and _46586_ (_15394_, _15393_, _15391_);
  or _46587_ (_15395_, _15394_, _15390_);
  or _46588_ (_15396_, _15395_, _09791_);
  or _46589_ (_15397_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _46590_ (_15398_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and _46591_ (_15399_, _15398_, _05549_);
  and _46592_ (_15400_, _15399_, _15397_);
  or _46593_ (_15401_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _46594_ (_15402_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and _46595_ (_15403_, _15402_, _09792_);
  and _46596_ (_15404_, _15403_, _15401_);
  or _46597_ (_15405_, _15404_, _15400_);
  or _46598_ (_15406_, _15405_, _05535_);
  and _46599_ (_15407_, _15406_, _05542_);
  and _46600_ (_15408_, _15407_, _15396_);
  or _46601_ (_15409_, _15408_, _15386_);
  and _46602_ (_15410_, _15409_, _09850_);
  and _46603_ (_15411_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _46604_ (_15412_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _46605_ (_15413_, _15412_, _15411_);
  and _46606_ (_15414_, _15413_, _09792_);
  and _46607_ (_15415_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _46608_ (_15416_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or _46609_ (_15417_, _15416_, _15415_);
  and _46610_ (_15418_, _15417_, _05549_);
  or _46611_ (_15419_, _15418_, _15414_);
  or _46612_ (_15420_, _15419_, _09791_);
  and _46613_ (_15421_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _46614_ (_15422_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or _46615_ (_15423_, _15422_, _15421_);
  and _46616_ (_15424_, _15423_, _09792_);
  and _46617_ (_15425_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _46618_ (_15426_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _46619_ (_15427_, _15426_, _15425_);
  and _46620_ (_15428_, _15427_, _05549_);
  or _46621_ (_15429_, _15428_, _15424_);
  or _46622_ (_15430_, _15429_, _05535_);
  and _46623_ (_15431_, _15430_, _09805_);
  and _46624_ (_15432_, _15431_, _15420_);
  or _46625_ (_15433_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _46626_ (_15434_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _46627_ (_15435_, _15434_, _15433_);
  and _46628_ (_15436_, _15435_, _09792_);
  or _46629_ (_15437_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or _46630_ (_15438_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _46631_ (_15439_, _15438_, _15437_);
  and _46632_ (_15440_, _15439_, _05549_);
  or _46633_ (_15441_, _15440_, _15436_);
  or _46634_ (_15442_, _15441_, _09791_);
  or _46635_ (_15443_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _46636_ (_15444_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _46637_ (_15445_, _15444_, _15443_);
  and _46638_ (_15446_, _15445_, _09792_);
  or _46639_ (_15447_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _46640_ (_15448_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _46641_ (_15449_, _15448_, _15447_);
  and _46642_ (_15450_, _15449_, _05549_);
  or _46643_ (_15451_, _15450_, _15446_);
  or _46644_ (_15452_, _15451_, _05535_);
  and _46645_ (_15453_, _15452_, _05542_);
  and _46646_ (_15454_, _15453_, _15442_);
  or _46647_ (_15455_, _15454_, _15432_);
  and _46648_ (_15456_, _15455_, _05518_);
  or _46649_ (_15457_, _15456_, _15410_);
  and _46650_ (_15458_, _15457_, _09790_);
  or _46651_ (_15459_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or _46652_ (_15460_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and _46653_ (_15461_, _15460_, _15459_);
  and _46654_ (_15462_, _15461_, _09792_);
  or _46655_ (_15463_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _46656_ (_15464_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _46657_ (_15465_, _15464_, _15463_);
  and _46658_ (_15466_, _15465_, _05549_);
  or _46659_ (_15467_, _15466_, _15462_);
  and _46660_ (_15468_, _15467_, _09791_);
  or _46661_ (_15469_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or _46662_ (_15470_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and _46663_ (_15471_, _15470_, _15469_);
  and _46664_ (_15472_, _15471_, _09792_);
  or _46665_ (_15473_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _46666_ (_15474_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _46667_ (_15475_, _15474_, _15473_);
  and _46668_ (_15476_, _15475_, _05549_);
  or _46669_ (_15477_, _15476_, _15472_);
  and _46670_ (_15478_, _15477_, _05535_);
  or _46671_ (_15479_, _15478_, _15468_);
  and _46672_ (_15480_, _15479_, _05542_);
  and _46673_ (_15481_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _46674_ (_15482_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _46675_ (_15483_, _15482_, _15481_);
  and _46676_ (_15484_, _15483_, _09792_);
  and _46677_ (_15485_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _46678_ (_15486_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or _46679_ (_15487_, _15486_, _15485_);
  and _46680_ (_15488_, _15487_, _05549_);
  or _46681_ (_15489_, _15488_, _15484_);
  and _46682_ (_15490_, _15489_, _09791_);
  and _46683_ (_15491_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _46684_ (_15492_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or _46685_ (_15493_, _15492_, _15491_);
  and _46686_ (_15494_, _15493_, _09792_);
  and _46687_ (_15495_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _46688_ (_15496_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _46689_ (_15497_, _15496_, _15495_);
  and _46690_ (_15498_, _15497_, _05549_);
  or _46691_ (_15499_, _15498_, _15494_);
  and _46692_ (_15500_, _15499_, _05535_);
  or _46693_ (_15501_, _15500_, _15490_);
  and _46694_ (_15502_, _15501_, _09805_);
  or _46695_ (_15503_, _15502_, _15480_);
  and _46696_ (_15504_, _15503_, _05518_);
  or _46697_ (_15505_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or _46698_ (_15506_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and _46699_ (_15507_, _15506_, _05549_);
  and _46700_ (_15508_, _15507_, _15505_);
  or _46701_ (_15509_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _46702_ (_15510_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and _46703_ (_15511_, _15510_, _09792_);
  and _46704_ (_15512_, _15511_, _15509_);
  or _46705_ (_15513_, _15512_, _15508_);
  and _46706_ (_15514_, _15513_, _09791_);
  or _46707_ (_15515_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or _46708_ (_15516_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and _46709_ (_15517_, _15516_, _05549_);
  and _46710_ (_15518_, _15517_, _15515_);
  or _46711_ (_15519_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _46712_ (_15520_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and _46713_ (_15521_, _15520_, _09792_);
  and _46714_ (_15522_, _15521_, _15519_);
  or _46715_ (_15523_, _15522_, _15518_);
  and _46716_ (_15524_, _15523_, _05535_);
  or _46717_ (_15525_, _15524_, _15514_);
  and _46718_ (_15526_, _15525_, _05542_);
  and _46719_ (_15527_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and _46720_ (_15528_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _46721_ (_15529_, _15528_, _15527_);
  and _46722_ (_15530_, _15529_, _09792_);
  and _46723_ (_15531_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and _46724_ (_15532_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _46725_ (_15533_, _15532_, _15531_);
  and _46726_ (_15534_, _15533_, _05549_);
  or _46727_ (_15535_, _15534_, _15530_);
  and _46728_ (_15536_, _15535_, _09791_);
  and _46729_ (_15537_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and _46730_ (_15538_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _46731_ (_15539_, _15538_, _15537_);
  and _46732_ (_15540_, _15539_, _09792_);
  and _46733_ (_15541_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and _46734_ (_15542_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or _46735_ (_15543_, _15542_, _15541_);
  and _46736_ (_15544_, _15543_, _05549_);
  or _46737_ (_15545_, _15544_, _15540_);
  and _46738_ (_15546_, _15545_, _05535_);
  or _46739_ (_15547_, _15546_, _15536_);
  and _46740_ (_15548_, _15547_, _09805_);
  or _46741_ (_15549_, _15548_, _15526_);
  and _46742_ (_15550_, _15549_, _09850_);
  or _46743_ (_15551_, _15550_, _15504_);
  and _46744_ (_15552_, _15551_, _05520_);
  or _46745_ (_15553_, _15552_, _15458_);
  or _46746_ (_15554_, _15553_, _10033_);
  and _46747_ (_15555_, _15554_, _15364_);
  or _46748_ (_15556_, _15555_, _04413_);
  and _46749_ (_15557_, _15556_, _15172_);
  or _46750_ (_15558_, _15557_, _05563_);
  or _46751_ (_15559_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _46752_ (_15560_, _15559_, _22731_);
  and _46753_ (_04805_, _15560_, _15558_);
  and _46754_ (_15561_, _24496_, _22974_);
  and _46755_ (_15562_, _15561_, _23996_);
  not _46756_ (_15563_, _15561_);
  and _46757_ (_15564_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _46758_ (_04811_, _15564_, _15562_);
  and _46759_ (_15565_, _24451_, _24089_);
  and _46760_ (_15566_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _46761_ (_04814_, _15566_, _15565_);
  and _46762_ (_15567_, _09779_, _24474_);
  and _46763_ (_15568_, _15567_, _23583_);
  not _46764_ (_15569_, _15567_);
  and _46765_ (_15570_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _46766_ (_04817_, _15570_, _15568_);
  and _46767_ (_15571_, _14778_, _23996_);
  and _46768_ (_15572_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or _46769_ (_04822_, _15572_, _15571_);
  and _46770_ (_15573_, _15567_, _24051_);
  and _46771_ (_15574_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _46772_ (_26992_, _15574_, _15573_);
  and _46773_ (_15575_, _14778_, _24134_);
  and _46774_ (_15576_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or _46775_ (_04834_, _15576_, _15575_);
  and _46776_ (_15577_, _14778_, _24051_);
  and _46777_ (_15578_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or _46778_ (_04836_, _15578_, _15577_);
  and _46779_ (_15579_, _15561_, _24134_);
  and _46780_ (_15580_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _46781_ (_04839_, _15580_, _15579_);
  and _46782_ (_15581_, _24365_, _24159_);
  and _46783_ (_15582_, _15581_, _24051_);
  not _46784_ (_15583_, _15581_);
  and _46785_ (_15584_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or _46786_ (_04842_, _15584_, _15582_);
  and _46787_ (_15585_, _15567_, _24089_);
  and _46788_ (_15586_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _46789_ (_04845_, _15586_, _15585_);
  and _46790_ (_15587_, _08435_, _24051_);
  and _46791_ (_15588_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or _46792_ (_04850_, _15588_, _15587_);
  and _46793_ (_15589_, _14778_, _24219_);
  and _46794_ (_15590_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or _46795_ (_04857_, _15590_, _15589_);
  and _46796_ (_15591_, _03236_, _24051_);
  and _46797_ (_15592_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _46798_ (_04863_, _15592_, _15591_);
  and _46799_ (_15593_, _08523_, _23583_);
  and _46800_ (_15594_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or _46801_ (_04870_, _15594_, _15593_);
  and _46802_ (_15595_, _10746_, _24134_);
  and _46803_ (_15596_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or _46804_ (_04873_, _15596_, _15595_);
  and _46805_ (_15597_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and _46806_ (_15598_, _03221_, _24219_);
  or _46807_ (_04883_, _15598_, _15597_);
  and _46808_ (_15599_, _15561_, _24051_);
  and _46809_ (_15600_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _46810_ (_04889_, _15600_, _15599_);
  and _46811_ (_15601_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and _46812_ (_15602_, _03319_, _24051_);
  or _46813_ (_04906_, _15602_, _15601_);
  and _46814_ (_15603_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  and _46815_ (_15604_, _03221_, _23996_);
  or _46816_ (_27093_, _15604_, _15603_);
  and _46817_ (_15605_, _24899_, _24476_);
  and _46818_ (_15606_, _15605_, _24089_);
  not _46819_ (_15607_, _15605_);
  and _46820_ (_15608_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or _46821_ (_04911_, _15608_, _15606_);
  and _46822_ (_15609_, _10746_, _23996_);
  and _46823_ (_15610_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or _46824_ (_04914_, _15610_, _15609_);
  and _46825_ (_15611_, _15567_, _23996_);
  and _46826_ (_15612_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _46827_ (_04917_, _15612_, _15611_);
  and _46828_ (_15613_, _15605_, _23583_);
  and _46829_ (_15614_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or _46830_ (_04919_, _15614_, _15613_);
  and _46831_ (_15615_, _15605_, _23887_);
  and _46832_ (_15616_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or _46833_ (_04922_, _15616_, _15615_);
  and _46834_ (_15617_, _15567_, _24134_);
  and _46835_ (_15618_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _46836_ (_04927_, _15618_, _15617_);
  and _46837_ (_15620_, _02432_, _23583_);
  and _46838_ (_15621_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  or _46839_ (_04929_, _15621_, _15620_);
  and _46840_ (_15622_, _03370_, _23548_);
  and _46841_ (_15623_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _46842_ (_04931_, _15623_, _15622_);
  and _46843_ (_15624_, _03370_, _23583_);
  and _46844_ (_15625_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _46845_ (_04934_, _15625_, _15624_);
  and _46846_ (_15626_, _04865_, _23548_);
  and _46847_ (_15627_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or _46848_ (_26963_, _15627_, _15626_);
  and _46849_ (_15628_, _15605_, _23996_);
  and _46850_ (_15629_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or _46851_ (_27181_, _15629_, _15628_);
  and _46852_ (_15630_, _03236_, _23583_);
  and _46853_ (_15631_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _46854_ (_04954_, _15631_, _15630_);
  and _46855_ (_15632_, _03236_, _24219_);
  and _46856_ (_15633_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _46857_ (_04958_, _15633_, _15632_);
  and _46858_ (_15634_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  and _46859_ (_15635_, _04614_, _23548_);
  or _46860_ (_04960_, _15635_, _15634_);
  and _46861_ (_15636_, _03236_, _23548_);
  and _46862_ (_15637_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _46863_ (_04962_, _15637_, _15636_);
  and _46864_ (_15638_, _15605_, _24134_);
  and _46865_ (_15639_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or _46866_ (_04963_, _15639_, _15638_);
  and _46867_ (_15640_, _09779_, _24056_);
  and _46868_ (_15641_, _15640_, _23996_);
  not _46869_ (_15642_, _15640_);
  and _46870_ (_15643_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or _46871_ (_04966_, _15643_, _15641_);
  and _46872_ (_15644_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _46873_ (_15645_, _03662_, _24219_);
  or _46874_ (_04968_, _15645_, _15644_);
  and _46875_ (_15646_, _15605_, _24051_);
  and _46876_ (_15647_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or _46877_ (_27180_, _15647_, _15646_);
  and _46878_ (_15648_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  and _46879_ (_15649_, _04614_, _24051_);
  or _46880_ (_04972_, _15649_, _15648_);
  and _46881_ (_15650_, _15640_, _24134_);
  and _46882_ (_15651_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or _46883_ (_26988_, _15651_, _15650_);
  and _46884_ (_15652_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _46885_ (_15653_, _03662_, _23996_);
  or _46886_ (_27096_, _15653_, _15652_);
  and _46887_ (_15654_, _03236_, _23887_);
  and _46888_ (_15655_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _46889_ (_05005_, _15655_, _15654_);
  and _46890_ (_15656_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  not _46891_ (_15657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _46892_ (_15658_, _02248_, _02237_);
  and _46893_ (_15659_, _15658_, _02264_);
  not _46894_ (_15660_, _02237_);
  and _46895_ (_15661_, _02248_, _02236_);
  and _46896_ (_15662_, _15661_, _15660_);
  and _46897_ (_15663_, _15662_, _02272_);
  nor _46898_ (_15664_, _15663_, _15659_);
  nand _46899_ (_15665_, _15664_, _15657_);
  or _46900_ (_15666_, _15664_, _15657_);
  nand _46901_ (_15667_, _15666_, _15665_);
  nor _46902_ (_15668_, _15667_, _02292_);
  and _46903_ (_15669_, _02292_, _23880_);
  or _46904_ (_15670_, _15669_, _15668_);
  and _46905_ (_15671_, _15670_, _02295_);
  or _46906_ (_05019_, _15671_, _15656_);
  and _46907_ (_15672_, _24478_, _24134_);
  and _46908_ (_15673_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _46909_ (_05024_, _15673_, _15672_);
  and _46910_ (_15674_, _08435_, _24089_);
  and _46911_ (_15675_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or _46912_ (_05027_, _15675_, _15674_);
  and _46913_ (_15676_, _24478_, _24051_);
  and _46914_ (_15677_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _46915_ (_05029_, _15677_, _15676_);
  and _46916_ (_15678_, _03370_, _23996_);
  and _46917_ (_15679_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _46918_ (_05052_, _15679_, _15678_);
  and _46919_ (_15680_, _15567_, _23548_);
  and _46920_ (_15681_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _46921_ (_26990_, _15681_, _15680_);
  and _46922_ (_15682_, _15567_, _24219_);
  and _46923_ (_15683_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _46924_ (_26989_, _15683_, _15682_);
  and _46925_ (_15684_, _15605_, _24219_);
  and _46926_ (_15685_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or _46927_ (_05064_, _15685_, _15684_);
  and _46928_ (_15686_, _10746_, _24051_);
  and _46929_ (_15687_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or _46930_ (_05089_, _15687_, _15686_);
  and _46931_ (_15688_, _24320_, _23548_);
  and _46932_ (_15689_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _46933_ (_05091_, _15689_, _15688_);
  and _46934_ (_15690_, _24478_, _23996_);
  and _46935_ (_15691_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _46936_ (_05093_, _15691_, _15690_);
  and _46937_ (_15692_, _10746_, _23583_);
  and _46938_ (_15693_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or _46939_ (_05113_, _15693_, _15692_);
  and _46940_ (_15694_, _24142_, _23583_);
  and _46941_ (_15695_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or _46942_ (_05116_, _15695_, _15694_);
  and _46943_ (_15696_, _07038_, _24051_);
  and _46944_ (_15697_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _46945_ (_05135_, _15697_, _15696_);
  and _46946_ (_15698_, _12429_, _23583_);
  and _46947_ (_15699_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or _46948_ (_05143_, _15699_, _15698_);
  and _46949_ (_15700_, _10746_, _24089_);
  and _46950_ (_15701_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or _46951_ (_27116_, _15701_, _15700_);
  and _46952_ (_15702_, _12429_, _23887_);
  and _46953_ (_15703_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or _46954_ (_27184_, _15703_, _15702_);
  and _46955_ (_15704_, _12429_, _23548_);
  and _46956_ (_15705_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or _46957_ (_27183_, _15705_, _15704_);
  and _46958_ (_15706_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _46959_ (_15707_, _04653_, _23548_);
  or _46960_ (_05154_, _15707_, _15706_);
  and _46961_ (_15708_, _24319_, _24141_);
  and _46962_ (_15709_, _15708_, _24051_);
  not _46963_ (_15710_, _15708_);
  and _46964_ (_15711_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _46965_ (_05163_, _15711_, _15709_);
  and _46966_ (_15712_, _15640_, _24219_);
  and _46967_ (_15713_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or _46968_ (_05166_, _15713_, _15712_);
  and _46969_ (_15714_, _03370_, _24089_);
  and _46970_ (_15715_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _46971_ (_05168_, _15715_, _15714_);
  and _46972_ (_15716_, _09779_, _24223_);
  and _46973_ (_15717_, _15716_, _23996_);
  not _46974_ (_15718_, _15716_);
  and _46975_ (_15719_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _46976_ (_05172_, _15719_, _15717_);
  and _46977_ (_15720_, _15708_, _23887_);
  and _46978_ (_15721_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _46979_ (_05175_, _15721_, _15720_);
  and _46980_ (_15722_, _12429_, _24051_);
  and _46981_ (_15723_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or _46982_ (_05187_, _15723_, _15722_);
  and _46983_ (_15724_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _46984_ (_15725_, _09705_, _24051_);
  or _46985_ (_05189_, _15725_, _15724_);
  and _46986_ (_15726_, _12429_, _24089_);
  and _46987_ (_15727_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or _46988_ (_05206_, _15727_, _15726_);
  and _46989_ (_15728_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _46990_ (_15729_, _09705_, _23548_);
  or _46991_ (_27023_, _15729_, _15728_);
  and _46992_ (_15730_, _08523_, _23887_);
  and _46993_ (_15731_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or _46994_ (_05217_, _15731_, _15730_);
  and _46995_ (_15732_, _15640_, _23583_);
  and _46996_ (_15733_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  or _46997_ (_05220_, _15733_, _15732_);
  and _46998_ (_15734_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _46999_ (_15735_, _09676_, _24134_);
  or _47000_ (_05222_, _15735_, _15734_);
  and _47001_ (_15736_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _47002_ (_15737_, _09676_, _24219_);
  or _47003_ (_05238_, _15737_, _15736_);
  and _47004_ (_15738_, _15640_, _23887_);
  and _47005_ (_15739_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or _47006_ (_05241_, _15739_, _15738_);
  and _47007_ (_15740_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and _47008_ (_15741_, _09645_, _24051_);
  or _47009_ (_05245_, _15741_, _15740_);
  and _47010_ (_15742_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and _47011_ (_15743_, _09645_, _23548_);
  or _47012_ (_05252_, _15743_, _15742_);
  and _47013_ (_15744_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and _47014_ (_15745_, _08591_, _24134_);
  or _47015_ (_05272_, _15745_, _15744_);
  and _47016_ (_15746_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and _47017_ (_15747_, _08591_, _23583_);
  or _47018_ (_27017_, _15747_, _15746_);
  and _47019_ (_15748_, _15708_, _23583_);
  and _47020_ (_15749_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _47021_ (_26926_, _15749_, _15748_);
  and _47022_ (_15750_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and _47023_ (_15751_, _06339_, _24089_);
  or _47024_ (_05283_, _15751_, _15750_);
  and _47025_ (_15752_, _24889_, _23548_);
  and _47026_ (_15753_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _47027_ (_05290_, _15753_, _15752_);
  and _47028_ (_15754_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _47029_ (_15755_, _06339_, _23548_);
  or _47030_ (_27014_, _15755_, _15754_);
  and _47031_ (_15756_, _15716_, _23887_);
  and _47032_ (_15757_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _47033_ (_05320_, _15757_, _15756_);
  and _47034_ (_15758_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and _47035_ (_15759_, _05596_, _24134_);
  or _47036_ (_05325_, _15759_, _15758_);
  and _47037_ (_15760_, _07779_, _24089_);
  and _47038_ (_15761_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  or _47039_ (_05330_, _15761_, _15760_);
  and _47040_ (_15762_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  and _47041_ (_15763_, _05596_, _23548_);
  or _47042_ (_05336_, _15763_, _15762_);
  and _47043_ (_15764_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _47044_ (_15765_, _05580_, _23996_);
  or _47045_ (_05346_, _15765_, _15764_);
  and _47046_ (_15766_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _47047_ (_15767_, _05580_, _23887_);
  or _47048_ (_05354_, _15767_, _15766_);
  and _47049_ (_15768_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and _47050_ (_15769_, _05567_, _23996_);
  or _47051_ (_05357_, _15769_, _15768_);
  and _47052_ (_15770_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and _47053_ (_15771_, _05567_, _23887_);
  or _47054_ (_05369_, _15771_, _15770_);
  and _47055_ (_15772_, _15708_, _23996_);
  and _47056_ (_15773_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _47057_ (_05379_, _15773_, _15772_);
  and _47058_ (_15774_, _09774_, _23548_);
  and _47059_ (_15775_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or _47060_ (_05383_, _15775_, _15774_);
  and _47061_ (_15776_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and _47062_ (_15777_, _04937_, _23583_);
  or _47063_ (_05390_, _15777_, _15776_);
  and _47064_ (_15778_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _47065_ (_15779_, _04905_, _24089_);
  or _47066_ (_05423_, _15779_, _15778_);
  and _47067_ (_15780_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _47068_ (_15781_, _04905_, _24219_);
  or _47069_ (_05433_, _15781_, _15780_);
  and _47070_ (_15782_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _47071_ (_15783_, _04897_, _24051_);
  or _47072_ (_05445_, _15783_, _15782_);
  and _47073_ (_15784_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _47074_ (_15785_, _04879_, _24134_);
  or _47075_ (_05447_, _15785_, _15784_);
  and _47076_ (_15786_, _09774_, _24219_);
  and _47077_ (_15787_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or _47078_ (_05450_, _15787_, _15786_);
  and _47079_ (_15788_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and _47080_ (_15789_, _04879_, _23583_);
  or _47081_ (_05452_, _15789_, _15788_);
  and _47082_ (_15790_, _09670_, _23548_);
  and _47083_ (_15791_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or _47084_ (_27203_, _15791_, _15790_);
  and _47085_ (_15792_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _47086_ (_15793_, _05580_, _24219_);
  or _47087_ (_27013_, _15793_, _15792_);
  nand _47088_ (_15794_, _25025_, _24004_);
  or _47089_ (_15795_, _15794_, _00883_);
  nand _47090_ (_15796_, _15794_, _04308_);
  and _47091_ (_15797_, _15796_, _24179_);
  and _47092_ (_15798_, _15797_, _15795_);
  nor _47093_ (_15799_, _24178_, _04308_);
  and _47094_ (_15800_, _00327_, _25017_);
  and _47095_ (_15801_, _15800_, _25481_);
  nand _47096_ (_15802_, _15801_, _23504_);
  or _47097_ (_15803_, _15801_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _47098_ (_15804_, _15803_, _24539_);
  and _47099_ (_15805_, _15804_, _15802_);
  or _47100_ (_15806_, _15805_, _15799_);
  or _47101_ (_15807_, _15806_, _15798_);
  and _47102_ (_05463_, _15807_, _22731_);
  and _47103_ (_15808_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and _47104_ (_15809_, _02836_, _24219_);
  or _47105_ (_05466_, _15809_, _15808_);
  and _47106_ (_15810_, _07038_, _24089_);
  and _47107_ (_15811_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _47108_ (_05470_, _15811_, _15810_);
  and _47109_ (_15812_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _47110_ (_15813_, _09676_, _23887_);
  or _47111_ (_05474_, _15813_, _15812_);
  and _47112_ (_15814_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not _47113_ (_15815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _47114_ (_15816_, _11153_, _15815_);
  and _47115_ (_15817_, _11153_, _15815_);
  nor _47116_ (_15818_, _15817_, _15816_);
  nor _47117_ (_15819_, _15818_, _02292_);
  and _47118_ (_15820_, _02292_, _02728_);
  or _47119_ (_15821_, _15820_, _15819_);
  and _47120_ (_15822_, _15821_, _02295_);
  or _47121_ (_05476_, _15822_, _15814_);
  or _47122_ (_15823_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _47123_ (_15824_, _15823_, _22731_);
  or _47124_ (_15825_, _11256_, _23577_);
  and _47125_ (_05477_, _15825_, _15824_);
  and _47126_ (_15826_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  and _47127_ (_15827_, _09645_, _23996_);
  or _47128_ (_05483_, _15827_, _15826_);
  and _47129_ (_15828_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and _47130_ (_15829_, _09645_, _23583_);
  or _47131_ (_05503_, _15829_, _15828_);
  and _47132_ (_15830_, _24223_, _24141_);
  and _47133_ (_15831_, _15830_, _24219_);
  not _47134_ (_15832_, _15830_);
  and _47135_ (_15833_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _47136_ (_26928_, _15833_, _15831_);
  and _47137_ (_15834_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and _47138_ (_15835_, _08591_, _24219_);
  or _47139_ (_27016_, _15835_, _15834_);
  and _47140_ (_15836_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  and _47141_ (_15837_, _05596_, _23583_);
  or _47142_ (_05557_, _15837_, _15836_);
  and _47143_ (_15838_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _47144_ (_15839_, _05580_, _24089_);
  or _47145_ (_05564_, _15839_, _15838_);
  and _47146_ (_15840_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and _47147_ (_15841_, _05567_, _24089_);
  or _47148_ (_05575_, _15841_, _15840_);
  and _47149_ (_15842_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and _47150_ (_15843_, _05567_, _24219_);
  or _47151_ (_05581_, _15843_, _15842_);
  and _47152_ (_15844_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and _47153_ (_15845_, _04937_, _24051_);
  or _47154_ (_05586_, _15845_, _15844_);
  and _47155_ (_15846_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and _47156_ (_15847_, _04937_, _23548_);
  or _47157_ (_05588_, _15847_, _15846_);
  and _47158_ (_15848_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _47159_ (_15849_, _04905_, _24134_);
  or _47160_ (_05590_, _15849_, _15848_);
  and _47161_ (_15850_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _47162_ (_15851_, _04905_, _23887_);
  or _47163_ (_27011_, _15851_, _15850_);
  and _47164_ (_15852_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _47165_ (_15853_, _04897_, _23996_);
  or _47166_ (_27009_, _15853_, _15852_);
  or _47167_ (_15854_, _11099_, _23880_);
  and _47168_ (_15855_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _47169_ (_15856_, _02256_, _02248_);
  or _47170_ (_15857_, _15856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _47171_ (_15858_, _11102_, _02281_);
  and _47172_ (_15859_, _15858_, _15857_);
  and _47173_ (_15860_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _47174_ (_15861_, _15860_, _15859_);
  nor _47175_ (_15862_, _15861_, _02616_);
  nor _47176_ (_15863_, _15862_, _15855_);
  nand _47177_ (_15864_, _15863_, _11099_);
  and _47178_ (_15865_, _15864_, _22731_);
  and _47179_ (_05602_, _15865_, _15854_);
  and _47180_ (_15866_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and _47181_ (_15867_, _09705_, _23887_);
  or _47182_ (_05607_, _15867_, _15866_);
  and _47183_ (_15868_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  and _47184_ (_15869_, _08591_, _24089_);
  or _47185_ (_05644_, _15869_, _15868_);
  and _47186_ (_15870_, _08435_, _23996_);
  and _47187_ (_15871_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or _47188_ (_05648_, _15871_, _15870_);
  and _47189_ (_15872_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _47190_ (_15873_, _06339_, _24051_);
  or _47191_ (_05650_, _15873_, _15872_);
  and _47192_ (_15874_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _47193_ (_15875_, _11134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47194_ (_15876_, _15856_, _02281_);
  and _47195_ (_15877_, _15876_, _15875_);
  and _47196_ (_15878_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _47197_ (_15879_, _15878_, _15877_);
  nor _47198_ (_15880_, _15879_, _02616_);
  or _47199_ (_15881_, _15880_, _15874_);
  and _47200_ (_15882_, _15881_, _02295_);
  and _47201_ (_15883_, _02440_, _02728_);
  or _47202_ (_05666_, _15883_, _15882_);
  and _47203_ (_15884_, _03355_, _24051_);
  and _47204_ (_15885_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _47205_ (_05676_, _15885_, _15884_);
  and _47206_ (_15886_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _47207_ (_15887_, _04879_, _23996_);
  or _47208_ (_05695_, _15887_, _15886_);
  and _47209_ (_15888_, _24496_, _24095_);
  and _47210_ (_15889_, _15888_, _23996_);
  not _47211_ (_15890_, _15888_);
  and _47212_ (_15891_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _47213_ (_05703_, _15891_, _15889_);
  and _47214_ (_15892_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _47215_ (_15893_, _09676_, _23583_);
  or _47216_ (_05714_, _15893_, _15892_);
  and _47217_ (_15894_, _15716_, _23548_);
  and _47218_ (_15895_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _47219_ (_05718_, _15895_, _15894_);
  and _47220_ (_15896_, _15830_, _23548_);
  and _47221_ (_15897_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _47222_ (_26929_, _15897_, _15896_);
  and _47223_ (_15898_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _47224_ (_15899_, _04879_, _24219_);
  or _47225_ (_05729_, _15899_, _15898_);
  and _47226_ (_15900_, _15716_, _24219_);
  and _47227_ (_15901_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _47228_ (_05740_, _15901_, _15900_);
  and _47229_ (_15902_, _09780_, _24051_);
  and _47230_ (_15903_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _47231_ (_05778_, _15903_, _15902_);
  and _47232_ (_15904_, _10797_, _23548_);
  and _47233_ (_15905_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or _47234_ (_05781_, _15905_, _15904_);
  and _47235_ (_15906_, _15888_, _24134_);
  and _47236_ (_15907_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _47237_ (_05783_, _15907_, _15906_);
  and _47238_ (_15908_, _10906_, _23583_);
  and _47239_ (_15909_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or _47240_ (_05786_, _15909_, _15908_);
  and _47241_ (_15910_, _15716_, _24051_);
  and _47242_ (_15911_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _47243_ (_05788_, _15911_, _15910_);
  and _47244_ (_15912_, _25319_, _24533_);
  nand _47245_ (_15913_, _15912_, _23504_);
  or _47246_ (_15914_, _15912_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _47247_ (_15915_, _15914_, _24539_);
  and _47248_ (_15916_, _15915_, _15913_);
  or _47249_ (_15917_, _25328_, _23577_);
  or _47250_ (_15918_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _47251_ (_15919_, _15918_, _24179_);
  and _47252_ (_15920_, _15919_, _15917_);
  nor _47253_ (_15921_, _24178_, _03939_);
  or _47254_ (_15922_, _15921_, rst);
  or _47255_ (_15923_, _15922_, _15920_);
  or _47256_ (_05791_, _15923_, _15916_);
  and _47257_ (_15924_, _15716_, _24089_);
  and _47258_ (_15925_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _47259_ (_05794_, _15925_, _15924_);
  and _47260_ (_15926_, _12372_, _24134_);
  and _47261_ (_15927_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or _47262_ (_26997_, _15927_, _15926_);
  and _47263_ (_15928_, _12372_, _24219_);
  and _47264_ (_15929_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or _47265_ (_26995_, _15929_, _15928_);
  and _47266_ (_15930_, _25220_, _24636_);
  nand _47267_ (_15931_, _15930_, _23504_);
  or _47268_ (_15932_, _15930_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47269_ (_15933_, _15932_, _24539_);
  and _47270_ (_15934_, _15933_, _15931_);
  nand _47271_ (_15935_, _25228_, _24082_);
  or _47272_ (_15936_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47273_ (_15937_, _15936_, _24179_);
  and _47274_ (_15938_, _15937_, _15935_);
  nor _47275_ (_15939_, _24178_, _03985_);
  or _47276_ (_15940_, _15939_, rst);
  or _47277_ (_15941_, _15940_, _15938_);
  or _47278_ (_05805_, _15941_, _15934_);
  and _47279_ (_15942_, _15640_, _24089_);
  and _47280_ (_15943_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  or _47281_ (_05812_, _15943_, _15942_);
  and _47282_ (_15944_, _25124_, _24594_);
  nand _47283_ (_15945_, _15944_, _23504_);
  or _47284_ (_15946_, _15944_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47285_ (_15947_, _15946_, _24539_);
  and _47286_ (_15948_, _15947_, _15945_);
  nand _47287_ (_15949_, _25130_, _24126_);
  or _47288_ (_15950_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47289_ (_15951_, _15950_, _24179_);
  and _47290_ (_15952_, _15951_, _15949_);
  nor _47291_ (_15953_, _24178_, _04230_);
  or _47292_ (_15954_, _15953_, rst);
  or _47293_ (_15955_, _15954_, _15952_);
  or _47294_ (_05816_, _15955_, _15948_);
  and _47295_ (_15956_, _09779_, _24319_);
  and _47296_ (_15957_, _15956_, _23887_);
  not _47297_ (_15958_, _15956_);
  and _47298_ (_15959_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _47299_ (_05820_, _15959_, _15957_);
  and _47300_ (_15960_, _09779_, _22974_);
  and _47301_ (_15961_, _15960_, _24089_);
  not _47302_ (_15962_, _15960_);
  and _47303_ (_15963_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  or _47304_ (_05825_, _15963_, _15961_);
  and _47305_ (_15964_, _15956_, _24089_);
  and _47306_ (_15965_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _47307_ (_05833_, _15965_, _15964_);
  and _47308_ (_15966_, _15956_, _23583_);
  and _47309_ (_15967_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _47310_ (_05840_, _15967_, _15966_);
  and _47311_ (_15968_, _25018_, _24636_);
  nand _47312_ (_15969_, _15968_, _23504_);
  or _47313_ (_15970_, _15968_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47314_ (_15971_, _15970_, _24539_);
  and _47315_ (_15972_, _15971_, _15969_);
  nand _47316_ (_15973_, _25026_, _24082_);
  or _47317_ (_15974_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47318_ (_15975_, _15974_, _24179_);
  and _47319_ (_15976_, _15975_, _15973_);
  nor _47320_ (_15977_, _24178_, _04134_);
  or _47321_ (_15978_, _15977_, rst);
  or _47322_ (_15979_, _15978_, _15976_);
  or _47323_ (_05843_, _15979_, _15972_);
  and _47324_ (_15980_, _03308_, _24159_);
  and _47325_ (_15981_, _15980_, _23583_);
  not _47326_ (_15982_, _15980_);
  and _47327_ (_15983_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or _47328_ (_26976_, _15983_, _15981_);
  and _47329_ (_15984_, _03308_, _24297_);
  and _47330_ (_15985_, _15984_, _24051_);
  not _47331_ (_15986_, _15984_);
  and _47332_ (_15987_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _47333_ (_26975_, _15987_, _15985_);
  and _47334_ (_15988_, _03308_, _24016_);
  and _47335_ (_15989_, _15988_, _23996_);
  not _47336_ (_15990_, _15988_);
  and _47337_ (_15991_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or _47338_ (_05859_, _15991_, _15989_);
  and _47339_ (_15992_, _03308_, _24236_);
  and _47340_ (_15993_, _15992_, _23887_);
  not _47341_ (_15994_, _15992_);
  and _47342_ (_15995_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or _47343_ (_05866_, _15995_, _15993_);
  and _47344_ (_15996_, _24141_, _24016_);
  and _47345_ (_15997_, _15996_, _24219_);
  not _47346_ (_15998_, _15996_);
  and _47347_ (_15999_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or _47348_ (_05892_, _15999_, _15997_);
  and _47349_ (_16000_, _03308_, _23941_);
  and _47350_ (_16001_, _16000_, _23887_);
  not _47351_ (_16002_, _16000_);
  and _47352_ (_16003_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or _47353_ (_05909_, _16003_, _16001_);
  and _47354_ (_16004_, _03308_, _24474_);
  and _47355_ (_16005_, _16004_, _23996_);
  not _47356_ (_16006_, _16004_);
  and _47357_ (_16007_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or _47358_ (_05913_, _16007_, _16005_);
  and _47359_ (_16008_, _03308_, _24319_);
  and _47360_ (_16009_, _16008_, _24051_);
  not _47361_ (_16010_, _16008_);
  and _47362_ (_16011_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or _47363_ (_05917_, _16011_, _16009_);
  and _47364_ (_16012_, _15956_, _24134_);
  and _47365_ (_16013_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _47366_ (_05928_, _16013_, _16012_);
  and _47367_ (_16014_, _03308_, _24095_);
  and _47368_ (_16015_, _16014_, _23583_);
  not _47369_ (_16016_, _16014_);
  and _47370_ (_16017_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _47371_ (_05932_, _16017_, _16015_);
  and _47372_ (_16018_, _11441_, _23996_);
  and _47373_ (_16019_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or _47374_ (_05935_, _16019_, _16018_);
  and _47375_ (_16020_, _03308_, _24146_);
  and _47376_ (_16021_, _16020_, _24134_);
  not _47377_ (_16022_, _16020_);
  and _47378_ (_16023_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or _47379_ (_26950_, _16023_, _16021_);
  and _47380_ (_16024_, _16020_, _23887_);
  and _47381_ (_16025_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or _47382_ (_05945_, _16025_, _16024_);
  and _47383_ (_16026_, _03308_, _24140_);
  and _47384_ (_16027_, _16026_, _23887_);
  not _47385_ (_16028_, _16026_);
  and _47386_ (_16029_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or _47387_ (_05951_, _16029_, _16027_);
  and _47388_ (_16030_, _03355_, _24134_);
  and _47389_ (_16031_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _47390_ (_05954_, _16031_, _16030_);
  and _47391_ (_16032_, _03355_, _23887_);
  and _47392_ (_16033_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _47393_ (_05960_, _16033_, _16032_);
  and _47394_ (_16034_, _24297_, _24141_);
  and _47395_ (_16035_, _16034_, _24051_);
  not _47396_ (_16036_, _16034_);
  and _47397_ (_16037_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or _47398_ (_05974_, _16037_, _16035_);
  and _47399_ (_16038_, _15830_, _23583_);
  and _47400_ (_16039_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _47401_ (_05978_, _16039_, _16038_);
  and _47402_ (_16040_, _15996_, _23887_);
  and _47403_ (_16041_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or _47404_ (_05981_, _16041_, _16040_);
  and _47405_ (_16042_, _15960_, _23996_);
  and _47406_ (_16043_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or _47407_ (_05998_, _16043_, _16042_);
  and _47408_ (_16044_, _15960_, _24134_);
  and _47409_ (_16045_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  or _47410_ (_06021_, _16045_, _16044_);
  and _47411_ (_16046_, _11046_, _24051_);
  and _47412_ (_16047_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _47413_ (_27000_, _16047_, _16046_);
  and _47414_ (_16048_, _24372_, _24141_);
  and _47415_ (_16049_, _16048_, _24219_);
  not _47416_ (_16050_, _16048_);
  and _47417_ (_16051_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _47418_ (_06045_, _16051_, _16049_);
  and _47419_ (_16052_, _12442_, _23548_);
  and _47420_ (_16053_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  or _47421_ (_26993_, _16053_, _16052_);
  and _47422_ (_16054_, _16048_, _23887_);
  and _47423_ (_16055_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _47424_ (_06054_, _16055_, _16054_);
  and _47425_ (_16056_, _15956_, _23548_);
  and _47426_ (_16057_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _47427_ (_06059_, _16057_, _16056_);
  and _47428_ (_16058_, _16048_, _23583_);
  and _47429_ (_16059_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _47430_ (_06065_, _16059_, _16058_);
  and _47431_ (_16060_, _09779_, _24146_);
  and _47432_ (_16061_, _16060_, _23548_);
  not _47433_ (_16062_, _16060_);
  and _47434_ (_16063_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _47435_ (_06068_, _16063_, _16061_);
  and _47436_ (_16064_, _25658_, _23996_);
  and _47437_ (_16065_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _47438_ (_06071_, _16065_, _16064_);
  and _47439_ (_16066_, _03308_, _22974_);
  and _47440_ (_16067_, _16066_, _23887_);
  not _47441_ (_16068_, _16066_);
  and _47442_ (_16069_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or _47443_ (_06086_, _16069_, _16067_);
  and _47444_ (_16070_, _06208_, _24219_);
  and _47445_ (_16071_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _47446_ (_06088_, _16071_, _16070_);
  and _47447_ (_16072_, _03308_, _24372_);
  and _47448_ (_16073_, _16072_, _23996_);
  not _47449_ (_16074_, _16072_);
  and _47450_ (_16075_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or _47451_ (_26956_, _16075_, _16073_);
  and _47452_ (_16076_, _16026_, _23996_);
  and _47453_ (_16077_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _47454_ (_06095_, _16077_, _16076_);
  and _47455_ (_16078_, _15960_, _23548_);
  and _47456_ (_16079_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or _47457_ (_06107_, _16079_, _16078_);
  and _47458_ (_16080_, _15996_, _24134_);
  and _47459_ (_16081_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or _47460_ (_26947_, _16081_, _16080_);
  and _47461_ (_16082_, _04865_, _24089_);
  and _47462_ (_16083_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or _47463_ (_26965_, _16083_, _16082_);
  and _47464_ (_16084_, _03309_, _24051_);
  and _47465_ (_16085_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  or _47466_ (_06120_, _16085_, _16084_);
  and _47467_ (_16086_, _15960_, _24219_);
  and _47468_ (_16087_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  or _47469_ (_06123_, _16087_, _16086_);
  and _47470_ (_16088_, _12372_, _23996_);
  and _47471_ (_16089_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  or _47472_ (_06147_, _16089_, _16088_);
  and _47473_ (_16090_, _15640_, _24051_);
  and _47474_ (_16091_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  or _47475_ (_06149_, _16091_, _16090_);
  and _47476_ (_16092_, _15960_, _24051_);
  and _47477_ (_16093_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or _47478_ (_06151_, _16093_, _16092_);
  and _47479_ (_16094_, _02438_, _24607_);
  nand _47480_ (_16095_, _16094_, _24043_);
  not _47481_ (_16096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47482_ (_16097_, _15658_, _02265_);
  and _47483_ (_16098_, _15662_, _02273_);
  or _47484_ (_16099_, _16098_, _16097_);
  and _47485_ (_16100_, _16099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _47486_ (_16101_, _16100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _47487_ (_16102_, _16101_, _16096_);
  and _47488_ (_16103_, _16101_, _16096_);
  or _47489_ (_16104_, _16103_, _16102_);
  or _47490_ (_16105_, _16104_, _02616_);
  and _47491_ (_16106_, _16105_, _02295_);
  and _47492_ (_16107_, _16106_, _16095_);
  and _47493_ (_16108_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _47494_ (_06161_, _16108_, _16107_);
  and _47495_ (_16109_, _25414_, _23583_);
  and _47496_ (_16110_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _47497_ (_27159_, _16110_, _16109_);
  and _47498_ (_16111_, _03308_, _24349_);
  and _47499_ (_16112_, _16111_, _24219_);
  not _47500_ (_16113_, _16111_);
  and _47501_ (_16114_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or _47502_ (_06169_, _16114_, _16112_);
  and _47503_ (_16115_, _16008_, _24134_);
  and _47504_ (_16116_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or _47505_ (_06179_, _16116_, _16115_);
  and _47506_ (_16117_, _15960_, _23583_);
  and _47507_ (_16118_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or _47508_ (_26985_, _16118_, _16117_);
  and _47509_ (_16119_, _15960_, _23887_);
  and _47510_ (_16120_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or _47511_ (_26984_, _16120_, _16119_);
  and _47512_ (_16121_, _24319_, _24301_);
  and _47513_ (_16122_, _16121_, _23996_);
  not _47514_ (_16123_, _16121_);
  and _47515_ (_16124_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _47516_ (_06207_, _16124_, _16122_);
  and _47517_ (_16125_, _16004_, _23548_);
  and _47518_ (_16126_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or _47519_ (_06214_, _16126_, _16125_);
  and _47520_ (_16127_, _16004_, _24219_);
  and _47521_ (_16128_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  or _47522_ (_06225_, _16128_, _16127_);
  and _47523_ (_16129_, _03309_, _23548_);
  and _47524_ (_16130_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or _47525_ (_06229_, _16130_, _16129_);
  and _47526_ (_16131_, _03309_, _24089_);
  and _47527_ (_16132_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or _47528_ (_06232_, _16132_, _16131_);
  and _47529_ (_16133_, _24134_, _24017_);
  and _47530_ (_16134_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or _47531_ (_06239_, _16134_, _16133_);
  and _47532_ (_16135_, _03309_, _24134_);
  and _47533_ (_16136_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or _47534_ (_06243_, _16136_, _16135_);
  and _47535_ (_16137_, _09779_, _24095_);
  and _47536_ (_16138_, _16137_, _23583_);
  not _47537_ (_16139_, _16137_);
  and _47538_ (_16140_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  or _47539_ (_26983_, _16140_, _16138_);
  and _47540_ (_16141_, _16137_, _23887_);
  and _47541_ (_16142_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  or _47542_ (_06248_, _16142_, _16141_);
  and _47543_ (_16143_, _04865_, _23583_);
  and _47544_ (_16144_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _47545_ (_26964_, _16144_, _16143_);
  and _47546_ (_16145_, _16137_, _23548_);
  and _47547_ (_16146_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  or _47548_ (_06266_, _16146_, _16145_);
  and _47549_ (_16147_, _06208_, _23548_);
  and _47550_ (_16148_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _47551_ (_06268_, _16148_, _16147_);
  and _47552_ (_16149_, _15996_, _23548_);
  and _47553_ (_16150_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or _47554_ (_06275_, _16150_, _16149_);
  and _47555_ (_16151_, _15996_, _24051_);
  and _47556_ (_16152_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or _47557_ (_06277_, _16152_, _16151_);
  and _47558_ (_16153_, _16137_, _24219_);
  and _47559_ (_16154_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or _47560_ (_06280_, _16154_, _16153_);
  and _47561_ (_16155_, _15996_, _24089_);
  and _47562_ (_16156_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or _47563_ (_06282_, _16156_, _16155_);
  and _47564_ (_16157_, _16034_, _23548_);
  and _47565_ (_16158_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or _47566_ (_06285_, _16158_, _16157_);
  and _47567_ (_16159_, _16034_, _23583_);
  and _47568_ (_16160_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or _47569_ (_06288_, _16160_, _16159_);
  and _47570_ (_16161_, _16026_, _24134_);
  and _47571_ (_16162_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or _47572_ (_06297_, _16162_, _16161_);
  and _47573_ (_16163_, _16020_, _24089_);
  and _47574_ (_16164_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or _47575_ (_06309_, _16164_, _16163_);
  and _47576_ (_16165_, _16072_, _23887_);
  and _47577_ (_16166_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or _47578_ (_26955_, _16166_, _16165_);
  and _47579_ (_16167_, _16137_, _24134_);
  and _47580_ (_16168_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or _47581_ (_06314_, _16168_, _16167_);
  and _47582_ (_16169_, _16137_, _24051_);
  and _47583_ (_16170_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or _47584_ (_06327_, _16170_, _16169_);
  and _47585_ (_16171_, _16137_, _24089_);
  and _47586_ (_16172_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or _47587_ (_06333_, _16172_, _16171_);
  and _47588_ (_16173_, _16014_, _23548_);
  and _47589_ (_16174_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or _47590_ (_06336_, _16174_, _16173_);
  and _47591_ (_16175_, _24302_, _23887_);
  and _47592_ (_16176_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or _47593_ (_06338_, _16176_, _16175_);
  and _47594_ (_16177_, _16066_, _23548_);
  and _47595_ (_16178_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or _47596_ (_06340_, _16178_, _16177_);
  and _47597_ (_16179_, _16066_, _24051_);
  and _47598_ (_16180_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or _47599_ (_06346_, _16180_, _16179_);
  and _47600_ (_16181_, _24219_, _24017_);
  and _47601_ (_16182_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or _47602_ (_06349_, _16182_, _16181_);
  and _47603_ (_16183_, _16008_, _23887_);
  and _47604_ (_16184_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or _47605_ (_06350_, _16184_, _16183_);
  and _47606_ (_16185_, _03308_, _24899_);
  and _47607_ (_16186_, _16185_, _24051_);
  not _47608_ (_16187_, _16185_);
  and _47609_ (_16188_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _47610_ (_06355_, _16188_, _16186_);
  and _47611_ (_16189_, _16000_, _23996_);
  and _47612_ (_16190_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or _47613_ (_06373_, _16190_, _16189_);
  and _47614_ (_16191_, _09779_, _24372_);
  and _47615_ (_16192_, _16191_, _23548_);
  not _47616_ (_16193_, _16191_);
  and _47617_ (_16194_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _47618_ (_06380_, _16194_, _16192_);
  and _47619_ (_16195_, _16111_, _24051_);
  and _47620_ (_16196_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or _47621_ (_06390_, _16196_, _16195_);
  and _47622_ (_16197_, _16111_, _23887_);
  and _47623_ (_16198_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or _47624_ (_26969_, _16198_, _16197_);
  and _47625_ (_16199_, _16191_, _23583_);
  and _47626_ (_16200_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _47627_ (_06396_, _16200_, _16199_);
  and _47628_ (_16201_, _15988_, _24219_);
  and _47629_ (_16202_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or _47630_ (_06401_, _16202_, _16201_);
  and _47631_ (_16203_, _15992_, _24134_);
  and _47632_ (_16204_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or _47633_ (_06403_, _16204_, _16203_);
  and _47634_ (_16205_, _16191_, _23887_);
  and _47635_ (_16206_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _47636_ (_06408_, _16206_, _16205_);
  and _47637_ (_16207_, _16048_, _24089_);
  and _47638_ (_16208_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _47639_ (_06414_, _16208_, _16207_);
  and _47640_ (_16209_, _16048_, _23996_);
  and _47641_ (_16210_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _47642_ (_06416_, _16210_, _16209_);
  and _47643_ (_16211_, _09779_, _24140_);
  and _47644_ (_16212_, _16211_, _23887_);
  not _47645_ (_16213_, _16211_);
  and _47646_ (_16214_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  or _47647_ (_06420_, _16214_, _16212_);
  and _47648_ (_16215_, _15980_, _23996_);
  and _47649_ (_16216_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or _47650_ (_26978_, _16216_, _16215_);
  and _47651_ (_16217_, _16060_, _24219_);
  and _47652_ (_16218_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _47653_ (_06428_, _16218_, _16217_);
  and _47654_ (_16219_, _16191_, _24219_);
  and _47655_ (_16220_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _47656_ (_06434_, _16220_, _16219_);
  and _47657_ (_16221_, _16060_, _24051_);
  and _47658_ (_16222_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _47659_ (_06436_, _16222_, _16221_);
  and _47660_ (_16223_, _16191_, _23996_);
  and _47661_ (_16224_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _47662_ (_06439_, _16224_, _16223_);
  and _47663_ (_16225_, _16191_, _24089_);
  and _47664_ (_16226_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _47665_ (_06444_, _16226_, _16225_);
  and _47666_ (_16227_, _16137_, _23996_);
  and _47667_ (_16228_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  or _47668_ (_06445_, _16228_, _16227_);
  and _47669_ (_16229_, _15956_, _24219_);
  and _47670_ (_16230_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _47671_ (_06457_, _16230_, _16229_);
  and _47672_ (_16231_, _15956_, _23996_);
  and _47673_ (_16232_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _47674_ (_06459_, _16232_, _16231_);
  and _47675_ (_16233_, _15956_, _24051_);
  and _47676_ (_16234_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _47677_ (_06462_, _16234_, _16233_);
  and _47678_ (_16235_, _16191_, _24134_);
  and _47679_ (_16236_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _47680_ (_06465_, _16236_, _16235_);
  and _47681_ (_16237_, _15716_, _24134_);
  and _47682_ (_16238_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _47683_ (_06467_, _16238_, _16237_);
  and _47684_ (_16239_, _15716_, _23583_);
  and _47685_ (_16240_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _47686_ (_26987_, _16240_, _16239_);
  and _47687_ (_16241_, _15640_, _23548_);
  and _47688_ (_16242_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or _47689_ (_06477_, _16242_, _16241_);
  and _47690_ (_16243_, _15567_, _23887_);
  and _47691_ (_16244_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _47692_ (_26991_, _16244_, _16243_);
  and _47693_ (_16245_, _16191_, _24051_);
  and _47694_ (_16246_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _47695_ (_26982_, _16246_, _16245_);
  and _47696_ (_16247_, _12442_, _24219_);
  and _47697_ (_16248_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  or _47698_ (_06485_, _16248_, _16247_);
  or _47699_ (_16249_, _15794_, _26570_);
  not _47700_ (_16250_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _47701_ (_16251_, _15794_, _16250_);
  and _47702_ (_16252_, _16251_, _24179_);
  and _47703_ (_16253_, _16252_, _16249_);
  nor _47704_ (_16254_, _24178_, _16250_);
  or _47705_ (_16255_, _15794_, _24531_);
  and _47706_ (_16256_, _16251_, _24539_);
  and _47707_ (_16257_, _16256_, _16255_);
  or _47708_ (_16258_, _16257_, _16254_);
  or _47709_ (_16259_, _16258_, _16253_);
  and _47710_ (_06501_, _16259_, _22731_);
  or _47711_ (_16260_, _15794_, _00473_);
  not _47712_ (_16261_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _47713_ (_16262_, _15794_, _16261_);
  and _47714_ (_16263_, _16262_, _24179_);
  and _47715_ (_16264_, _16263_, _16260_);
  nor _47716_ (_16265_, _24178_, _16261_);
  and _47717_ (_16266_, _15800_, _24562_);
  nand _47718_ (_16267_, _16266_, _23504_);
  or _47719_ (_16268_, _16266_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _47720_ (_16269_, _16268_, _24539_);
  and _47721_ (_16270_, _16269_, _16267_);
  or _47722_ (_16271_, _16270_, _16265_);
  or _47723_ (_16272_, _16271_, _16264_);
  and _47724_ (_06504_, _16272_, _22731_);
  or _47725_ (_16273_, _15794_, _00393_);
  not _47726_ (_16274_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _47727_ (_16275_, _15794_, _16274_);
  and _47728_ (_16276_, _16275_, _24179_);
  and _47729_ (_16277_, _16276_, _16273_);
  nor _47730_ (_16278_, _24178_, _16274_);
  and _47731_ (_16279_, _15800_, _24177_);
  nand _47732_ (_16280_, _16279_, _23504_);
  or _47733_ (_16281_, _16279_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _47734_ (_16282_, _16281_, _24539_);
  and _47735_ (_16283_, _16282_, _16280_);
  or _47736_ (_16284_, _16283_, _16278_);
  or _47737_ (_16285_, _16284_, _16277_);
  and _47738_ (_06506_, _16285_, _22731_);
  or _47739_ (_16286_, _15794_, _00569_);
  not _47740_ (_16287_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _47741_ (_16288_, _15794_, _16287_);
  and _47742_ (_16289_, _16288_, _24179_);
  and _47743_ (_16290_, _16289_, _16286_);
  nor _47744_ (_16291_, _24178_, _16287_);
  and _47745_ (_16292_, _15800_, _24533_);
  nand _47746_ (_16293_, _16292_, _23504_);
  or _47747_ (_16294_, _16292_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _47748_ (_16295_, _16294_, _24539_);
  and _47749_ (_16296_, _16295_, _16293_);
  or _47750_ (_16297_, _16296_, _16291_);
  or _47751_ (_16298_, _16297_, _16290_);
  and _47752_ (_06511_, _16298_, _22731_);
  or _47753_ (_16299_, _15794_, _00747_);
  nand _47754_ (_16300_, _15794_, _04315_);
  and _47755_ (_16301_, _16300_, _24179_);
  and _47756_ (_16302_, _16301_, _16299_);
  nor _47757_ (_16303_, _24178_, _04315_);
  and _47758_ (_16304_, _15800_, _24607_);
  nand _47759_ (_16305_, _16304_, _23504_);
  or _47760_ (_16306_, _16304_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _47761_ (_16307_, _16306_, _24539_);
  and _47762_ (_16308_, _16307_, _16305_);
  or _47763_ (_16309_, _16308_, _16303_);
  or _47764_ (_16310_, _16309_, _16302_);
  and _47765_ (_06514_, _16310_, _22731_);
  or _47766_ (_16311_, _15794_, _00654_);
  nand _47767_ (_16312_, _15794_, _04325_);
  and _47768_ (_16313_, _16312_, _24179_);
  and _47769_ (_16314_, _16313_, _16311_);
  nor _47770_ (_16315_, _24178_, _04325_);
  and _47771_ (_16316_, _15800_, _24636_);
  nand _47772_ (_16317_, _16316_, _23504_);
  or _47773_ (_16318_, _16316_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _47774_ (_16319_, _16318_, _24539_);
  and _47775_ (_16320_, _16319_, _16317_);
  or _47776_ (_16321_, _16320_, _16315_);
  or _47777_ (_16322_, _16321_, _16314_);
  and _47778_ (_06517_, _16322_, _22731_);
  and _47779_ (_16323_, _11264_, _24051_);
  and _47780_ (_16324_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _47781_ (_06519_, _16324_, _16323_);
  or _47782_ (_16325_, _15794_, _00814_);
  nand _47783_ (_16326_, _15794_, _04329_);
  and _47784_ (_16327_, _16326_, _24179_);
  and _47785_ (_16328_, _16327_, _16325_);
  nor _47786_ (_16329_, _24178_, _04329_);
  and _47787_ (_16330_, _15800_, _24594_);
  nand _47788_ (_16331_, _16330_, _23504_);
  or _47789_ (_16332_, _16330_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _47790_ (_16333_, _16332_, _24539_);
  and _47791_ (_16334_, _16333_, _16331_);
  or _47792_ (_16335_, _16334_, _16329_);
  or _47793_ (_16336_, _16335_, _16328_);
  and _47794_ (_06526_, _16336_, _22731_);
  and _47795_ (_16337_, _11046_, _24089_);
  and _47796_ (_16338_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _47797_ (_06530_, _16338_, _16337_);
  and _47798_ (_16339_, _16060_, _23887_);
  and _47799_ (_16340_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _47800_ (_26980_, _16340_, _16339_);
  and _47801_ (_16341_, _16060_, _24089_);
  and _47802_ (_16342_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _47803_ (_06541_, _16342_, _16341_);
  and _47804_ (_16343_, _16060_, _23583_);
  and _47805_ (_16344_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _47806_ (_06547_, _16344_, _16343_);
  and _47807_ (_16345_, _11311_, _23548_);
  and _47808_ (_16346_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or _47809_ (_06555_, _16346_, _16345_);
  and _47810_ (_16347_, _09780_, _23887_);
  and _47811_ (_16348_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _47812_ (_06558_, _16348_, _16347_);
  and _47813_ (_16349_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and _47814_ (_16350_, _04853_, _23996_);
  or _47815_ (_06564_, _16350_, _16349_);
  and _47816_ (_16351_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and _47817_ (_16352_, _04853_, _24089_);
  or _47818_ (_06569_, _16352_, _16351_);
  and _47819_ (_16353_, _02478_, _23548_);
  and _47820_ (_16354_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or _47821_ (_06574_, _16354_, _16353_);
  and _47822_ (_16355_, _11311_, _23583_);
  and _47823_ (_16356_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or _47824_ (_06604_, _16356_, _16355_);
  and _47825_ (_16357_, _16060_, _24134_);
  and _47826_ (_16358_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _47827_ (_26981_, _16358_, _16357_);
  and _47828_ (_16359_, _09670_, _24051_);
  and _47829_ (_16360_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or _47830_ (_06614_, _16360_, _16359_);
  and _47831_ (_16361_, _02996_, _24134_);
  and _47832_ (_16362_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  or _47833_ (_27211_, _16362_, _16361_);
  and _47834_ (_16363_, _16060_, _23996_);
  and _47835_ (_16364_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _47836_ (_06627_, _16364_, _16363_);
  and _47837_ (_16365_, _16211_, _23583_);
  and _47838_ (_16366_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  or _47839_ (_06667_, _16366_, _16365_);
  and _47840_ (_26864_, _00143_, _22731_);
  and _47841_ (_16367_, _26687_, _22731_);
  and _47842_ (_26889_, _16367_, _26716_);
  and _47843_ (_06681_, _26889_, _26811_);
  nor _47844_ (_06701_, _00104_, rst);
  and _47845_ (_16368_, _16211_, _24089_);
  and _47846_ (_16369_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  or _47847_ (_06707_, _16369_, _16368_);
  nor _47848_ (_26865_[4], _25834_, rst);
  and _47849_ (_26866_[7], _00124_, _22731_);
  and _47850_ (_16370_, _16211_, _24051_);
  and _47851_ (_16371_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or _47852_ (_06744_, _16371_, _16370_);
  and _47853_ (_26887_, _02050_, _22731_);
  and _47854_ (_26880_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _22731_);
  and _47855_ (_16372_, _26880_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _47856_ (_26886_, _16372_, _26887_);
  and _47857_ (_16373_, _16211_, _23996_);
  and _47858_ (_16374_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or _47859_ (_26979_, _16374_, _16373_);
  nor _47860_ (_16375_, _26605_, rst);
  and _47861_ (_26868_, _16375_, _00339_);
  and _47862_ (_26869_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _22731_);
  and _47863_ (_16376_, _16211_, _24134_);
  and _47864_ (_16377_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  or _47865_ (_06760_, _16377_, _16376_);
  and _47866_ (_16378_, _15561_, _24219_);
  and _47867_ (_16379_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _47868_ (_06787_, _16379_, _16378_);
  and _47869_ (_16380_, _02996_, _24051_);
  and _47870_ (_16381_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or _47871_ (_06806_, _16381_, _16380_);
  and _47872_ (_16382_, _00883_, _26605_);
  and _47873_ (_16383_, _03853_, _26574_);
  and _47874_ (_16384_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _47875_ (_16385_, _26606_, _00885_);
  or _47876_ (_16386_, _16385_, _16384_);
  or _47877_ (_16387_, _16386_, _16383_);
  or _47878_ (_16388_, _16387_, _16382_);
  or _47879_ (_16389_, _01362_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _47880_ (_16390_, _01364_, _23057_);
  or _47881_ (_16391_, _16390_, _00892_);
  and _47882_ (_16392_, _16391_, _16389_);
  nand _47883_ (_16393_, _16392_, _23003_);
  or _47884_ (_16394_, _16392_, _23003_);
  and _47885_ (_16395_, _16394_, _16393_);
  and _47886_ (_16396_, _16395_, _26662_);
  or _47887_ (_16397_, _16396_, _16388_);
  nand _47888_ (_16398_, _01306_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _47889_ (_16399_, _01306_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _47890_ (_16400_, _16399_, _26665_);
  nand _47891_ (_16401_, _16400_, _16398_);
  nand _47892_ (_16402_, _16401_, _00339_);
  or _47893_ (_16403_, _16402_, _16397_);
  and _47894_ (_16404_, _01377_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _47895_ (_16405_, _01377_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _47896_ (_16406_, _16405_, _16404_);
  or _47897_ (_16407_, _16406_, _00339_);
  and _47898_ (_16408_, _16407_, _22731_);
  and _47899_ (_26870_[15], _16408_, _16403_);
  and _47900_ (_16409_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _47901_ (_16410_, _01751_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _47902_ (_16411_, _01751_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _47903_ (_16412_, _16411_, _16410_);
  not _47904_ (_16413_, _16412_);
  nor _47905_ (_16414_, _16413_, _01754_);
  and _47906_ (_16415_, _16413_, _01754_);
  or _47907_ (_16416_, _16415_, _16414_);
  or _47908_ (_16417_, _16416_, _24471_);
  or _47909_ (_16418_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _47910_ (_16419_, _16418_, _01554_);
  and _47911_ (_16420_, _16419_, _16417_);
  or _47912_ (_26871_[15], _16420_, _16409_);
  nor _47913_ (_16421_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _47914_ (_26872_, _16421_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _47915_ (_16422_, _15980_, _24089_);
  and _47916_ (_16423_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or _47917_ (_26977_, _16423_, _16422_);
  and _47918_ (_16424_, _15980_, _24134_);
  and _47919_ (_16425_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or _47920_ (_06817_, _16425_, _16424_);
  and _47921_ (_16426_, _15980_, _24051_);
  and _47922_ (_16427_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  or _47923_ (_06823_, _16427_, _16426_);
  and _47924_ (_16428_, _25672_, _24089_);
  and _47925_ (_16429_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _47926_ (_06869_, _16429_, _16428_);
  and _47927_ (_16430_, _16211_, _23548_);
  and _47928_ (_16431_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  or _47929_ (_06881_, _16431_, _16430_);
  and _47930_ (_16432_, _16211_, _24219_);
  and _47931_ (_16433_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or _47932_ (_06886_, _16433_, _16432_);
  and _47933_ (_16434_, _06356_, _24134_);
  and _47934_ (_16435_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _47935_ (_06897_, _16435_, _16434_);
  and _47936_ (_16436_, _07779_, _24219_);
  and _47937_ (_16437_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  or _47938_ (_06923_, _16437_, _16436_);
  and _47939_ (_16438_, _06356_, _24051_);
  and _47940_ (_16439_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _47941_ (_06928_, _16439_, _16438_);
  and _47942_ (_16440_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _47943_ (_16441_, _04897_, _24219_);
  or _47944_ (_06948_, _16441_, _16440_);
  and _47945_ (_16442_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and _47946_ (_16443_, _04897_, _23548_);
  or _47947_ (_06955_, _16443_, _16442_);
  and _47948_ (_16444_, _16034_, _23887_);
  and _47949_ (_16445_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or _47950_ (_26948_, _16445_, _16444_);
  and _47951_ (_16446_, _15984_, _23996_);
  and _47952_ (_16447_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or _47953_ (_06960_, _16447_, _16446_);
  and _47954_ (_16448_, _15984_, _24134_);
  and _47955_ (_16449_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or _47956_ (_06964_, _16449_, _16448_);
  and _47957_ (_26873_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _22731_);
  nand _47958_ (_16450_, _22737_, _01621_);
  nand _47959_ (_16451_, _16450_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _47960_ (_16452_, _16451_, _01773_);
  and _47961_ (_26874_, _16452_, _22731_);
  and _47962_ (_16453_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _22731_);
  and _47963_ (_16454_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _22731_);
  and _47964_ (_16455_, _16454_, _01773_);
  or _47965_ (_26875_[7], _16455_, _16453_);
  nand _47966_ (_06974_, _00166_, _22731_);
  nor _47967_ (_16456_, _25694_, _25454_);
  nand _47968_ (_16457_, _01797_, _01794_);
  and _47969_ (_16458_, _16457_, _22737_);
  and _47970_ (_16459_, _16458_, _23588_);
  nor _47971_ (_16460_, _16458_, _23588_);
  nor _47972_ (_16461_, _16460_, _16459_);
  nor _47973_ (_16462_, _16461_, _16456_);
  and _47974_ (_16463_, _23600_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _47975_ (_16464_, _16463_, _16456_);
  and _47976_ (_16465_, _16464_, _01544_);
  or _47977_ (_16466_, _16465_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _47978_ (_16467_, _16466_, _16462_);
  and _47979_ (_26876_[2], _16467_, _22731_);
  and _47980_ (_16468_, _24236_, _24141_);
  and _47981_ (_16469_, _16468_, _24089_);
  not _47982_ (_16470_, _16468_);
  and _47983_ (_16471_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _47984_ (_06978_, _16471_, _16469_);
  nand _47985_ (_06980_, _00187_, _22731_);
  and _47986_ (_16472_, _16468_, _23887_);
  and _47987_ (_16473_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _47988_ (_06983_, _16473_, _16472_);
  nor _47989_ (_06988_, _26804_, rst);
  nor _47990_ (_06990_, _00014_, rst);
  nand _47991_ (_06992_, _00204_, _22731_);
  and _47992_ (_16474_, _03313_, _24089_);
  and _47993_ (_16475_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or _47994_ (_06994_, _16475_, _16474_);
  nor _47995_ (_06997_, _00084_, rst);
  nor _47996_ (_06999_, _00046_, rst);
  and _47997_ (_16476_, _24349_, _24141_);
  and _47998_ (_16477_, _16476_, _23583_);
  not _47999_ (_16478_, _16476_);
  and _48000_ (_16479_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _48001_ (_07003_, _16479_, _16477_);
  and _48002_ (_16480_, _23890_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or _48003_ (_16481_, _24244_, _23930_);
  or _48004_ (_16482_, _16481_, _24275_);
  or _48005_ (_16483_, _23842_, _23815_);
  or _48006_ (_16484_, _23904_, _23897_);
  or _48007_ (_16485_, _16484_, _16483_);
  or _48008_ (_16486_, _16485_, _16482_);
  or _48009_ (_16487_, _16486_, _23795_);
  or _48010_ (_16488_, _01980_, _23913_);
  or _48011_ (_16489_, _16488_, _09759_);
  or _48012_ (_16490_, _16489_, _23835_);
  or _48013_ (_16491_, _16490_, _11472_);
  or _48014_ (_16492_, _16491_, _16487_);
  and _48015_ (_16493_, _16492_, _24295_);
  or _48016_ (_26851_[1], _16493_, _16480_);
  and _48017_ (_16494_, _24141_, _23941_);
  and _48018_ (_16495_, _16494_, _23996_);
  not _48019_ (_16496_, _16494_);
  and _48020_ (_16497_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or _48021_ (_26937_, _16497_, _16495_);
  and _48022_ (_16498_, _15980_, _24219_);
  and _48023_ (_16499_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  or _48024_ (_07010_, _16499_, _16498_);
  and _48025_ (_16500_, _23720_, _23635_);
  and _48026_ (_16501_, _16500_, _23761_);
  and _48027_ (_16502_, _23699_, _23675_);
  and _48028_ (_16503_, _16502_, _23740_);
  and _48029_ (_16504_, _22738_, _22731_);
  and _48030_ (_16505_, _16504_, _23656_);
  and _48031_ (_16506_, _16505_, _23612_);
  and _48032_ (_16507_, _16506_, _16503_);
  and _48033_ (_26878_, _16507_, _16501_);
  and _48034_ (_16508_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _01836_);
  and _48035_ (_16509_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _48036_ (_16510_, _16509_, _16508_);
  and _48037_ (_26879_[7], _16510_, _22731_);
  and _48038_ (_16511_, _16494_, _23887_);
  and _48039_ (_16512_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or _48040_ (_07033_, _16512_, _16511_);
  and _48041_ (_16513_, _24899_, _24141_);
  and _48042_ (_16514_, _16513_, _23996_);
  not _48043_ (_16515_, _16513_);
  and _48044_ (_16516_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or _48045_ (_07037_, _16516_, _16514_);
  and _48046_ (_16517_, _15980_, _23887_);
  and _48047_ (_16518_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or _48048_ (_07039_, _16518_, _16517_);
  and _48049_ (_16519_, _16513_, _23887_);
  and _48050_ (_16520_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or _48051_ (_07043_, _16520_, _16519_);
  and _48052_ (_16521_, _15980_, _23548_);
  and _48053_ (_16522_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or _48054_ (_07049_, _16522_, _16521_);
  and _48055_ (_16523_, _24141_, _24095_);
  and _48056_ (_16524_, _16523_, _23548_);
  not _48057_ (_16525_, _16523_);
  and _48058_ (_16526_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or _48059_ (_07051_, _16526_, _16524_);
  and _48060_ (_16527_, _16523_, _23583_);
  and _48061_ (_16528_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or _48062_ (_07054_, _16528_, _16527_);
  and _48063_ (_16529_, _24474_, _24141_);
  and _48064_ (_16530_, _16529_, _23583_);
  not _48065_ (_16531_, _16529_);
  and _48066_ (_16532_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _48067_ (_07059_, _16532_, _16530_);
  and _48068_ (_16533_, _16529_, _23548_);
  and _48069_ (_16534_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _48070_ (_07061_, _16534_, _16533_);
  and _48071_ (_16535_, _24141_, _24056_);
  and _48072_ (_16536_, _16535_, _23996_);
  not _48073_ (_16537_, _16535_);
  and _48074_ (_16538_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or _48075_ (_26931_, _16538_, _16536_);
  and _48076_ (_16539_, _16535_, _23583_);
  and _48077_ (_16540_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or _48078_ (_07075_, _16540_, _16539_);
  and _48079_ (_16541_, _24301_, _23941_);
  and _48080_ (_16542_, _16541_, _24051_);
  not _48081_ (_16543_, _16541_);
  and _48082_ (_16544_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or _48083_ (_27225_, _16544_, _16542_);
  and _48084_ (_16545_, _15708_, _24219_);
  and _48085_ (_16546_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _48086_ (_07081_, _16546_, _16545_);
  and _48087_ (_16547_, _06356_, _23548_);
  and _48088_ (_16548_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _48089_ (_07083_, _16548_, _16547_);
  and _48090_ (_16549_, _15984_, _23887_);
  and _48091_ (_16550_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or _48092_ (_07089_, _16550_, _16549_);
  and _48093_ (_16551_, _24141_, _22974_);
  and _48094_ (_16552_, _16551_, _23996_);
  not _48095_ (_16553_, _16551_);
  and _48096_ (_16554_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or _48097_ (_07092_, _16554_, _16552_);
  and _48098_ (_16555_, _16551_, _24051_);
  and _48099_ (_16556_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or _48100_ (_07094_, _16556_, _16555_);
  and _48101_ (_16557_, _11441_, _24134_);
  and _48102_ (_16558_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _48103_ (_07100_, _16558_, _16557_);
  and _48104_ (_16559_, _15561_, _23548_);
  and _48105_ (_16560_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or _48106_ (_07103_, _16560_, _16559_);
  and _48107_ (_16561_, _16523_, _24134_);
  and _48108_ (_16562_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or _48109_ (_07107_, _16562_, _16561_);
  nand _48110_ (_16563_, _01816_, _24043_);
  and _48111_ (_16564_, _08221_, _08217_);
  and _48112_ (_16565_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _48113_ (_16566_, _16565_, _16564_);
  and _48114_ (_16567_, _16566_, _02193_);
  and _48115_ (_16568_, _08221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _48116_ (_16569_, _16568_, _16567_);
  or _48117_ (_16570_, _16569_, _01816_);
  and _48118_ (_16571_, _16570_, _22731_);
  and _48119_ (_07109_, _16571_, _16563_);
  and _48120_ (_16572_, _16523_, _23887_);
  and _48121_ (_16573_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or _48122_ (_26924_, _16573_, _16572_);
  and _48123_ (_16574_, _16523_, _24219_);
  and _48124_ (_16575_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or _48125_ (_07113_, _16575_, _16574_);
  and _48126_ (_16576_, _15984_, _23548_);
  and _48127_ (_16577_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or _48128_ (_07115_, _16577_, _16576_);
  and _48129_ (_16578_, _06356_, _24219_);
  and _48130_ (_16579_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _48131_ (_07117_, _16579_, _16578_);
  and _48132_ (_16580_, _08523_, _24134_);
  and _48133_ (_16581_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or _48134_ (_07123_, _16581_, _16580_);
  and _48135_ (_16582_, _15984_, _24219_);
  and _48136_ (_16583_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _48137_ (_07125_, _16583_, _16582_);
  and _48138_ (_16584_, _16048_, _24051_);
  and _48139_ (_16585_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _48140_ (_07130_, _16585_, _16584_);
  and _48141_ (_16586_, _16048_, _23548_);
  and _48142_ (_16587_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _48143_ (_07141_, _16587_, _16586_);
  and _48144_ (_16588_, _15830_, _23887_);
  and _48145_ (_16589_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _48146_ (_26930_, _16589_, _16588_);
  and _48147_ (_16590_, _16523_, _24051_);
  and _48148_ (_16591_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or _48149_ (_07145_, _16591_, _16590_);
  and _48150_ (_16592_, _15708_, _24089_);
  and _48151_ (_16593_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _48152_ (_07164_, _16593_, _16592_);
  and _48153_ (_16594_, _15708_, _24134_);
  and _48154_ (_16595_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _48155_ (_26927_, _16595_, _16594_);
  not _48156_ (_16596_, _01862_);
  and _48157_ (_16597_, _01865_, _16596_);
  or _48158_ (_16598_, _01867_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _48159_ (_26882_[3], _16598_, _22731_);
  and _48160_ (_16599_, _26882_[3], _01870_);
  and _48161_ (_26881_, _16599_, _16597_);
  and _48162_ (_16600_, _16523_, _23996_);
  and _48163_ (_16601_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or _48164_ (_07177_, _16601_, _16600_);
  and _48165_ (_16602_, _16541_, _24089_);
  and _48166_ (_16603_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or _48167_ (_07180_, _16603_, _16602_);
  and _48168_ (_16604_, _15984_, _24089_);
  and _48169_ (_16605_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or _48170_ (_07185_, _16605_, _16604_);
  and _48171_ (_16606_, _16476_, _24051_);
  and _48172_ (_16607_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _48173_ (_07188_, _16607_, _16606_);
  and _48174_ (_16608_, _16494_, _24089_);
  and _48175_ (_16609_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or _48176_ (_07194_, _16609_, _16608_);
  and _48177_ (_16610_, _16513_, _24089_);
  and _48178_ (_16611_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or _48179_ (_07197_, _16611_, _16610_);
  and _48180_ (_16612_, _16513_, _24219_);
  and _48181_ (_16613_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or _48182_ (_26934_, _16613_, _16612_);
  and _48183_ (_16614_, _16529_, _24051_);
  and _48184_ (_16615_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _48185_ (_07201_, _16615_, _16614_);
  and _48186_ (_16616_, _15984_, _23583_);
  and _48187_ (_16617_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or _48188_ (_07204_, _16617_, _16616_);
  and _48189_ (_16618_, _06356_, _23583_);
  and _48190_ (_16619_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _48191_ (_27178_, _16619_, _16618_);
  and _48192_ (_16620_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _48193_ (_16621_, _01218_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _48194_ (_16622_, _16621_, _16620_);
  and _48195_ (_26883_[31], _16622_, _22731_);
  and _48196_ (_16623_, _07779_, _23887_);
  and _48197_ (_16624_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or _48198_ (_07214_, _16624_, _16623_);
  and _48199_ (_16625_, _16535_, _24219_);
  and _48200_ (_16626_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or _48201_ (_07216_, _16626_, _16625_);
  and _48202_ (_16627_, _16551_, _24219_);
  and _48203_ (_16628_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or _48204_ (_07221_, _16628_, _16627_);
  and _48205_ (_16629_, _24017_, _23887_);
  and _48206_ (_16630_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or _48207_ (_07226_, _16630_, _16629_);
  and _48208_ (_16631_, _16551_, _23887_);
  and _48209_ (_16632_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or _48210_ (_07232_, _16632_, _16631_);
  and _48211_ (_16633_, _16523_, _24089_);
  and _48212_ (_16634_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or _48213_ (_26925_, _16634_, _16633_);
  and _48214_ (_16635_, _15830_, _24089_);
  and _48215_ (_16636_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _48216_ (_07245_, _16636_, _16635_);
  and _48217_ (_16637_, _08523_, _24051_);
  and _48218_ (_16638_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or _48219_ (_27082_, _16638_, _16637_);
  and _48220_ (_16639_, _15988_, _23583_);
  and _48221_ (_16640_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _48222_ (_07251_, _16640_, _16639_);
  and _48223_ (_16641_, _15988_, _23887_);
  and _48224_ (_16642_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or _48225_ (_07266_, _16642_, _16641_);
  and _48226_ (_16643_, _15988_, _23548_);
  and _48227_ (_16644_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or _48228_ (_07270_, _16644_, _16643_);
  or _48229_ (_16645_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _48230_ (_16646_, _25694_, _25457_);
  and _48231_ (_16647_, _16646_, _22731_);
  and _48232_ (_26884_[31], _16647_, _16645_);
  and _48233_ (_16648_, _16551_, _23548_);
  and _48234_ (_16649_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or _48235_ (_07293_, _16649_, _16648_);
  and _48236_ (_16650_, _16535_, _24089_);
  and _48237_ (_16651_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or _48238_ (_07297_, _16651_, _16650_);
  and _48239_ (_16652_, _15708_, _23548_);
  and _48240_ (_16653_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _48241_ (_07300_, _16653_, _16652_);
  and _48242_ (_16654_, _03241_, _23996_);
  and _48243_ (_16655_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or _48244_ (_07306_, _16655_, _16654_);
  and _48245_ (_16656_, _16048_, _24134_);
  and _48246_ (_16657_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _48247_ (_07309_, _16657_, _16656_);
  and _48248_ (_16658_, _03241_, _24134_);
  and _48249_ (_16659_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  or _48250_ (_27173_, _16659_, _16658_);
  and _48251_ (_16660_, _16494_, _24219_);
  and _48252_ (_16661_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or _48253_ (_07317_, _16661_, _16660_);
  and _48254_ (_16662_, _15830_, _24051_);
  and _48255_ (_16663_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _48256_ (_07324_, _16663_, _16662_);
  and _48257_ (_16664_, _15988_, _24134_);
  and _48258_ (_16665_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or _48259_ (_26974_, _16665_, _16664_);
  and _48260_ (_16666_, _24394_, _23548_);
  and _48261_ (_16667_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _48262_ (_07338_, _16667_, _16666_);
  and _48263_ (_16668_, _15988_, _24051_);
  and _48264_ (_16669_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or _48265_ (_07341_, _16669_, _16668_);
  and _48266_ (_16670_, _24496_, _24159_);
  and _48267_ (_16671_, _16670_, _24134_);
  not _48268_ (_16672_, _16670_);
  and _48269_ (_16673_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or _48270_ (_07344_, _16673_, _16671_);
  and _48271_ (_16674_, _16670_, _24219_);
  and _48272_ (_16675_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or _48273_ (_07346_, _16675_, _16674_);
  and _48274_ (_16676_, _15988_, _24089_);
  and _48275_ (_16677_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or _48276_ (_07349_, _16677_, _16676_);
  and _48277_ (_16678_, _24496_, _24297_);
  and _48278_ (_16679_, _16678_, _23887_);
  not _48279_ (_16680_, _16678_);
  and _48280_ (_16681_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or _48281_ (_07353_, _16681_, _16679_);
  and _48282_ (_16682_, _03043_, _24134_);
  and _48283_ (_16683_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or _48284_ (_07355_, _16683_, _16682_);
  and _48285_ (_16684_, _05478_, _24219_);
  and _48286_ (_16685_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or _48287_ (_27249_, _16685_, _16684_);
  and _48288_ (_16686_, _02502_, _23548_);
  and _48289_ (_16687_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or _48290_ (_07360_, _16687_, _16686_);
  and _48291_ (_16688_, _02478_, _23887_);
  and _48292_ (_16689_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or _48293_ (_27246_, _16689_, _16688_);
  and _48294_ (_16690_, _06129_, _24219_);
  and _48295_ (_16691_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or _48296_ (_07370_, _16691_, _16690_);
  and _48297_ (_16692_, _15561_, _23887_);
  and _48298_ (_16693_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or _48299_ (_27241_, _16693_, _16692_);
  and _48300_ (_16694_, _15888_, _24051_);
  and _48301_ (_16695_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _48302_ (_07391_, _16695_, _16694_);
  and _48303_ (_16696_, _15992_, _24051_);
  and _48304_ (_16697_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  or _48305_ (_07394_, _16697_, _16696_);
  and _48306_ (_16698_, _24496_, _24372_);
  and _48307_ (_16699_, _16698_, _23583_);
  not _48308_ (_16700_, _16698_);
  and _48309_ (_16701_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or _48310_ (_07397_, _16701_, _16699_);
  and _48311_ (_16702_, _02767_, _23887_);
  and _48312_ (_16703_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _48313_ (_07399_, _16703_, _16702_);
  nor _48314_ (_26867_[0], _26630_, rst);
  and _48315_ (_16704_, _24496_, _24140_);
  and _48316_ (_16705_, _16704_, _24089_);
  not _48317_ (_16706_, _16704_);
  and _48318_ (_16707_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or _48319_ (_07403_, _16707_, _16705_);
  and _48320_ (_16708_, _02767_, _23548_);
  and _48321_ (_16709_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _48322_ (_27174_, _16709_, _16708_);
  and _48323_ (_16710_, _15992_, _24089_);
  and _48324_ (_16711_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or _48325_ (_07407_, _16711_, _16710_);
  or _48326_ (_16712_, _08401_, _23880_);
  and _48327_ (_16713_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48328_ (_16714_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _48329_ (_16715_, _16714_, _16713_);
  or _48330_ (_16716_, _16715_, _25608_);
  and _48331_ (_16717_, _16716_, _25617_);
  and _48332_ (_16718_, _16717_, _16712_);
  and _48333_ (_16719_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _48334_ (_16720_, _16719_, _16718_);
  and _48335_ (_07409_, _16720_, _22731_);
  and _48336_ (_16721_, _15992_, _23583_);
  and _48337_ (_16722_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or _48338_ (_26973_, _16722_, _16721_);
  and _48339_ (_16723_, _02045_, _24134_);
  and _48340_ (_16724_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _48341_ (_07414_, _16724_, _16723_);
  and _48342_ (_16725_, _16551_, _23583_);
  and _48343_ (_16726_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or _48344_ (_07418_, _16726_, _16725_);
  and _48345_ (_16727_, _02767_, _24219_);
  and _48346_ (_16728_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _48347_ (_07425_, _16728_, _16727_);
  and _48348_ (_16729_, _11311_, _23887_);
  and _48349_ (_16730_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or _48350_ (_07427_, _16730_, _16729_);
  and _48351_ (_16731_, _24899_, _24301_);
  and _48352_ (_16732_, _16731_, _24134_);
  not _48353_ (_16733_, _16731_);
  and _48354_ (_16734_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or _48355_ (_07433_, _16734_, _16732_);
  and _48356_ (_16735_, _05485_, _23996_);
  and _48357_ (_16736_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _48358_ (_07444_, _16736_, _16735_);
  and _48359_ (_16737_, _11441_, _24051_);
  and _48360_ (_16738_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _48361_ (_07449_, _16738_, _16737_);
  and _48362_ (_16739_, _16551_, _24089_);
  and _48363_ (_16740_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or _48364_ (_07456_, _16740_, _16739_);
  and _48365_ (_16741_, _24451_, _24051_);
  and _48366_ (_16742_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _48367_ (_07462_, _16742_, _16741_);
  and _48368_ (_16743_, _16551_, _24134_);
  and _48369_ (_16744_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or _48370_ (_07469_, _16744_, _16743_);
  and _48371_ (_16745_, _15992_, _23996_);
  and _48372_ (_16746_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or _48373_ (_07471_, _16746_, _16745_);
  and _48374_ (_16747_, _25672_, _23996_);
  and _48375_ (_16748_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _48376_ (_27206_, _16748_, _16747_);
  and _48377_ (_16749_, _25672_, _23583_);
  and _48378_ (_16750_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _48379_ (_07499_, _16750_, _16749_);
  and _48380_ (_16751_, _03241_, _23548_);
  and _48381_ (_16752_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or _48382_ (_07501_, _16752_, _16751_);
  and _48383_ (_16753_, _09670_, _24134_);
  and _48384_ (_16754_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or _48385_ (_07503_, _16754_, _16753_);
  and _48386_ (_16755_, _06208_, _23583_);
  and _48387_ (_16756_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _48388_ (_07506_, _16756_, _16755_);
  and _48389_ (_16757_, _03241_, _24219_);
  and _48390_ (_16758_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  or _48391_ (_07511_, _16758_, _16757_);
  and _48392_ (_16759_, _16541_, _23996_);
  and _48393_ (_16760_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or _48394_ (_07513_, _16760_, _16759_);
  and _48395_ (_16761_, _25637_, _23548_);
  and _48396_ (_16762_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _48397_ (_07515_, _16762_, _16761_);
  and _48398_ (_16763_, _16111_, _23996_);
  and _48399_ (_16764_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or _48400_ (_07528_, _16764_, _16763_);
  and _48401_ (_16765_, _15830_, _24134_);
  and _48402_ (_16766_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _48403_ (_07535_, _16766_, _16765_);
  and _48404_ (_16767_, _25658_, _24051_);
  and _48405_ (_16768_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _48406_ (_07540_, _16768_, _16767_);
  and _48407_ (_16769_, _16111_, _24134_);
  and _48408_ (_16770_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or _48409_ (_07542_, _16770_, _16769_);
  and _48410_ (_16771_, _15888_, _24219_);
  and _48411_ (_16772_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _48412_ (_07544_, _16772_, _16771_);
  and _48413_ (_16773_, _24496_, _24146_);
  and _48414_ (_16774_, _16773_, _23583_);
  not _48415_ (_16775_, _16773_);
  and _48416_ (_16776_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or _48417_ (_07546_, _16776_, _16774_);
  and _48418_ (_16777_, _03241_, _23887_);
  and _48419_ (_16778_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  or _48420_ (_07550_, _16778_, _16777_);
  and _48421_ (_16779_, _03241_, _24089_);
  and _48422_ (_16780_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or _48423_ (_07554_, _16780_, _16779_);
  and _48424_ (_16781_, _25479_, _24636_);
  and _48425_ (_16782_, _16781_, _23504_);
  nor _48426_ (_16783_, _16781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _48427_ (_16784_, _16783_, _16782_);
  nand _48428_ (_16785_, _16784_, _08541_);
  nand _48429_ (_16786_, _25489_, _24082_);
  and _48430_ (_16787_, _16786_, _22731_);
  and _48431_ (_07558_, _16787_, _16785_);
  and _48432_ (_16788_, _25479_, _24533_);
  nand _48433_ (_16789_, _16788_, _23504_);
  or _48434_ (_16790_, _16788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _48435_ (_16791_, _16790_, _08541_);
  and _48436_ (_16792_, _16791_, _16789_);
  and _48437_ (_16793_, _25489_, _23577_);
  or _48438_ (_16794_, _16793_, _16792_);
  and _48439_ (_07562_, _16794_, _22731_);
  and _48440_ (_16795_, _03001_, _24089_);
  and _48441_ (_16796_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _48442_ (_07565_, _16796_, _16795_);
  and _48443_ (_16797_, _03241_, _23583_);
  and _48444_ (_16798_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  or _48445_ (_27172_, _16798_, _16797_);
  and _48446_ (_16799_, _25479_, _24562_);
  nand _48447_ (_16800_, _16799_, _23504_);
  or _48448_ (_16801_, _16799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _48449_ (_16802_, _16801_, _08541_);
  and _48450_ (_16803_, _16802_, _16800_);
  and _48451_ (_16804_, _25489_, _23880_);
  or _48452_ (_16805_, _16804_, _16803_);
  and _48453_ (_07577_, _16805_, _22731_);
  and _48454_ (_16806_, _24451_, _23548_);
  and _48455_ (_16807_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _48456_ (_07580_, _16807_, _16806_);
  and _48457_ (_16808_, _15992_, _23548_);
  and _48458_ (_16809_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or _48459_ (_07586_, _16809_, _16808_);
  and _48460_ (_16810_, _15581_, _23548_);
  and _48461_ (_16811_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or _48462_ (_07588_, _16811_, _16810_);
  nand _48463_ (_16812_, _03797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _48464_ (_16813_, _16812_, _25479_);
  or _48465_ (_16814_, _16813_, _03798_);
  not _48466_ (_16815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _48467_ (_16816_, _25528_, _16815_);
  or _48468_ (_16817_, _16816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _48469_ (_16818_, _16817_, _25479_);
  and _48470_ (_16819_, _16818_, _16814_);
  or _48471_ (_16820_, _16819_, _25489_);
  nand _48472_ (_16821_, _25489_, _24126_);
  and _48473_ (_16822_, _16821_, _22731_);
  and _48474_ (_07603_, _16822_, _16820_);
  and _48475_ (_16823_, _15992_, _24219_);
  and _48476_ (_16824_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  or _48477_ (_07607_, _16824_, _16823_);
  or _48478_ (_16825_, _25550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _48479_ (_16826_, _25541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _48480_ (_16827_, _25543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _48481_ (_16828_, _25544_, _25531_);
  or _48482_ (_16829_, _16828_, _25499_);
  and _48483_ (_16830_, _16829_, _16827_);
  or _48484_ (_16831_, _16830_, _16826_);
  and _48485_ (_16832_, _16831_, _16825_);
  or _48486_ (_16833_, _16832_, _25558_);
  nand _48487_ (_16834_, _25558_, _24126_);
  and _48488_ (_16835_, _16834_, _22731_);
  and _48489_ (_07624_, _16835_, _16833_);
  and _48490_ (_16836_, _24394_, _23887_);
  and _48491_ (_16837_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _48492_ (_07626_, _16837_, _16836_);
  and _48493_ (_16838_, _25479_, _24577_);
  nand _48494_ (_16839_, _16838_, _23504_);
  or _48495_ (_16840_, _16838_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _48496_ (_16841_, _16840_, _08541_);
  and _48497_ (_16842_, _16841_, _16839_);
  and _48498_ (_16843_, _25489_, _24671_);
  or _48499_ (_16844_, _16843_, _16842_);
  and _48500_ (_07639_, _16844_, _22731_);
  and _48501_ (_16845_, _05478_, _23548_);
  and _48502_ (_16846_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or _48503_ (_27250_, _16846_, _16845_);
  and _48504_ (_16847_, _03245_, _23583_);
  and _48505_ (_16848_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or _48506_ (_07646_, _16848_, _16847_);
  and _48507_ (_16849_, _16111_, _23548_);
  and _48508_ (_16850_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or _48509_ (_07648_, _16850_, _16849_);
  and _48510_ (_16851_, _03245_, _23887_);
  and _48511_ (_16852_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or _48512_ (_07868_, _16852_, _16851_);
  and _48513_ (_16853_, _15561_, _23583_);
  and _48514_ (_16854_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or _48515_ (_07870_, _16854_, _16853_);
  and _48516_ (_16855_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _48517_ (_16856_, _16855_, _25523_);
  and _48518_ (_16857_, _25514_, _25507_);
  or _48519_ (_16858_, _16857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _48520_ (_16859_, _16857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _48521_ (_16860_, _16859_, _16858_);
  or _48522_ (_16861_, _16860_, _25531_);
  or _48523_ (_16862_, _16861_, _16856_);
  or _48524_ (_16863_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _48525_ (_16864_, _16863_, _25502_);
  and _48526_ (_16865_, _16864_, _16862_);
  and _48527_ (_16866_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _48528_ (_16867_, _25558_, _24671_);
  or _48529_ (_16868_, _16867_, _16866_);
  or _48530_ (_16869_, _16868_, _16865_);
  and _48531_ (_07875_, _16869_, _22731_);
  and _48532_ (_16870_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _48533_ (_16871_, _16870_, _25523_);
  nand _48534_ (_16872_, _25518_, _25507_);
  and _48535_ (_16873_, _16872_, _08420_);
  nor _48536_ (_16874_, _16873_, _08458_);
  or _48537_ (_16875_, _16874_, _25531_);
  or _48538_ (_16876_, _16875_, _16871_);
  or _48539_ (_16877_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _48540_ (_16878_, _16877_, _25502_);
  and _48541_ (_16879_, _16878_, _16876_);
  and _48542_ (_16880_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _48543_ (_16881_, _16880_, _16879_);
  and _48544_ (_16882_, _08468_, _02700_);
  or _48545_ (_16883_, _16882_, _16881_);
  and _48546_ (_07877_, _16883_, _22731_);
  and _48547_ (_16884_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _48548_ (_16885_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _48549_ (_16886_, _16885_, _25523_);
  and _48550_ (_16887_, _25517_, _25507_);
  or _48551_ (_16888_, _16887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _48552_ (_16889_, _16888_, _16872_);
  or _48553_ (_16890_, _16889_, _25531_);
  or _48554_ (_16891_, _16890_, _16886_);
  or _48555_ (_16892_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _48556_ (_16893_, _16892_, _25502_);
  and _48557_ (_16894_, _16893_, _16891_);
  or _48558_ (_16895_, _16894_, _16884_);
  and _48559_ (_16896_, _08468_, _23577_);
  or _48560_ (_16897_, _16896_, _16895_);
  and _48561_ (_07879_, _16897_, _22731_);
  and _48562_ (_16898_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _48563_ (_16899_, _16898_, _25523_);
  and _48564_ (_16900_, _25516_, _25507_);
  nor _48565_ (_16901_, _16900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _48566_ (_16902_, _16901_, _16887_);
  or _48567_ (_16903_, _16902_, _25531_);
  or _48568_ (_16904_, _16903_, _16899_);
  or _48569_ (_16905_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _48570_ (_16906_, _16905_, _25502_);
  and _48571_ (_16907_, _16906_, _16904_);
  and _48572_ (_16908_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _48573_ (_16909_, _16908_, _16907_);
  and _48574_ (_16910_, _08468_, _23880_);
  or _48575_ (_16911_, _16910_, _16909_);
  and _48576_ (_07881_, _16911_, _22731_);
  and _48577_ (_16912_, _07038_, _24219_);
  and _48578_ (_16913_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _48579_ (_27226_, _16913_, _16912_);
  and _48580_ (_16914_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _48581_ (_16915_, _16914_, _25523_);
  and _48582_ (_16916_, _25515_, _25507_);
  nor _48583_ (_16917_, _16916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _48584_ (_16918_, _16917_, _16900_);
  or _48585_ (_16919_, _16918_, _25531_);
  or _48586_ (_16920_, _16919_, _16915_);
  or _48587_ (_16921_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _48588_ (_16922_, _16921_, _25502_);
  and _48589_ (_16923_, _16922_, _16920_);
  and _48590_ (_16924_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _48591_ (_16925_, _25558_, _02728_);
  or _48592_ (_16926_, _16925_, _16924_);
  or _48593_ (_16927_, _16926_, _16923_);
  and _48594_ (_07884_, _16927_, _22731_);
  and _48595_ (_16928_, _25499_, _23880_);
  and _48596_ (_16929_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48597_ (_16930_, _16929_, _25523_);
  and _48598_ (_16931_, _25508_, _25507_);
  or _48599_ (_16932_, _16931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _48600_ (_16933_, _16932_, _08442_);
  or _48601_ (_16934_, _16933_, _25531_);
  or _48602_ (_16935_, _16934_, _16930_);
  or _48603_ (_16936_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48604_ (_16937_, _16936_, _25502_);
  and _48605_ (_16938_, _16937_, _16935_);
  and _48606_ (_16939_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _48607_ (_16940_, _16939_, _16938_);
  or _48608_ (_16941_, _16940_, _16928_);
  and _48609_ (_07889_, _16941_, _22731_);
  and _48610_ (_16942_, _25507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  not _48611_ (_16943_, _16942_);
  nor _48612_ (_16944_, _16943_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _48613_ (_16945_, _16943_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _48614_ (_16946_, _16945_, _25531_);
  or _48615_ (_16947_, _16946_, _16944_);
  and _48616_ (_16948_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _48617_ (_16949_, _16948_, _25523_);
  or _48618_ (_16950_, _16949_, _16947_);
  or _48619_ (_16951_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _48620_ (_16952_, _16951_, _25502_);
  and _48621_ (_16953_, _16952_, _16950_);
  nor _48622_ (_16954_, _25550_, _23542_);
  and _48623_ (_16955_, _25558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _48624_ (_16956_, _16955_, _16954_);
  or _48625_ (_16957_, _16956_, _16953_);
  and _48626_ (_07891_, _16957_, _22731_);
  or _48627_ (_16958_, _25507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _48628_ (_16959_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _48629_ (_16960_, _16959_, _25522_);
  or _48630_ (_16961_, _16960_, _16943_);
  and _48631_ (_16962_, _16961_, _16958_);
  or _48632_ (_16963_, _16962_, _25531_);
  or _48633_ (_16964_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _48634_ (_16965_, _16964_, _25502_);
  and _48635_ (_16966_, _16965_, _16963_);
  and _48636_ (_16967_, _25499_, _24671_);
  and _48637_ (_16968_, _25558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _48638_ (_16969_, _16968_, _16967_);
  or _48639_ (_16970_, _16969_, _16966_);
  and _48640_ (_07896_, _16970_, _22731_);
  and _48641_ (_16971_, _02996_, _24219_);
  and _48642_ (_16972_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or _48643_ (_07898_, _16972_, _16971_);
  and _48644_ (_16973_, _16111_, _24089_);
  and _48645_ (_16974_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or _48646_ (_07902_, _16974_, _16973_);
  and _48647_ (_16975_, _03245_, _24134_);
  and _48648_ (_16976_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or _48649_ (_07904_, _16976_, _16975_);
  nor _48650_ (_16977_, _25550_, _24043_);
  and _48651_ (_16978_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48652_ (_16979_, _16978_, _25523_);
  nand _48653_ (_16980_, _25511_, _25507_);
  nor _48654_ (_16981_, _16980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _48655_ (_16982_, _16980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _48656_ (_16983_, _16982_, _25531_);
  or _48657_ (_16984_, _16983_, _16981_);
  or _48658_ (_16985_, _16984_, _16979_);
  or _48659_ (_16986_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48660_ (_16987_, _16986_, _25502_);
  and _48661_ (_16988_, _16987_, _16985_);
  and _48662_ (_16989_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _48663_ (_16990_, _16989_, _16988_);
  or _48664_ (_16991_, _16990_, _16977_);
  and _48665_ (_07905_, _16991_, _22731_);
  and _48666_ (_16992_, _16111_, _23583_);
  and _48667_ (_16993_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  or _48668_ (_07908_, _16993_, _16992_);
  and _48669_ (_16994_, _06208_, _24089_);
  and _48670_ (_16995_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _48671_ (_07910_, _16995_, _16994_);
  and _48672_ (_16996_, _25637_, _23996_);
  and _48673_ (_16997_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _48674_ (_07912_, _16997_, _16996_);
  nor _48675_ (_16998_, _25550_, _24126_);
  and _48676_ (_16999_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _48677_ (_17000_, _16999_, _25523_);
  and _48678_ (_17001_, _25512_, _25507_);
  nor _48679_ (_17002_, _17001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _48680_ (_17003_, _17002_, _25582_);
  or _48681_ (_17004_, _17003_, _25531_);
  or _48682_ (_17005_, _17004_, _17000_);
  or _48683_ (_17006_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _48684_ (_17007_, _17006_, _25502_);
  and _48685_ (_17008_, _17007_, _17005_);
  and _48686_ (_17009_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _48687_ (_17010_, _17009_, _17008_);
  or _48688_ (_17011_, _17010_, _16998_);
  and _48689_ (_07914_, _17011_, _22731_);
  nor _48690_ (_17012_, _25550_, _24082_);
  and _48691_ (_17013_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _48692_ (_17014_, _17013_, _25523_);
  and _48693_ (_17015_, _25510_, _25507_);
  or _48694_ (_17016_, _17015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _48695_ (_17017_, _17016_, _16980_);
  or _48696_ (_17018_, _17017_, _25531_);
  or _48697_ (_17019_, _17018_, _17014_);
  or _48698_ (_17020_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _48699_ (_17021_, _17020_, _25502_);
  and _48700_ (_17022_, _17021_, _17019_);
  and _48701_ (_17023_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _48702_ (_17024_, _17023_, _17022_);
  or _48703_ (_17025_, _17024_, _17012_);
  and _48704_ (_07917_, _17025_, _22731_);
  and _48705_ (_17026_, _15830_, _23996_);
  and _48706_ (_17027_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _48707_ (_07952_, _17027_, _17026_);
  and _48708_ (_17028_, _16535_, _23548_);
  and _48709_ (_17029_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or _48710_ (_07959_, _17029_, _17028_);
  and _48711_ (_17030_, _15561_, _24089_);
  and _48712_ (_17031_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or _48713_ (_07961_, _17031_, _17030_);
  and _48714_ (_17032_, _24372_, _24098_);
  and _48715_ (_17033_, _17032_, _24219_);
  not _48716_ (_17034_, _17032_);
  and _48717_ (_17035_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or _48718_ (_07965_, _17035_, _17033_);
  and _48719_ (_17036_, _24146_, _24098_);
  and _48720_ (_17037_, _17036_, _23996_);
  not _48721_ (_17038_, _17036_);
  and _48722_ (_17039_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or _48723_ (_07968_, _17039_, _17037_);
  and _48724_ (_17040_, _17036_, _23548_);
  and _48725_ (_17041_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or _48726_ (_07972_, _17041_, _17040_);
  and _48727_ (_17042_, _24140_, _24098_);
  and _48728_ (_17043_, _17042_, _24089_);
  not _48729_ (_17044_, _17042_);
  and _48730_ (_17045_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _48731_ (_07975_, _17045_, _17043_);
  and _48732_ (_17046_, _24159_, _22982_);
  and _48733_ (_17047_, _17046_, _24089_);
  not _48734_ (_17048_, _17046_);
  and _48735_ (_17049_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _48736_ (_07981_, _17049_, _17047_);
  and _48737_ (_17050_, _17046_, _23887_);
  and _48738_ (_17051_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _48739_ (_07983_, _17051_, _17050_);
  and _48740_ (_17052_, _24297_, _22982_);
  and _48741_ (_17053_, _17052_, _24089_);
  not _48742_ (_17054_, _17052_);
  and _48743_ (_17055_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or _48744_ (_07988_, _17055_, _17053_);
  and _48745_ (_17056_, _17052_, _23887_);
  and _48746_ (_17057_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or _48747_ (_07990_, _17057_, _17056_);
  and _48748_ (_17058_, _24016_, _22982_);
  and _48749_ (_17059_, _17058_, _24051_);
  not _48750_ (_17060_, _17058_);
  and _48751_ (_17061_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or _48752_ (_07993_, _17061_, _17059_);
  and _48753_ (_17062_, _17058_, _23583_);
  and _48754_ (_17063_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or _48755_ (_07995_, _17063_, _17062_);
  and _48756_ (_17064_, _17058_, _24219_);
  and _48757_ (_17065_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or _48758_ (_07997_, _17065_, _17064_);
  and _48759_ (_17066_, _24236_, _22982_);
  and _48760_ (_17067_, _17066_, _24134_);
  not _48761_ (_17068_, _17066_);
  and _48762_ (_17069_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _48763_ (_08002_, _17069_, _17067_);
  and _48764_ (_17070_, _17066_, _23887_);
  and _48765_ (_17071_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _48766_ (_08005_, _17071_, _17070_);
  and _48767_ (_17072_, _24899_, _22982_);
  and _48768_ (_17073_, _17072_, _24134_);
  not _48769_ (_17074_, _17072_);
  and _48770_ (_17075_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or _48771_ (_08012_, _17075_, _17073_);
  and _48772_ (_17076_, _11360_, _24051_);
  and _48773_ (_17077_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _48774_ (_27079_, _17077_, _17076_);
  and _48775_ (_17078_, _24474_, _22982_);
  and _48776_ (_17079_, _17078_, _24134_);
  not _48777_ (_17080_, _17078_);
  and _48778_ (_17081_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _48779_ (_08020_, _17081_, _17079_);
  and _48780_ (_17082_, _17078_, _24089_);
  and _48781_ (_17083_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _48782_ (_27285_, _17083_, _17082_);
  and _48783_ (_17084_, _17078_, _24219_);
  and _48784_ (_17085_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _48785_ (_08023_, _17085_, _17084_);
  nand _48786_ (_17086_, _25603_, _24126_);
  and _48787_ (_17087_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _48788_ (_17088_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _48789_ (_17089_, _17088_, _17087_);
  or _48790_ (_17090_, _17089_, _25603_);
  and _48791_ (_17091_, _17090_, _22731_);
  and _48792_ (_08237_, _17091_, _17086_);
  and _48793_ (_17092_, _24057_, _23996_);
  and _48794_ (_17093_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or _48795_ (_08238_, _17093_, _17092_);
  and _48796_ (_17094_, _03245_, _24051_);
  and _48797_ (_17095_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or _48798_ (_08240_, _17095_, _17094_);
  nand _48799_ (_17096_, _25603_, _24043_);
  and _48800_ (_17097_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _48801_ (_17098_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _48802_ (_17099_, _17098_, _17097_);
  or _48803_ (_17100_, _17099_, _25603_);
  and _48804_ (_17101_, _17100_, _22731_);
  and _48805_ (_08242_, _17101_, _17096_);
  and _48806_ (_17102_, _24349_, _22982_);
  and _48807_ (_17103_, _17102_, _24089_);
  not _48808_ (_17104_, _17102_);
  and _48809_ (_17105_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _48810_ (_08247_, _17105_, _17103_);
  and _48811_ (_17106_, _16000_, _24089_);
  and _48812_ (_17107_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or _48813_ (_08249_, _17107_, _17106_);
  and _48814_ (_17108_, _16000_, _23583_);
  and _48815_ (_17109_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or _48816_ (_08253_, _17109_, _17108_);
  and _48817_ (_17110_, _23941_, _22982_);
  and _48818_ (_17111_, _17110_, _24051_);
  not _48819_ (_17112_, _17110_);
  and _48820_ (_17113_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or _48821_ (_27291_, _17113_, _17111_);
  and _48822_ (_17114_, _03255_, _24134_);
  and _48823_ (_17115_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or _48824_ (_08256_, _17115_, _17114_);
  and _48825_ (_17116_, _16535_, _23887_);
  and _48826_ (_17117_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or _48827_ (_08259_, _17117_, _17116_);
  and _48828_ (_17118_, _03255_, _24051_);
  and _48829_ (_17119_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _48830_ (_08261_, _17119_, _17118_);
  or _48831_ (_17120_, _25617_, _23577_);
  and _48832_ (_17121_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _48833_ (_17122_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _48834_ (_17123_, _17122_, _17121_);
  or _48835_ (_17124_, _17123_, _25603_);
  and _48836_ (_17125_, _17124_, _22731_);
  and _48837_ (_08266_, _17125_, _17120_);
  or _48838_ (_17126_, _25617_, _23880_);
  and _48839_ (_17127_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _48840_ (_17128_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _48841_ (_17129_, _17128_, _17127_);
  or _48842_ (_17130_, _17129_, _25603_);
  and _48843_ (_17131_, _17130_, _22731_);
  and _48844_ (_08268_, _17131_, _17126_);
  and _48845_ (_17132_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _48846_ (_17133_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _48847_ (_17134_, _17133_, _17132_);
  or _48848_ (_17135_, _17134_, _25603_);
  nand _48849_ (_17136_, _25603_, _23542_);
  and _48850_ (_17137_, _17136_, _22731_);
  and _48851_ (_08270_, _17137_, _17135_);
  and _48852_ (_17138_, _03255_, _24089_);
  and _48853_ (_17139_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or _48854_ (_08272_, _17139_, _17138_);
  and _48855_ (_17140_, _17036_, _23583_);
  and _48856_ (_17141_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or _48857_ (_08275_, _17141_, _17140_);
  and _48858_ (_17142_, _16000_, _24134_);
  and _48859_ (_17143_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or _48860_ (_08278_, _17143_, _17142_);
  and _48861_ (_17144_, _16000_, _24051_);
  and _48862_ (_17145_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _48863_ (_08280_, _17145_, _17144_);
  and _48864_ (_17146_, _16535_, _24051_);
  and _48865_ (_17147_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or _48866_ (_08284_, _17147_, _17146_);
  and _48867_ (_17148_, _17042_, _23548_);
  and _48868_ (_17149_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _48869_ (_27301_, _17149_, _17148_);
  nor _48870_ (_17150_, _08401_, _24043_);
  and _48871_ (_17151_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48872_ (_17152_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _48873_ (_17153_, _17152_, _17151_);
  nor _48874_ (_17154_, _17153_, _25608_);
  or _48875_ (_17155_, _17154_, _08404_);
  or _48876_ (_17156_, _17155_, _17150_);
  or _48877_ (_17157_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48878_ (_17158_, _17157_, _22731_);
  and _48879_ (_08288_, _17158_, _17156_);
  and _48880_ (_17159_, _17046_, _24134_);
  and _48881_ (_17160_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _48882_ (_08290_, _17160_, _17159_);
  and _48883_ (_17161_, _02364_, _24219_);
  and _48884_ (_17162_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _48885_ (_08369_, _17162_, _17161_);
  and _48886_ (_17163_, _02364_, _23548_);
  and _48887_ (_17164_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _48888_ (_08381_, _17164_, _17163_);
  not _48889_ (_17165_, _23855_);
  or _48890_ (_26842_[1], _02006_, _17165_);
  and _48891_ (_17166_, _24142_, _24051_);
  and _48892_ (_17167_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or _48893_ (_08393_, _17167_, _17166_);
  and _48894_ (_17168_, _22734_, _22735_);
  and _48895_ (_17169_, _17168_, _26571_);
  and _48896_ (_17170_, _01432_, _01411_);
  or _48897_ (_17171_, _17170_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _48898_ (_17172_, _01391_, _01402_);
  and _48899_ (_17173_, _01475_, _17172_);
  and _48900_ (_17174_, _01432_, _01526_);
  and _48901_ (_17175_, _01502_, _01420_);
  or _48902_ (_17176_, _17175_, _17174_);
  or _48903_ (_17177_, _17176_, _17173_);
  or _48904_ (_17178_, _17177_, _17171_);
  and _48905_ (_17179_, _17178_, _17169_);
  nor _48906_ (_17180_, _17168_, _26571_);
  or _48907_ (_17181_, _17180_, rst);
  or _48908_ (_26843_[0], _17181_, _17179_);
  or _48909_ (_17182_, _01985_, _24253_);
  or _48910_ (_17183_, _02385_, _24275_);
  or _48911_ (_17184_, _17183_, _17182_);
  and _48912_ (_17185_, _17184_, _22737_);
  and _48913_ (_17186_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _48914_ (_17187_, _17186_, _02359_);
  or _48915_ (_17188_, _17187_, _17185_);
  and _48916_ (_26846_[1], _17188_, _22731_);
  and _48917_ (_17189_, _23890_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or _48918_ (_17190_, _26576_, _00287_);
  or _48919_ (_17191_, _17190_, _01979_);
  or _48920_ (_17192_, _00240_, _04800_);
  or _48921_ (_17193_, _26584_, _23894_);
  or _48922_ (_17194_, _26742_, _23923_);
  or _48923_ (_17195_, _17194_, _17193_);
  or _48924_ (_17196_, _17195_, _17192_);
  or _48925_ (_17197_, _17196_, _17191_);
  and _48926_ (_17198_, _17197_, _23855_);
  or _48927_ (_26845_, _17198_, _17189_);
  and _48928_ (_17199_, _05478_, _23887_);
  and _48929_ (_17200_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or _48930_ (_08400_, _17200_, _17199_);
  and _48931_ (_17201_, _05478_, _23583_);
  and _48932_ (_17202_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or _48933_ (_08408_, _17202_, _17201_);
  and _48934_ (_17203_, _24409_, _24051_);
  and _48935_ (_17204_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or _48936_ (_08410_, _17204_, _17203_);
  and _48937_ (_17205_, _09717_, _24134_);
  and _48938_ (_17206_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _48939_ (_08597_, _17206_, _17205_);
  or _48940_ (_17207_, _04786_, _01978_);
  or _48941_ (_17208_, _24267_, _23917_);
  or _48942_ (_17209_, _17208_, _17207_);
  or _48943_ (_17210_, _23815_, _23790_);
  or _48944_ (_17211_, _26694_, _23919_);
  or _48945_ (_17212_, _17211_, _17210_);
  nand _48946_ (_17213_, _23838_, _01990_);
  nand _48947_ (_17214_, _17213_, _26699_);
  or _48948_ (_17215_, _17214_, _03906_);
  or _48949_ (_17216_, _23836_, _23833_);
  or _48950_ (_17217_, _17216_, _17215_);
  or _48951_ (_17218_, _17217_, _17212_);
  or _48952_ (_17219_, _26754_, _26731_);
  and _48953_ (_17220_, _23927_, _23687_);
  or _48954_ (_17221_, _17220_, _01979_);
  or _48955_ (_17222_, _17221_, _17219_);
  or _48956_ (_17223_, _17222_, _09756_);
  or _48957_ (_17224_, _17223_, _17218_);
  or _48958_ (_17225_, _17224_, _17209_);
  and _48959_ (_17226_, _17225_, _22737_);
  and _48960_ (_17227_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _48961_ (_17228_, _17227_, _02010_);
  or _48962_ (_17229_, _17228_, _17226_);
  and _48963_ (_26846_[0], _17229_, _22731_);
  and _48964_ (_17230_, _09717_, _23996_);
  and _48965_ (_17231_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _48966_ (_08602_, _17231_, _17230_);
  or _48967_ (_17232_, _23703_, _26679_);
  or _48968_ (_17233_, _22736_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _48969_ (_17234_, _17233_, _22731_);
  and _48970_ (_26844_[4], _17234_, _17232_);
  and _48971_ (_17235_, _09717_, _24051_);
  and _48972_ (_17236_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _48973_ (_27072_, _17236_, _17235_);
  and _48974_ (_26841_[0], _26713_, _22731_);
  or _48975_ (_17237_, _23765_, _26679_);
  or _48976_ (_17238_, _22736_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _48977_ (_17239_, _17238_, _22731_);
  and _48978_ (_26844_[5], _17239_, _17237_);
  and _48979_ (_17240_, _24350_, _23548_);
  and _48980_ (_17241_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _48981_ (_27057_, _17241_, _17240_);
  or _48982_ (_17242_, _23660_, _26679_);
  or _48983_ (_17243_, _22736_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _48984_ (_17244_, _17243_, _22731_);
  and _48985_ (_26844_[1], _17244_, _17242_);
  and _48986_ (_17245_, _02364_, _24051_);
  and _48987_ (_17246_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _48988_ (_08629_, _17246_, _17245_);
  or _48989_ (_17247_, _23639_, _26679_);
  or _48990_ (_17248_, _22736_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _48991_ (_17249_, _17248_, _22731_);
  and _48992_ (_26844_[2], _17249_, _17247_);
  and _48993_ (_17250_, _02364_, _24134_);
  and _48994_ (_17251_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _48995_ (_08634_, _17251_, _17250_);
  and _48996_ (_17252_, _05460_, _24134_);
  and _48997_ (_17253_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _48998_ (_08650_, _17253_, _17252_);
  and _48999_ (_17254_, _05460_, _23996_);
  and _49000_ (_17255_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or _49001_ (_08655_, _17255_, _17254_);
  and _49002_ (_17256_, _03001_, _24051_);
  and _49003_ (_17257_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _49004_ (_27216_, _17257_, _17256_);
  nand _49005_ (_17258_, _16094_, _24082_);
  nor _49006_ (_17259_, _16100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _49007_ (_17260_, _17259_, _16101_);
  or _49008_ (_17261_, _17260_, _02616_);
  and _49009_ (_17262_, _17261_, _02295_);
  and _49010_ (_17263_, _17262_, _17258_);
  and _49011_ (_17264_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _49012_ (_08662_, _17264_, _17263_);
  and _49013_ (_17265_, _24442_, _24219_);
  and _49014_ (_17266_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or _49015_ (_08667_, _17266_, _17265_);
  and _49016_ (_17267_, _17052_, _24134_);
  and _49017_ (_17268_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or _49018_ (_08694_, _17268_, _17267_);
  and _49019_ (_17269_, _17058_, _23996_);
  and _49020_ (_17270_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or _49021_ (_27297_, _17270_, _17269_);
  nor _49022_ (_17271_, _08401_, _24082_);
  and _49023_ (_17272_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49024_ (_17273_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _49025_ (_17274_, _17273_, _17272_);
  nor _49026_ (_17275_, _17274_, _25608_);
  or _49027_ (_17276_, _17275_, _08404_);
  or _49028_ (_17277_, _17276_, _17271_);
  or _49029_ (_17278_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49030_ (_17279_, _17278_, _22731_);
  and _49031_ (_08701_, _17279_, _17277_);
  or _49032_ (_17280_, _08401_, _23577_);
  and _49033_ (_17281_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49034_ (_17282_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _49035_ (_17283_, _17282_, _17281_);
  or _49036_ (_17284_, _17283_, _25608_);
  and _49037_ (_17285_, _17284_, _25617_);
  and _49038_ (_17286_, _17285_, _17280_);
  and _49039_ (_17287_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _49040_ (_17288_, _17287_, _17286_);
  and _49041_ (_08711_, _17288_, _22731_);
  and _49042_ (_17289_, _24142_, _23887_);
  and _49043_ (_17290_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or _49044_ (_08728_, _17290_, _17289_);
  or _49045_ (_17291_, _23681_, _26679_);
  or _49046_ (_17292_, _22736_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _49047_ (_17293_, _17292_, _22731_);
  and _49048_ (_26844_[0], _17293_, _17291_);
  and _49049_ (_17294_, _05460_, _24089_);
  and _49050_ (_17295_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _49051_ (_08738_, _17295_, _17294_);
  nand _49052_ (_17296_, _23615_, _22736_);
  or _49053_ (_17297_, _22736_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _49054_ (_17298_, _17297_, _22731_);
  and _49055_ (_26844_[3], _17298_, _17296_);
  or _49056_ (_17299_, _23745_, _26679_);
  or _49057_ (_17300_, _22736_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _49058_ (_17301_, _17300_, _22731_);
  and _49059_ (_26844_[6], _17301_, _17299_);
  and _49060_ (_17302_, _03355_, _24219_);
  and _49061_ (_17303_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _49062_ (_08780_, _17303_, _17302_);
  and _49063_ (_17304_, _11360_, _24089_);
  and _49064_ (_17305_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _49065_ (_08782_, _17305_, _17304_);
  and _49066_ (_17306_, _17110_, _23548_);
  and _49067_ (_17307_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or _49068_ (_08799_, _17307_, _17306_);
  and _49069_ (_17308_, _17072_, _23583_);
  and _49070_ (_17309_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or _49071_ (_08802_, _17309_, _17308_);
  and _49072_ (_17310_, _17102_, _24134_);
  and _49073_ (_17311_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _49074_ (_08809_, _17311_, _17310_);
  and _49075_ (_17312_, _17032_, _23548_);
  and _49076_ (_17313_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or _49077_ (_08812_, _17313_, _17312_);
  and _49078_ (_17314_, _17042_, _24051_);
  and _49079_ (_17315_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _49080_ (_08814_, _17315_, _17314_);
  and _49081_ (_17316_, _24237_, _23548_);
  and _49082_ (_17317_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _49083_ (_08817_, _17317_, _17316_);
  and _49084_ (_17318_, _03245_, _24219_);
  and _49085_ (_17319_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or _49086_ (_27169_, _17319_, _17318_);
  and _49087_ (_17320_, _16731_, _23996_);
  and _49088_ (_17321_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or _49089_ (_08825_, _17321_, _17320_);
  nor _49090_ (_26867_[7], _00139_, rst);
  and _49091_ (_17322_, _17072_, _24219_);
  and _49092_ (_17323_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or _49093_ (_08847_, _17323_, _17322_);
  and _49094_ (_17324_, _17102_, _24219_);
  and _49095_ (_17325_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _49096_ (_08851_, _17325_, _17324_);
  and _49097_ (_17326_, _17052_, _23996_);
  and _49098_ (_17327_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or _49099_ (_08855_, _17327_, _17326_);
  and _49100_ (_17328_, _16185_, _23996_);
  and _49101_ (_17329_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or _49102_ (_08862_, _17329_, _17328_);
  and _49103_ (_17330_, _08523_, _24219_);
  and _49104_ (_17331_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or _49105_ (_08865_, _17331_, _17330_);
  and _49106_ (_17332_, _11360_, _23996_);
  and _49107_ (_17333_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or _49108_ (_08873_, _17333_, _17332_);
  and _49109_ (_17334_, _24297_, _24098_);
  and _49110_ (_17335_, _17334_, _24089_);
  not _49111_ (_17336_, _17334_);
  and _49112_ (_17337_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _49113_ (_08887_, _17337_, _17335_);
  and _49114_ (_17338_, _24098_, _24016_);
  and _49115_ (_17339_, _17338_, _24134_);
  not _49116_ (_17340_, _17338_);
  and _49117_ (_17341_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _49118_ (_08892_, _17341_, _17339_);
  and _49119_ (_17342_, _17338_, _23548_);
  and _49120_ (_17343_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _49121_ (_08896_, _17343_, _17342_);
  and _49122_ (_17344_, _24236_, _24098_);
  and _49123_ (_17345_, _17344_, _23996_);
  not _49124_ (_17346_, _17344_);
  and _49125_ (_17347_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or _49126_ (_26910_, _17347_, _17345_);
  and _49127_ (_17348_, _03255_, _23996_);
  and _49128_ (_17349_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _49129_ (_08903_, _17349_, _17348_);
  and _49130_ (_17350_, _16185_, _24134_);
  and _49131_ (_17351_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or _49132_ (_08905_, _17351_, _17350_);
  nand _49133_ (_17352_, _25608_, _24210_);
  or _49134_ (_17353_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _49135_ (_17354_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49136_ (_17355_, _17354_, _17353_);
  or _49137_ (_17356_, _17355_, _25608_);
  and _49138_ (_17357_, _17356_, _17352_);
  or _49139_ (_17358_, _17357_, _08404_);
  or _49140_ (_17359_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _49141_ (_17360_, _17359_, _22731_);
  and _49142_ (_08907_, _17360_, _17358_);
  and _49143_ (_17361_, _16535_, _24134_);
  and _49144_ (_17362_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or _49145_ (_08912_, _17362_, _17361_);
  and _49146_ (_17363_, _24349_, _24098_);
  and _49147_ (_17364_, _17363_, _24134_);
  not _49148_ (_17365_, _17363_);
  and _49149_ (_17366_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or _49150_ (_08923_, _17366_, _17364_);
  and _49151_ (_17367_, _17363_, _23583_);
  and _49152_ (_17368_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or _49153_ (_08925_, _17368_, _17367_);
  and _49154_ (_17369_, _24098_, _23941_);
  and _49155_ (_17370_, _17369_, _24089_);
  not _49156_ (_17371_, _17369_);
  and _49157_ (_17372_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _49158_ (_08932_, _17372_, _17370_);
  and _49159_ (_17373_, _15581_, _23887_);
  and _49160_ (_17374_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or _49161_ (_08947_, _17374_, _17373_);
  and _49162_ (_17375_, _05478_, _24089_);
  and _49163_ (_17376_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or _49164_ (_08949_, _17376_, _17375_);
  and _49165_ (_17377_, _24518_, _24134_);
  and _49166_ (_17378_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or _49167_ (_27220_, _17378_, _17377_);
  and _49168_ (_26840_[7], _23724_, _22731_);
  and _49169_ (_17379_, _24899_, _24098_);
  and _49170_ (_17380_, _17379_, _24051_);
  not _49171_ (_17381_, _17379_);
  and _49172_ (_17382_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _49173_ (_26903_, _17382_, _17380_);
  and _49174_ (_17383_, _17379_, _24219_);
  and _49175_ (_17384_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _49176_ (_08986_, _17384_, _17383_);
  and _49177_ (_17385_, _24474_, _24098_);
  and _49178_ (_17386_, _17385_, _24134_);
  not _49179_ (_17387_, _17385_);
  and _49180_ (_17388_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or _49181_ (_08989_, _17388_, _17386_);
  and _49182_ (_17389_, _17385_, _23548_);
  and _49183_ (_17390_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or _49184_ (_08992_, _17390_, _17389_);
  and _49185_ (_17391_, _24223_, _24098_);
  and _49186_ (_17392_, _17391_, _24089_);
  not _49187_ (_17393_, _17391_);
  and _49188_ (_17394_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or _49189_ (_08995_, _17394_, _17392_);
  and _49190_ (_17395_, _24319_, _24098_);
  and _49191_ (_17396_, _17395_, _23996_);
  not _49192_ (_17397_, _17395_);
  and _49193_ (_17398_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or _49194_ (_08999_, _17398_, _17396_);
  and _49195_ (_17399_, _16000_, _23548_);
  and _49196_ (_17400_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or _49197_ (_09002_, _17400_, _17399_);
  and _49198_ (_17401_, _03269_, _23996_);
  and _49199_ (_17402_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or _49200_ (_09004_, _17402_, _17401_);
  and _49201_ (_17403_, _17395_, _24089_);
  and _49202_ (_17404_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or _49203_ (_09009_, _17404_, _17403_);
  and _49204_ (_17405_, _16541_, _23887_);
  and _49205_ (_17406_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or _49206_ (_09014_, _17406_, _17405_);
  and _49207_ (_17407_, _16541_, _23548_);
  and _49208_ (_17408_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or _49209_ (_09017_, _17408_, _17407_);
  and _49210_ (_17409_, _17395_, _23548_);
  and _49211_ (_17410_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or _49212_ (_09034_, _17410_, _17409_);
  and _49213_ (_17411_, _24098_, _22974_);
  and _49214_ (_17412_, _17411_, _24134_);
  not _49215_ (_17413_, _17411_);
  and _49216_ (_17414_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _49217_ (_09038_, _17414_, _17412_);
  and _49218_ (_17415_, _17411_, _23583_);
  and _49219_ (_17416_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _49220_ (_09042_, _17416_, _17415_);
  and _49221_ (_17417_, _24098_, _24056_);
  and _49222_ (_17418_, _17417_, _24051_);
  not _49223_ (_17419_, _17417_);
  and _49224_ (_17420_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _49225_ (_26900_, _17420_, _17418_);
  and _49226_ (_17421_, _17417_, _23583_);
  and _49227_ (_17422_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _49228_ (_09048_, _17422_, _17421_);
  and _49229_ (_17423_, _16000_, _24219_);
  and _49230_ (_17424_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _49231_ (_09056_, _17424_, _17423_);
  and _49232_ (_17425_, _17334_, _23548_);
  and _49233_ (_17426_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _49234_ (_09057_, _17426_, _17425_);
  and _49235_ (_17427_, _03269_, _24134_);
  and _49236_ (_17428_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or _49237_ (_09059_, _17428_, _17427_);
  and _49238_ (_17429_, _03269_, _24051_);
  and _49239_ (_17430_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  or _49240_ (_09061_, _17430_, _17429_);
  and _49241_ (_17431_, _16121_, _23583_);
  and _49242_ (_17432_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _49243_ (_09063_, _17432_, _17431_);
  and _49244_ (_17433_, _16185_, _23548_);
  and _49245_ (_17434_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or _49246_ (_09069_, _17434_, _17433_);
  and _49247_ (_17435_, _17338_, _23583_);
  and _49248_ (_17436_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _49249_ (_26913_, _17436_, _17435_);
  nand _49250_ (_17437_, _16094_, _23989_);
  or _49251_ (_17438_, _02267_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _49252_ (_17439_, _02268_, _15660_);
  and _49253_ (_17440_, _17439_, _17438_);
  and _49254_ (_17441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _49255_ (_17442_, _02277_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not _49256_ (_17443_, _02271_);
  nor _49257_ (_17444_, _02278_, _17443_);
  and _49258_ (_17445_, _17444_, _17442_);
  or _49259_ (_17446_, _17445_, _17441_);
  or _49260_ (_17447_, _17446_, _17440_);
  or _49261_ (_17448_, _17447_, _02616_);
  and _49262_ (_17449_, _17448_, _02295_);
  and _49263_ (_17450_, _17449_, _17437_);
  and _49264_ (_17451_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _49265_ (_09079_, _17451_, _17450_);
  and _49266_ (_17452_, _11360_, _24219_);
  and _49267_ (_17453_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or _49268_ (_09096_, _17453_, _17452_);
  and _49269_ (_17454_, _08435_, _23887_);
  and _49270_ (_17455_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or _49271_ (_09103_, _17455_, _17454_);
  and _49272_ (_17456_, _17344_, _23887_);
  and _49273_ (_17457_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or _49274_ (_26907_, _17457_, _17456_);
  and _49275_ (_17458_, _17363_, _24219_);
  and _49276_ (_17459_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or _49277_ (_09108_, _17459_, _17458_);
  and _49278_ (_17460_, _17369_, _23548_);
  and _49279_ (_17461_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _49280_ (_26904_, _17461_, _17460_);
  and _49281_ (_17462_, _17379_, _23887_);
  and _49282_ (_17463_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _49283_ (_09112_, _17463_, _17462_);
  and _49284_ (_17464_, _17385_, _23583_);
  and _49285_ (_17465_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or _49286_ (_09113_, _17465_, _17464_);
  and _49287_ (_17466_, _16529_, _24219_);
  and _49288_ (_17467_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _49289_ (_09119_, _17467_, _17466_);
  and _49290_ (_17468_, _16185_, _24219_);
  and _49291_ (_17469_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or _49292_ (_09122_, _17469_, _17468_);
  and _49293_ (_17470_, _17417_, _23996_);
  and _49294_ (_17471_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _49295_ (_09130_, _17471_, _17470_);
  and _49296_ (_17472_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _49297_ (_17473_, _17472_, _26165_);
  and _49298_ (_17474_, _17472_, _26165_);
  or _49299_ (_17475_, _17474_, _17473_);
  and _49300_ (_09133_, _17475_, _22731_);
  or _49301_ (_17476_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _49302_ (_17477_, _17476_, _22731_);
  nand _49303_ (_17478_, _24189_, _24043_);
  and _49304_ (_09136_, _17478_, _17477_);
  and _49305_ (_17479_, _17334_, _24051_);
  and _49306_ (_17480_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _49307_ (_09139_, _17480_, _17479_);
  and _49308_ (_09141_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _22731_);
  and _49309_ (_09145_, _00855_, _22731_);
  and _49310_ (_09148_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _22731_);
  or _49311_ (_17481_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _49312_ (_17482_, _17472_, rst);
  and _49313_ (_09152_, _17482_, _17481_);
  and _49314_ (_17483_, _16529_, _23887_);
  and _49315_ (_17484_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _49316_ (_09157_, _17484_, _17483_);
  and _49317_ (_17485_, _03255_, _23887_);
  and _49318_ (_17486_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _49319_ (_09159_, _17486_, _17485_);
  and _49320_ (_17487_, _17363_, _24089_);
  and _49321_ (_17488_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or _49322_ (_09177_, _17488_, _17487_);
  and _49323_ (_17489_, _17369_, _24051_);
  and _49324_ (_17490_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _49325_ (_09180_, _17490_, _17489_);
  and _49326_ (_17491_, _17385_, _23996_);
  and _49327_ (_17492_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or _49328_ (_09183_, _17492_, _17491_);
  and _49329_ (_17493_, _17395_, _23887_);
  and _49330_ (_17494_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or _49331_ (_09188_, _17494_, _17493_);
  and _49332_ (_17495_, _17417_, _24219_);
  and _49333_ (_17496_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _49334_ (_09191_, _17496_, _17495_);
  and _49335_ (_17497_, _16529_, _24089_);
  and _49336_ (_17498_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _49337_ (_09196_, _17498_, _17497_);
  and _49338_ (_17499_, _17379_, _24134_);
  and _49339_ (_17500_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _49340_ (_09198_, _17500_, _17499_);
  and _49341_ (_17501_, _16529_, _24134_);
  and _49342_ (_17502_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _49343_ (_09201_, _17502_, _17501_);
  and _49344_ (_17503_, _25637_, _24134_);
  and _49345_ (_17504_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _49346_ (_09207_, _17504_, _17503_);
  and _49347_ (_17505_, _17391_, _23996_);
  and _49348_ (_17506_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or _49349_ (_09209_, _17506_, _17505_);
  and _49350_ (_17507_, _17110_, _23996_);
  and _49351_ (_17508_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or _49352_ (_09211_, _17508_, _17507_);
  and _49353_ (_17509_, _25637_, _24089_);
  and _49354_ (_17510_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _49355_ (_09214_, _17510_, _17509_);
  and _49356_ (_17511_, _17391_, _24051_);
  and _49357_ (_17512_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or _49358_ (_09216_, _17512_, _17511_);
  and _49359_ (_17513_, _16121_, _24134_);
  and _49360_ (_17514_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _49361_ (_09218_, _17514_, _17513_);
  and _49362_ (_17515_, _03255_, _23548_);
  and _49363_ (_17516_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _49364_ (_09220_, _17516_, _17515_);
  and _49365_ (_17517_, _03255_, _24219_);
  and _49366_ (_17518_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or _49367_ (_09224_, _17518_, _17517_);
  and _49368_ (_17519_, _17110_, _24089_);
  and _49369_ (_17520_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or _49370_ (_09226_, _17520_, _17519_);
  and _49371_ (_17521_, _16185_, _24089_);
  and _49372_ (_17522_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or _49373_ (_09228_, _17522_, _17521_);
  and _49374_ (_17523_, _25672_, _24134_);
  and _49375_ (_17524_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _49376_ (_09230_, _17524_, _17523_);
  and _49377_ (_17525_, _16185_, _23583_);
  and _49378_ (_17526_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _49379_ (_09232_, _17526_, _17525_);
  and _49380_ (_17527_, _16731_, _23887_);
  and _49381_ (_17528_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or _49382_ (_09256_, _17528_, _17527_);
  and _49383_ (_17529_, _16731_, _23548_);
  and _49384_ (_17530_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or _49385_ (_09268_, _17530_, _17529_);
  and _49386_ (_17531_, _08559_, _23996_);
  and _49387_ (_17532_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or _49388_ (_09270_, _17532_, _17531_);
  and _49389_ (_17533_, _16731_, _24051_);
  and _49390_ (_17534_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or _49391_ (_09276_, _17534_, _17533_);
  and _49392_ (_17535_, _16731_, _24089_);
  and _49393_ (_17536_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or _49394_ (_27223_, _17536_, _17535_);
  and _49395_ (_17537_, _24155_, _23996_);
  and _49396_ (_17538_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or _49397_ (_09287_, _17538_, _17537_);
  and _49398_ (_17539_, _11360_, _23887_);
  and _49399_ (_17540_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _49400_ (_27078_, _17540_, _17539_);
  and _49401_ (_17541_, _11360_, _23548_);
  and _49402_ (_17542_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _49403_ (_09317_, _17542_, _17541_);
  and _49404_ (_17543_, _04812_, _24219_);
  and _49405_ (_17544_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _49406_ (_09328_, _17544_, _17543_);
  and _49407_ (_17545_, _24496_, _24016_);
  and _49408_ (_17546_, _17545_, _23548_);
  not _49409_ (_17547_, _17545_);
  and _49410_ (_17548_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or _49411_ (_09331_, _17548_, _17546_);
  and _49412_ (_17549_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  and _49413_ (_17550_, _02513_, _24051_);
  or _49414_ (_09347_, _17550_, _17549_);
  and _49415_ (_17551_, _06208_, _24134_);
  and _49416_ (_17552_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _49417_ (_09357_, _17552_, _17551_);
  and _49418_ (_17553_, _06208_, _24051_);
  and _49419_ (_17554_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _49420_ (_09367_, _17554_, _17553_);
  and _49421_ (_17555_, _08559_, _23887_);
  and _49422_ (_17556_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or _49423_ (_09391_, _17556_, _17555_);
  and _49424_ (_17557_, _08559_, _23548_);
  and _49425_ (_17558_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or _49426_ (_09402_, _17558_, _17557_);
  and _49427_ (_17559_, _02996_, _23996_);
  and _49428_ (_17560_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  or _49429_ (_09412_, _17560_, _17559_);
  and _49430_ (_17561_, _08559_, _24219_);
  and _49431_ (_17562_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or _49432_ (_09416_, _17562_, _17561_);
  and _49433_ (_17563_, _17545_, _23887_);
  and _49434_ (_17564_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or _49435_ (_09427_, _17564_, _17563_);
  not _49436_ (_17565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _49437_ (_17566_, _02205_, _17565_);
  or _49438_ (_17567_, _02321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _49439_ (_17568_, _17567_, _08225_);
  nor _49440_ (_17569_, _17568_, _02219_);
  nor _49441_ (_17570_, _17569_, _02323_);
  nor _49442_ (_17571_, _17570_, _17566_);
  nor _49443_ (_17572_, _17571_, _01816_);
  and _49444_ (_09462_, _17572_, _01815_);
  and _49445_ (_17573_, _06208_, _23996_);
  and _49446_ (_17574_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _49447_ (_27221_, _17574_, _17573_);
  and _49448_ (_17575_, _12429_, _24134_);
  and _49449_ (_17576_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or _49450_ (_09513_, _17576_, _17575_);
  and _49451_ (_17577_, _08559_, _24051_);
  and _49452_ (_17578_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or _49453_ (_09544_, _17578_, _17577_);
  nor _49454_ (_26867_[6], _00069_, rst);
  and _49455_ (_17579_, _11311_, _24134_);
  and _49456_ (_17580_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or _49457_ (_09613_, _17580_, _17579_);
  and _49458_ (_17581_, _24301_, _22974_);
  and _49459_ (_17582_, _17581_, _23996_);
  not _49460_ (_17583_, _17581_);
  and _49461_ (_17584_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or _49462_ (_09630_, _17584_, _17582_);
  and _49463_ (_17585_, _03043_, _23887_);
  and _49464_ (_17586_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or _49465_ (_09649_, _17586_, _17585_);
  and _49466_ (_17587_, _03043_, _23548_);
  and _49467_ (_17588_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or _49468_ (_09662_, _17588_, _17587_);
  and _49469_ (_17589_, _17581_, _24134_);
  and _49470_ (_17590_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or _49471_ (_09664_, _17590_, _17589_);
  and _49472_ (_17591_, _03043_, _24219_);
  and _49473_ (_17592_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or _49474_ (_09666_, _17592_, _17591_);
  and _49475_ (_17593_, _08435_, _23548_);
  and _49476_ (_17594_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or _49477_ (_09686_, _17594_, _17593_);
  and _49478_ (_17595_, _15888_, _23887_);
  and _49479_ (_17596_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or _49480_ (_09688_, _17596_, _17595_);
  and _49481_ (_17597_, _15888_, _23548_);
  and _49482_ (_17598_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or _49483_ (_09691_, _17598_, _17597_);
  and _49484_ (_17599_, _15888_, _24089_);
  and _49485_ (_17600_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _49486_ (_09721_, _17600_, _17599_);
  and _49487_ (_17601_, _16121_, _24089_);
  and _49488_ (_17602_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _49489_ (_09735_, _17602_, _17601_);
  and _49490_ (_17603_, _24179_, _22867_);
  and _49491_ (_17604_, _17603_, _24174_);
  nand _49492_ (_17605_, _17604_, _24533_);
  and _49493_ (_17606_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _49494_ (_17607_, _15912_, _24178_);
  and _49495_ (_17608_, _17607_, _22869_);
  and _49496_ (_17609_, _17608_, _00747_);
  or _49497_ (_17610_, _17609_, _17606_);
  or _49498_ (_17611_, _17610_, _04433_);
  nand _49499_ (_17612_, _04433_, _01281_);
  and _49500_ (_17613_, _17612_, _22731_);
  and _49501_ (_09741_, _17613_, _17611_);
  and _49502_ (_17614_, _08559_, _24089_);
  and _49503_ (_17615_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or _49504_ (_09743_, _17615_, _17614_);
  and _49505_ (_17616_, _17391_, _24134_);
  and _49506_ (_17617_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or _49507_ (_26898_, _17617_, _17616_);
  and _49508_ (_17619_, _17110_, _24134_);
  and _49509_ (_17620_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or _49510_ (_09748_, _17620_, _17619_);
  and _49511_ (_17621_, _16529_, _23996_);
  and _49512_ (_17622_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _49513_ (_09755_, _17622_, _17621_);
  and _49514_ (_17623_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _49515_ (_17624_, _17608_, _00883_);
  or _49516_ (_17625_, _17624_, _17623_);
  or _49517_ (_17626_, _17625_, _04433_);
  not _49518_ (_17627_, _04433_);
  or _49519_ (_17628_, _17627_, _03853_);
  and _49520_ (_17629_, _17628_, _22731_);
  and _49521_ (_09766_, _17629_, _17626_);
  and _49522_ (_17630_, _17417_, _23548_);
  and _49523_ (_17631_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _49524_ (_09768_, _17631_, _17630_);
  and _49525_ (_17632_, _17102_, _23548_);
  and _49526_ (_17633_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _49527_ (_09770_, _17633_, _17632_);
  and _49528_ (_17634_, _17604_, _24562_);
  nor _49529_ (_17635_, _17634_, _04433_);
  or _49530_ (_17636_, _17635_, _26570_);
  not _49531_ (_17637_, _17635_);
  or _49532_ (_17638_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _49533_ (_17639_, _17638_, _22731_);
  and _49534_ (_09776_, _17639_, _17636_);
  not _49535_ (_17640_, _01520_);
  or _49536_ (_17641_, _17176_, _17640_);
  or _49537_ (_17642_, _17641_, _17171_);
  and _49538_ (_17643_, _01434_, _01384_);
  and _49539_ (_17644_, _01475_, _01424_);
  or _49540_ (_17645_, _01431_, _01387_);
  and _49541_ (_17646_, _17645_, _01488_);
  or _49542_ (_17647_, _17646_, _17644_);
  or _49543_ (_17648_, _17647_, _17643_);
  or _49544_ (_17649_, _01528_, _01492_);
  or _49545_ (_17650_, _17173_, _01522_);
  or _49546_ (_17651_, _17650_, _17649_);
  not _49547_ (_17652_, _01448_);
  nor _49548_ (_17653_, _01539_, _17652_);
  nand _49549_ (_17654_, _17653_, _01414_);
  or _49550_ (_17655_, _17654_, _17651_);
  or _49551_ (_17656_, _17655_, _17648_);
  or _49552_ (_17657_, _17656_, _17642_);
  and _49553_ (_17658_, _17657_, _22738_);
  nor _49554_ (_17659_, _17169_, _02002_);
  or _49555_ (_17660_, _17659_, rst);
  or _49556_ (_26843_[1], _17660_, _17658_);
  and _49557_ (_17661_, _16185_, _23887_);
  and _49558_ (_17662_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or _49559_ (_09788_, _17662_, _17661_);
  or _49560_ (_17663_, _17635_, _00569_);
  or _49561_ (_17664_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _49562_ (_17665_, _17664_, _22731_);
  and _49563_ (_09800_, _17665_, _17663_);
  and _49564_ (_17666_, _17102_, _23887_);
  and _49565_ (_17667_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _49566_ (_27292_, _17667_, _17666_);
  or _49567_ (_17668_, _24246_, _17165_);
  or _49568_ (_26842_[2], _17668_, _02008_);
  and _49569_ (_17669_, _24518_, _24051_);
  and _49570_ (_17670_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or _49571_ (_09807_, _17670_, _17669_);
  and _49572_ (_17671_, _17417_, _23887_);
  and _49573_ (_17672_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _49574_ (_09810_, _17672_, _17671_);
  and _49575_ (_17673_, _03269_, _23548_);
  and _49576_ (_17674_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  or _49577_ (_27166_, _17674_, _17673_);
  not _49578_ (_17675_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _49579_ (_17676_, _25481_, _17675_);
  or _49580_ (_17677_, _17676_, _25482_);
  and _49581_ (_17678_, _17677_, _00308_);
  and _49582_ (_17679_, _00312_, _23504_);
  and _49583_ (_17680_, _00311_, _17675_);
  or _49584_ (_17681_, _17680_, _00308_);
  or _49585_ (_17682_, _17681_, _17679_);
  nand _49586_ (_17683_, _17682_, _25684_);
  or _49587_ (_17684_, _17683_, _17678_);
  nand _49588_ (_17685_, _25683_, _23989_);
  and _49589_ (_17686_, _17685_, _22731_);
  and _49590_ (_09826_, _17686_, _17684_);
  and _49591_ (_17687_, _17417_, _24089_);
  and _49592_ (_17688_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _49593_ (_26899_, _17688_, _17687_);
  nand _49594_ (_17689_, _17637_, _00813_);
  or _49595_ (_17690_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _49596_ (_17691_, _17690_, _22731_);
  and _49597_ (_09835_, _17691_, _17689_);
  or _49598_ (_17692_, _17635_, _00473_);
  or _49599_ (_17693_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _49600_ (_17694_, _17693_, _22731_);
  and _49601_ (_09837_, _17694_, _17692_);
  and _49602_ (_17695_, _17102_, _23583_);
  and _49603_ (_17696_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _49604_ (_09844_, _17696_, _17695_);
  and _49605_ (_17697_, _24518_, _23996_);
  and _49606_ (_17698_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or _49607_ (_09846_, _17698_, _17697_);
  and _49608_ (_17699_, _17417_, _24134_);
  and _49609_ (_17700_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _49610_ (_09854_, _17700_, _17699_);
  and _49611_ (_17701_, _17102_, _24051_);
  and _49612_ (_17702_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _49613_ (_27293_, _17702_, _17701_);
  and _49614_ (_17703_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _49615_ (_17704_, _17608_, _00654_);
  or _49616_ (_17705_, _17704_, _17703_);
  or _49617_ (_17706_, _17705_, _04433_);
  nand _49618_ (_17707_, _04433_, _01192_);
  and _49619_ (_17708_, _17707_, _22731_);
  and _49620_ (_09864_, _17708_, _17706_);
  and _49621_ (_17709_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _49622_ (_17710_, _17608_, _00569_);
  or _49623_ (_17711_, _17710_, _17709_);
  or _49624_ (_17712_, _17711_, _04433_);
  nand _49625_ (_17713_, _04433_, _01121_);
  and _49626_ (_17714_, _17713_, _22731_);
  and _49627_ (_09875_, _17714_, _17712_);
  and _49628_ (_17715_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _49629_ (_17716_, _17608_, _00473_);
  or _49630_ (_17717_, _17716_, _17715_);
  or _49631_ (_17718_, _17717_, _04433_);
  nand _49632_ (_17719_, _04433_, _01061_);
  and _49633_ (_17720_, _17719_, _22731_);
  and _49634_ (_09881_, _17720_, _17718_);
  and _49635_ (_17721_, _24099_, _23996_);
  and _49636_ (_17722_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _49637_ (_09884_, _17722_, _17721_);
  and _49638_ (_17723_, _24057_, _24051_);
  and _49639_ (_17724_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or _49640_ (_09886_, _17724_, _17723_);
  and _49641_ (_17725_, _09670_, _23887_);
  and _49642_ (_17726_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or _49643_ (_09891_, _17726_, _17725_);
  and _49644_ (_17727_, _03269_, _23887_);
  and _49645_ (_17728_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  or _49646_ (_27167_, _17728_, _17727_);
  and _49647_ (_17729_, _09670_, _24219_);
  and _49648_ (_17730_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or _49649_ (_09896_, _17730_, _17729_);
  and _49650_ (_17731_, _17411_, _24219_);
  and _49651_ (_17732_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _49652_ (_26895_, _17732_, _17731_);
  and _49653_ (_17733_, _24134_, _24057_);
  and _49654_ (_17734_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or _49655_ (_09908_, _17734_, _17733_);
  or _49656_ (_17735_, _17635_, _00393_);
  or _49657_ (_17736_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _49658_ (_17737_, _17736_, _22731_);
  and _49659_ (_09911_, _17737_, _17735_);
  or _49660_ (_17738_, _17635_, _00747_);
  or _49661_ (_17739_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _49662_ (_17740_, _17739_, _22731_);
  and _49663_ (_09914_, _17740_, _17738_);
  or _49664_ (_17741_, _17635_, _00654_);
  or _49665_ (_17742_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _49666_ (_17743_, _17742_, _22731_);
  and _49667_ (_09916_, _17743_, _17741_);
  and _49668_ (_17744_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _49669_ (_17745_, _17608_, _00393_);
  or _49670_ (_17746_, _17745_, _17744_);
  or _49671_ (_17747_, _17746_, _04433_);
  nand _49672_ (_17748_, _04433_, _01009_);
  and _49673_ (_17749_, _17748_, _22731_);
  and _49674_ (_09918_, _17749_, _17747_);
  and _49675_ (_17750_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _49676_ (_17751_, _17608_, _26570_);
  or _49677_ (_17753_, _17751_, _17750_);
  or _49678_ (_17754_, _17753_, _04433_);
  or _49679_ (_17755_, _17627_, _00939_);
  and _49680_ (_17756_, _17755_, _22731_);
  and _49681_ (_09920_, _17756_, _17754_);
  and _49682_ (_17757_, _09670_, _24089_);
  and _49683_ (_17758_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or _49684_ (_27204_, _17758_, _17757_);
  and _49685_ (_17759_, _16004_, _23583_);
  and _49686_ (_17760_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  or _49687_ (_26967_, _17760_, _17759_);
  or _49688_ (_17761_, _17635_, _00883_);
  or _49689_ (_17762_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _49690_ (_17763_, _17762_, _22731_);
  and _49691_ (_09929_, _17763_, _17761_);
  and _49692_ (_17764_, _17411_, _23548_);
  and _49693_ (_17765_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _49694_ (_09939_, _17765_, _17764_);
  and _49695_ (_17766_, _16004_, _23887_);
  and _49696_ (_17767_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or _49697_ (_26966_, _17767_, _17766_);
  and _49698_ (_17769_, _25672_, _24219_);
  and _49699_ (_17770_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _49700_ (_27205_, _17770_, _17769_);
  and _49701_ (_17771_, _17078_, _23548_);
  and _49702_ (_17772_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _49703_ (_09950_, _17772_, _17771_);
  and _49704_ (_17773_, _17411_, _23887_);
  and _49705_ (_17774_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _49706_ (_09953_, _17774_, _17773_);
  nand _49707_ (_17775_, _16094_, _25951_);
  nor _49708_ (_17776_, _16099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _49709_ (_17777_, _17776_, _16100_);
  or _49710_ (_17778_, _17777_, _02616_);
  and _49711_ (_17779_, _17778_, _02295_);
  and _49712_ (_17780_, _17779_, _17775_);
  and _49713_ (_17781_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _49714_ (_09955_, _17781_, _17780_);
  nor _49715_ (_17782_, _17605_, _00813_);
  and _49716_ (_17783_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _49717_ (_17784_, _17783_, _04433_);
  or _49718_ (_17785_, _17784_, _17782_);
  nand _49719_ (_17786_, _04433_, _01353_);
  and _49720_ (_17787_, _17786_, _22731_);
  and _49721_ (_09959_, _17787_, _17785_);
  and _49722_ (_17788_, _17411_, _24089_);
  and _49723_ (_17789_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _49724_ (_09961_, _17789_, _17788_);
  and _49725_ (_17790_, _17078_, _23887_);
  and _49726_ (_17791_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _49727_ (_09966_, _17791_, _17790_);
  and _49728_ (_17792_, _02364_, _23887_);
  and _49729_ (_17793_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _49730_ (_27207_, _17793_, _17792_);
  and _49731_ (_17794_, _15581_, _24219_);
  and _49732_ (_17795_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or _49733_ (_09970_, _17795_, _17794_);
  and _49734_ (_17796_, _17411_, _24051_);
  and _49735_ (_17797_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _49736_ (_09972_, _17797_, _17796_);
  and _49737_ (_17798_, _17078_, _23583_);
  and _49738_ (_17799_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _49739_ (_09974_, _17799_, _17798_);
  and _49740_ (_17800_, _17581_, _24051_);
  and _49741_ (_17801_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or _49742_ (_09977_, _17801_, _17800_);
  and _49743_ (_17802_, _02364_, _23996_);
  and _49744_ (_17803_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _49745_ (_09980_, _17803_, _17802_);
  and _49746_ (_17804_, _16121_, _24051_);
  and _49747_ (_17805_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _49748_ (_09996_, _17805_, _17804_);
  and _49749_ (_17806_, _15581_, _24089_);
  and _49750_ (_17807_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or _49751_ (_10001_, _17807_, _17806_);
  and _49752_ (_17808_, _16004_, _24089_);
  and _49753_ (_17809_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or _49754_ (_10003_, _17809_, _17808_);
  and _49755_ (_17810_, _17411_, _23996_);
  and _49756_ (_17811_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _49757_ (_10006_, _17811_, _17810_);
  and _49758_ (_17812_, _17078_, _24051_);
  and _49759_ (_17813_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _49760_ (_10008_, _17813_, _17812_);
  and _49761_ (_17814_, _15581_, _23583_);
  and _49762_ (_17815_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or _49763_ (_27209_, _17815_, _17814_);
  and _49764_ (_17816_, _17078_, _23996_);
  and _49765_ (_17817_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _49766_ (_27286_, _17817_, _17816_);
  and _49767_ (_17819_, _17395_, _24219_);
  and _49768_ (_17820_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or _49769_ (_10018_, _17820_, _17819_);
  and _49770_ (_17821_, _16004_, _24134_);
  and _49771_ (_17822_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or _49772_ (_26968_, _17822_, _17821_);
  and _49773_ (_17823_, _17072_, _23548_);
  and _49774_ (_17824_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or _49775_ (_10040_, _17824_, _17823_);
  and _49776_ (_17825_, _02996_, _24089_);
  and _49777_ (_17826_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or _49778_ (_10043_, _17826_, _17825_);
  and _49779_ (_17827_, _17395_, _23583_);
  and _49780_ (_17828_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or _49781_ (_10045_, _17828_, _17827_);
  and _49782_ (_17829_, _08559_, _23583_);
  and _49783_ (_17830_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or _49784_ (_10048_, _17830_, _17829_);
  and _49785_ (_17831_, _16004_, _24051_);
  and _49786_ (_17832_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or _49787_ (_10050_, _17832_, _17831_);
  and _49788_ (_17833_, _17395_, _24051_);
  and _49789_ (_17834_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or _49790_ (_10055_, _17834_, _17833_);
  and _49791_ (_17835_, _24451_, _24219_);
  and _49792_ (_17836_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _49793_ (_10059_, _17836_, _17835_);
  and _49794_ (_17837_, _17072_, _23887_);
  and _49795_ (_17838_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or _49796_ (_10061_, _17838_, _17837_);
  and _49797_ (_17839_, _17072_, _24089_);
  and _49798_ (_17840_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or _49799_ (_10070_, _17840_, _17839_);
  and _49800_ (_17841_, _17395_, _24134_);
  and _49801_ (_17842_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or _49802_ (_26896_, _17842_, _17841_);
  and _49803_ (_17843_, _24451_, _23583_);
  and _49804_ (_17844_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _49805_ (_27212_, _17844_, _17843_);
  and _49806_ (_17845_, _03001_, _23583_);
  and _49807_ (_17846_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _49808_ (_27215_, _17846_, _17845_);
  and _49809_ (_17847_, _17072_, _24051_);
  and _49810_ (_17848_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or _49811_ (_27287_, _17848_, _17847_);
  and _49812_ (_17849_, _03269_, _23583_);
  and _49813_ (_17850_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  or _49814_ (_27168_, _17850_, _17849_);
  and _49815_ (_17851_, _03001_, _24219_);
  and _49816_ (_17852_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _49817_ (_27214_, _17852_, _17851_);
  and _49818_ (_17854_, _01810_, _23548_);
  and _49819_ (_17855_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or _49820_ (_10090_, _17855_, _17854_);
  and _49821_ (_17856_, _17391_, _24219_);
  and _49822_ (_17857_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or _49823_ (_10093_, _17857_, _17856_);
  and _49824_ (_17858_, _17072_, _23996_);
  and _49825_ (_17859_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or _49826_ (_27288_, _17859_, _17858_);
  and _49827_ (_17860_, _03001_, _23996_);
  and _49828_ (_17861_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _49829_ (_10097_, _17861_, _17860_);
  and _49830_ (_17862_, _00308_, _24636_);
  nand _49831_ (_17863_, _17862_, _23504_);
  or _49832_ (_17864_, _17862_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _49833_ (_17865_, _17864_, _25684_);
  and _49834_ (_17866_, _17865_, _17863_);
  or _49835_ (_17867_, _17866_, _25833_);
  and _49836_ (_10102_, _17867_, _22731_);
  and _49837_ (_17868_, _01810_, _23996_);
  and _49838_ (_17869_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or _49839_ (_10111_, _17869_, _17868_);
  and _49840_ (_17870_, _17391_, _23548_);
  and _49841_ (_17871_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or _49842_ (_10113_, _17871_, _17870_);
  and _49843_ (_17872_, _17110_, _24219_);
  and _49844_ (_17873_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or _49845_ (_10115_, _17873_, _17872_);
  and _49846_ (_17874_, _00308_, _24533_);
  nand _49847_ (_17875_, _17874_, _23504_);
  or _49848_ (_17876_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _49849_ (_17877_, _17876_, _25684_);
  and _49850_ (_17878_, _17877_, _17875_);
  or _49851_ (_17879_, _17878_, _25686_);
  and _49852_ (_10118_, _17879_, _22731_);
  and _49853_ (_17880_, _00308_, _24607_);
  nand _49854_ (_17881_, _17880_, _23504_);
  or _49855_ (_17882_, _17880_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _49856_ (_17883_, _17882_, _25684_);
  and _49857_ (_17884_, _17883_, _17881_);
  nor _49858_ (_17885_, _25684_, _24043_);
  or _49859_ (_17886_, _17885_, _17884_);
  and _49860_ (_10120_, _17886_, _22731_);
  and _49861_ (_17887_, _17110_, _23887_);
  and _49862_ (_17888_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or _49863_ (_10126_, _17888_, _17887_);
  or _49864_ (_17889_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _49865_ (_17890_, _23382_, _23380_);
  not _49866_ (_17891_, _23051_);
  nand _49867_ (_17892_, _23380_, _17891_);
  and _49868_ (_17893_, _17892_, _22995_);
  and _49869_ (_17894_, _17893_, _17890_);
  nand _49870_ (_17895_, _23427_, _23392_);
  or _49871_ (_17896_, _23427_, _23053_);
  and _49872_ (_17897_, _17896_, _23390_);
  and _49873_ (_17898_, _17897_, _17895_);
  and _49874_ (_17899_, _23528_, _23120_);
  and _49875_ (_17900_, _17899_, _23323_);
  and _49876_ (_17901_, _01104_, _26163_);
  and _49877_ (_17902_, _17901_, _01258_);
  nand _49878_ (_17903_, _17902_, _17900_);
  nand _49879_ (_17904_, _17903_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _49880_ (_17905_, _17904_, _17898_);
  nor _49881_ (_17906_, _17905_, _17894_);
  nand _49882_ (_17907_, _17906_, _00788_);
  or _49883_ (_17908_, _00364_, _26560_);
  or _49884_ (_17909_, _17908_, _00449_);
  or _49885_ (_17910_, _17909_, _00530_);
  or _49886_ (_17911_, _00715_, _00627_);
  or _49887_ (_17912_, _17911_, _17910_);
  and _49888_ (_17913_, _17912_, _23531_);
  or _49889_ (_17914_, _17913_, _17907_);
  or _49890_ (_17915_, _17914_, _00862_);
  and _49891_ (_17916_, _17915_, _17889_);
  or _49892_ (_17917_, _17916_, _00308_);
  and _49893_ (_17918_, _02578_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _49894_ (_17919_, _17918_, _02580_);
  or _49895_ (_17920_, _17919_, _00309_);
  and _49896_ (_17921_, _17920_, _17917_);
  or _49897_ (_17923_, _17921_, _25683_);
  or _49898_ (_17924_, _25684_, _23880_);
  and _49899_ (_17925_, _17924_, _22731_);
  and _49900_ (_10130_, _17925_, _17923_);
  and _49901_ (_17926_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _49902_ (_17927_, _17926_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _49903_ (_17928_, _23376_, _22995_);
  and _49904_ (_17929_, _23413_, _23390_);
  nand _49905_ (_17930_, _23484_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _49906_ (_17931_, _17930_, _17926_);
  or _49907_ (_17932_, _17931_, _17929_);
  or _49908_ (_17933_, _17932_, _17928_);
  and _49909_ (_17934_, _17933_, _17927_);
  or _49910_ (_17935_, _17934_, _00308_);
  or _49911_ (_17936_, _24594_, _00546_);
  nand _49912_ (_17937_, _17936_, _00308_);
  or _49913_ (_17938_, _17937_, _03798_);
  and _49914_ (_17939_, _17938_, _17935_);
  or _49915_ (_17940_, _17939_, _25683_);
  nand _49916_ (_17941_, _25683_, _24126_);
  and _49917_ (_17943_, _17941_, _22731_);
  and _49918_ (_10132_, _17943_, _17940_);
  and _49919_ (_17944_, _17391_, _23887_);
  and _49920_ (_17945_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or _49921_ (_26897_, _17945_, _17944_);
  and _49922_ (_17946_, _17110_, _23583_);
  and _49923_ (_17947_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or _49924_ (_10140_, _17947_, _17946_);
  and _49925_ (_17948_, _17391_, _23583_);
  and _49926_ (_17949_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or _49927_ (_10144_, _17949_, _17948_);
  and _49928_ (_10147_, _03857_, _22731_);
  and _49929_ (_17950_, _16008_, _23548_);
  and _49930_ (_17951_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or _49931_ (_10151_, _17951_, _17950_);
  and _49932_ (_17952_, _11441_, _24219_);
  and _49933_ (_17953_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or _49934_ (_10154_, _17953_, _17952_);
  and _49935_ (_17954_, _00308_, _24177_);
  nand _49936_ (_17955_, _17954_, _23504_);
  or _49937_ (_17957_, _17954_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _49938_ (_17958_, _17957_, _25684_);
  and _49939_ (_17959_, _17958_, _17955_);
  nor _49940_ (_17960_, _25684_, _23542_);
  or _49941_ (_17961_, _17960_, _17959_);
  and _49942_ (_10161_, _17961_, _22731_);
  and _49943_ (_17962_, _16731_, _24219_);
  and _49944_ (_17963_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or _49945_ (_27222_, _17963_, _17962_);
  and _49946_ (_17964_, _17385_, _24219_);
  and _49947_ (_17965_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or _49948_ (_10166_, _17965_, _17964_);
  and _49949_ (_17966_, _16008_, _24219_);
  and _49950_ (_17967_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  or _49951_ (_26960_, _17967_, _17966_);
  and _49952_ (_17968_, _17102_, _23996_);
  and _49953_ (_17969_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _49954_ (_27294_, _17969_, _17968_);
  and _49955_ (_17970_, _17385_, _23887_);
  and _49956_ (_17971_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or _49957_ (_10170_, _17971_, _17970_);
  and _49958_ (_17972_, _17066_, _24219_);
  and _49959_ (_17973_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _49960_ (_10173_, _17973_, _17972_);
  and _49961_ (_17974_, _03275_, _24051_);
  and _49962_ (_17975_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _49963_ (_10175_, _17975_, _17974_);
  and _49964_ (_17976_, _16731_, _23583_);
  and _49965_ (_17977_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or _49966_ (_10177_, _17977_, _17976_);
  and _49967_ (_17978_, _17385_, _24089_);
  and _49968_ (_17979_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or _49969_ (_10179_, _17979_, _17978_);
  and _49970_ (_17980_, _16541_, _23583_);
  and _49971_ (_17981_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or _49972_ (_10181_, _17981_, _17980_);
  and _49973_ (_17982_, _17066_, _23548_);
  and _49974_ (_17983_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _49975_ (_27295_, _17983_, _17982_);
  and _49976_ (_17984_, _16541_, _24219_);
  and _49977_ (_17985_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or _49978_ (_27224_, _17985_, _17984_);
  and _49979_ (_17986_, _17066_, _23583_);
  and _49980_ (_17987_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _49981_ (_10186_, _17987_, _17986_);
  and _49982_ (_17988_, _17385_, _24051_);
  and _49983_ (_17989_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or _49984_ (_26901_, _17989_, _17988_);
  and _49985_ (_17990_, _16541_, _24134_);
  and _49986_ (_17991_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or _49987_ (_10190_, _17991_, _17990_);
  and _49988_ (_17992_, _16008_, _24089_);
  and _49989_ (_17993_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or _49990_ (_10194_, _17993_, _17992_);
  and _49991_ (_17994_, _17066_, _24089_);
  and _49992_ (_17995_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _49993_ (_10196_, _17995_, _17994_);
  and _49994_ (_17996_, _07038_, _24134_);
  and _49995_ (_17997_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _49996_ (_10198_, _17997_, _17996_);
  and _49997_ (_17999_, _17379_, _23548_);
  and _49998_ (_18000_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _49999_ (_10201_, _18000_, _17999_);
  and _50000_ (_18001_, _04920_, _24089_);
  and _50001_ (_18002_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _50002_ (_10214_, _18002_, _18001_);
  nor _50003_ (_10220_, _03809_, rst);
  and _50004_ (_18003_, _17066_, _24051_);
  and _50005_ (_18004_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _50006_ (_10242_, _18004_, _18003_);
  and _50007_ (_18005_, _04920_, _23548_);
  and _50008_ (_18006_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _50009_ (_10244_, _18006_, _18005_);
  and _50010_ (_18007_, _16008_, _23583_);
  and _50011_ (_18008_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or _50012_ (_26961_, _18008_, _18007_);
  and _50013_ (_18009_, _17379_, _23583_);
  and _50014_ (_18010_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _50015_ (_26902_, _18010_, _18009_);
  and _50016_ (_18011_, _17066_, _23996_);
  and _50017_ (_18012_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _50018_ (_10260_, _18012_, _18011_);
  and _50019_ (_10266_, _03732_, _22731_);
  nor _50020_ (_10304_, _03721_, rst);
  and _50021_ (_10324_, _03792_, _22731_);
  and _50022_ (_18013_, _17379_, _24089_);
  and _50023_ (_18014_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _50024_ (_10337_, _18014_, _18013_);
  and _50025_ (_10358_, _03779_, _22731_);
  and _50026_ (_18015_, _02970_, _24089_);
  and _50027_ (_18016_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or _50028_ (_10366_, _18016_, _18015_);
  and _50029_ (_18017_, _03275_, _23996_);
  and _50030_ (_18018_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _50031_ (_27165_, _18018_, _18017_);
  and _50032_ (_18019_, _17379_, _23996_);
  and _50033_ (_18020_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _50034_ (_10375_, _18020_, _18019_);
  and _50035_ (_18021_, _17058_, _23548_);
  and _50036_ (_18022_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or _50037_ (_10379_, _18022_, _18021_);
  and _50038_ (_18023_, _16034_, _24089_);
  and _50039_ (_18024_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or _50040_ (_10420_, _18024_, _18023_);
  and _50041_ (_18025_, _17369_, _24219_);
  and _50042_ (_18026_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _50043_ (_10428_, _18026_, _18025_);
  and _50044_ (_18027_, _16066_, _23583_);
  and _50045_ (_18028_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or _50046_ (_10431_, _18028_, _18027_);
  and _50047_ (_18029_, _16066_, _24089_);
  and _50048_ (_18030_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or _50049_ (_10434_, _18030_, _18029_);
  nor _50050_ (_10442_, _03759_, rst);
  and _50051_ (_18031_, _17058_, _23887_);
  and _50052_ (_18032_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or _50053_ (_10446_, _18032_, _18031_);
  and _50054_ (_10454_, _03746_, _22731_);
  and _50055_ (_18033_, _17369_, _23887_);
  and _50056_ (_18034_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _50057_ (_10461_, _18034_, _18033_);
  and _50058_ (_18035_, _17058_, _24089_);
  and _50059_ (_18036_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or _50060_ (_27296_, _18036_, _18035_);
  and _50061_ (_18037_, _16704_, _24219_);
  and _50062_ (_18038_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _50063_ (_27234_, _18038_, _18037_);
  and _50064_ (_18039_, _16513_, _23548_);
  and _50065_ (_18040_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or _50066_ (_10506_, _18040_, _18039_);
  and _50067_ (_18041_, _17058_, _24134_);
  and _50068_ (_18042_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or _50069_ (_10508_, _18042_, _18041_);
  and _50070_ (_18043_, _16773_, _23887_);
  and _50071_ (_18044_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or _50072_ (_10513_, _18044_, _18043_);
  and _50073_ (_18045_, _17369_, _23583_);
  and _50074_ (_18046_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _50075_ (_10523_, _18046_, _18045_);
  and _50076_ (_18047_, _17369_, _24134_);
  and _50077_ (_18048_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _50078_ (_10528_, _18048_, _18047_);
  and _50079_ (_18049_, _17052_, _24219_);
  and _50080_ (_18050_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or _50081_ (_10534_, _18050_, _18049_);
  and _50082_ (_18051_, _16513_, _23583_);
  and _50083_ (_18052_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or _50084_ (_10539_, _18052_, _18051_);
  and _50085_ (_18053_, _16121_, _23887_);
  and _50086_ (_18054_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _50087_ (_10551_, _18054_, _18053_);
  and _50088_ (_18055_, _17369_, _23996_);
  and _50089_ (_18056_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _50090_ (_26905_, _18056_, _18055_);
  and _50091_ (_18057_, _03360_, _23548_);
  and _50092_ (_18058_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or _50093_ (_10560_, _18058_, _18057_);
  and _50094_ (_18059_, _17052_, _23548_);
  and _50095_ (_18060_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or _50096_ (_10562_, _18060_, _18059_);
  and _50097_ (_18061_, _16513_, _24051_);
  and _50098_ (_18062_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or _50099_ (_10569_, _18062_, _18061_);
  and _50100_ (_18063_, _17363_, _23548_);
  and _50101_ (_18064_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or _50102_ (_10572_, _18064_, _18063_);
  and _50103_ (_18065_, _16698_, _24051_);
  and _50104_ (_18066_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or _50105_ (_10574_, _18066_, _18065_);
  and _50106_ (_18067_, _16121_, _23548_);
  and _50107_ (_18068_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _50108_ (_10577_, _18068_, _18067_);
  and _50109_ (_18069_, _17052_, _23583_);
  and _50110_ (_18070_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or _50111_ (_10583_, _18070_, _18069_);
  and _50112_ (_18071_, _15888_, _23583_);
  and _50113_ (_18072_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or _50114_ (_10589_, _18072_, _18071_);
  and _50115_ (_18073_, _17052_, _24051_);
  and _50116_ (_18074_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or _50117_ (_27298_, _18074_, _18073_);
  and _50118_ (_18075_, _16513_, _24134_);
  and _50119_ (_18076_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or _50120_ (_26935_, _18076_, _18075_);
  and _50121_ (_18077_, _16698_, _24089_);
  and _50122_ (_18078_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or _50123_ (_10599_, _18078_, _18077_);
  and _50124_ (_18079_, _17363_, _23887_);
  and _50125_ (_18080_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or _50126_ (_10601_, _18080_, _18079_);
  and _50127_ (_18081_, _17046_, _24219_);
  and _50128_ (_18082_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _50129_ (_10607_, _18082_, _18081_);
  and _50130_ (_18083_, _09774_, _23887_);
  and _50131_ (_18084_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or _50132_ (_10609_, _18084_, _18083_);
  and _50133_ (_18085_, _16121_, _24219_);
  and _50134_ (_18086_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _50135_ (_10613_, _18086_, _18085_);
  and _50136_ (_18087_, _17363_, _24051_);
  and _50137_ (_18088_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or _50138_ (_10618_, _18088_, _18087_);
  and _50139_ (_18089_, _02617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _50140_ (_18090_, _02260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _50141_ (_18091_, _18090_, _02284_);
  and _50142_ (_18092_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _50143_ (_18093_, _18092_, _02263_);
  or _50144_ (_18094_, _18093_, _18091_);
  nor _50145_ (_18095_, _02248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _50146_ (_18096_, _18095_, _02615_);
  nand _50147_ (_18097_, _18096_, _18094_);
  nor _50148_ (_18098_, _18097_, _02616_);
  or _50149_ (_18099_, _18098_, _18089_);
  and _50150_ (_18100_, _18099_, _02295_);
  and _50151_ (_18101_, _02440_, _02450_);
  or _50152_ (_10620_, _18101_, _18100_);
  and _50153_ (_18102_, _11441_, _23887_);
  and _50154_ (_18103_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _50155_ (_10622_, _18103_, _18102_);
  and _50156_ (_18104_, _17363_, _23996_);
  and _50157_ (_18106_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or _50158_ (_10624_, _18106_, _18104_);
  and _50159_ (_18107_, _08578_, _24089_);
  and _50160_ (_18108_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or _50161_ (_10630_, _18108_, _18107_);
  and _50162_ (_18109_, _16494_, _23548_);
  and _50163_ (_18110_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or _50164_ (_10639_, _18110_, _18109_);
  and _50165_ (_18111_, _16494_, _23583_);
  and _50166_ (_18112_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or _50167_ (_26936_, _18112_, _18111_);
  and _50168_ (_18113_, _17046_, _23548_);
  and _50169_ (_18114_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _50170_ (_27299_, _18114_, _18113_);
  and _50171_ (_18115_, _17344_, _24219_);
  and _50172_ (_18116_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or _50173_ (_10645_, _18116_, _18115_);
  and _50174_ (_18117_, _16494_, _24051_);
  and _50175_ (_18118_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or _50176_ (_10648_, _18118_, _18117_);
  and _50177_ (_18120_, _06129_, _24134_);
  and _50178_ (_18121_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or _50179_ (_10650_, _18121_, _18120_);
  and _50180_ (_18122_, _03309_, _23996_);
  and _50181_ (_18123_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or _50182_ (_10653_, _18123_, _18122_);
  and _50183_ (_18124_, _17046_, _23583_);
  and _50184_ (_18125_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _50185_ (_10656_, _18125_, _18124_);
  and _50186_ (_18126_, _06129_, _23583_);
  and _50187_ (_18127_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or _50188_ (_10658_, _18127_, _18126_);
  and _50189_ (_18128_, _11441_, _23583_);
  and _50190_ (_18129_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or _50191_ (_10668_, _18129_, _18128_);
  and _50192_ (_18130_, _17046_, _24051_);
  and _50193_ (_18131_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _50194_ (_10671_, _18131_, _18130_);
  and _50195_ (_18132_, _25658_, _24089_);
  and _50196_ (_18133_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or _50197_ (_10675_, _18133_, _18132_);
  and _50198_ (_18135_, _17344_, _23548_);
  and _50199_ (_18136_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or _50200_ (_26906_, _18136_, _18135_);
  and _50201_ (_18137_, _25658_, _23548_);
  and _50202_ (_18138_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or _50203_ (_10681_, _18138_, _18137_);
  and _50204_ (_18139_, _17344_, _23583_);
  and _50205_ (_18140_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or _50206_ (_26908_, _18140_, _18139_);
  and _50207_ (_18141_, _24497_, _24089_);
  and _50208_ (_18142_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or _50209_ (_10686_, _18142_, _18141_);
  and _50210_ (_18143_, _17046_, _23996_);
  and _50211_ (_18144_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _50212_ (_10688_, _18144_, _18143_);
  and _50213_ (_18145_, _05485_, _23548_);
  and _50214_ (_18146_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _50215_ (_10690_, _18146_, _18145_);
  and _50216_ (_18147_, _16494_, _24134_);
  and _50217_ (_18148_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or _50218_ (_10692_, _18148_, _18147_);
  and _50219_ (_18149_, _16034_, _23996_);
  and _50220_ (_18150_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or _50221_ (_10694_, _18150_, _18149_);
  and _50222_ (_18151_, _17344_, _24089_);
  and _50223_ (_18152_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or _50224_ (_10696_, _18152_, _18151_);
  and _50225_ (_18153_, _17042_, _24219_);
  and _50226_ (_18154_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _50227_ (_27300_, _18154_, _18153_);
  and _50228_ (_18156_, _03275_, _23548_);
  and _50229_ (_18157_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _50230_ (_10703_, _18157_, _18156_);
  and _50231_ (_18158_, _03275_, _24219_);
  and _50232_ (_18159_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _50233_ (_10705_, _18159_, _18158_);
  and _50234_ (_18160_, _16698_, _23996_);
  and _50235_ (_18161_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or _50236_ (_10711_, _18161_, _18160_);
  and _50237_ (_18162_, _24497_, _23996_);
  and _50238_ (_18163_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or _50239_ (_10713_, _18163_, _18162_);
  and _50240_ (_18164_, _16698_, _24134_);
  and _50241_ (_18165_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or _50242_ (_10716_, _18165_, _18164_);
  and _50243_ (_18166_, _17344_, _24051_);
  and _50244_ (_18167_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or _50245_ (_26909_, _18167_, _18166_);
  and _50246_ (_18168_, _17042_, _23887_);
  and _50247_ (_18169_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _50248_ (_10720_, _18169_, _18168_);
  and _50249_ (_18170_, _16476_, _24219_);
  and _50250_ (_18171_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _50251_ (_10723_, _18171_, _18170_);
  and _50252_ (_18172_, _16476_, _23548_);
  and _50253_ (_18173_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _50254_ (_10734_, _18173_, _18172_);
  and _50255_ (_18174_, _08578_, _23583_);
  and _50256_ (_18175_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or _50257_ (_10736_, _18175_, _18174_);
  and _50258_ (_18177_, _16066_, _24134_);
  and _50259_ (_18178_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or _50260_ (_10739_, _18178_, _18177_);
  and _50261_ (_18179_, _17344_, _24134_);
  and _50262_ (_18180_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or _50263_ (_10747_, _18180_, _18179_);
  and _50264_ (_18181_, _17042_, _23583_);
  and _50265_ (_18182_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _50266_ (_27302_, _18182_, _18181_);
  and _50267_ (_18183_, _25124_, _25481_);
  nand _50268_ (_18184_, _18183_, _23504_);
  or _50269_ (_18185_, _18183_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _50270_ (_18186_, _18185_, _24539_);
  and _50271_ (_18187_, _18186_, _18184_);
  nand _50272_ (_18188_, _25130_, _23989_);
  or _50273_ (_18189_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _50274_ (_18190_, _18189_, _24179_);
  and _50275_ (_18191_, _18190_, _18188_);
  nor _50276_ (_18192_, _24178_, _04206_);
  or _50277_ (_18193_, _18192_, rst);
  or _50278_ (_18194_, _18193_, _18191_);
  or _50279_ (_10753_, _18194_, _18187_);
  and _50280_ (_18195_, _17042_, _24134_);
  and _50281_ (_18196_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _50282_ (_27303_, _18196_, _18195_);
  and _50283_ (_18197_, _16066_, _23996_);
  and _50284_ (_18198_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or _50285_ (_26959_, _18198_, _18197_);
  and _50286_ (_18199_, _17338_, _24219_);
  and _50287_ (_18200_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _50288_ (_26911_, _18200_, _18199_);
  and _50289_ (_18201_, _16476_, _23887_);
  and _50290_ (_18202_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _50291_ (_26938_, _18202_, _18201_);
  and _50292_ (_18203_, _16476_, _24089_);
  and _50293_ (_18204_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _50294_ (_26939_, _18204_, _18203_);
  and _50295_ (_18205_, _17338_, _23887_);
  and _50296_ (_18206_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _50297_ (_26912_, _18206_, _18205_);
  and _50298_ (_18207_, _11419_, _24089_);
  and _50299_ (_18208_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _50300_ (_27087_, _18208_, _18207_);
  and _50301_ (_18209_, _16476_, _24134_);
  and _50302_ (_18210_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _50303_ (_26940_, _18210_, _18209_);
  and _50304_ (_18211_, _17042_, _23996_);
  and _50305_ (_18212_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _50306_ (_27304_, _18212_, _18211_);
  and _50307_ (_18213_, _03043_, _23583_);
  and _50308_ (_18214_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or _50309_ (_27251_, _18214_, _18213_);
  and _50310_ (_18215_, _17338_, _24089_);
  and _50311_ (_18216_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _50312_ (_26914_, _18216_, _18215_);
  and _50313_ (_18217_, _17545_, _23583_);
  and _50314_ (_18218_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or _50315_ (_27254_, _18218_, _18217_);
  and _50316_ (_18219_, _17036_, _24219_);
  and _50317_ (_18220_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or _50318_ (_27305_, _18220_, _18219_);
  and _50319_ (_18221_, _17545_, _24219_);
  and _50320_ (_18222_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _50321_ (_27253_, _18222_, _18221_);
  and _50322_ (_18223_, _16476_, _23996_);
  and _50323_ (_18224_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _50324_ (_26941_, _18224_, _18223_);
  and _50325_ (_18225_, _17036_, _23887_);
  and _50326_ (_18226_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or _50327_ (_27306_, _18226_, _18225_);
  and _50328_ (_18227_, _16468_, _24219_);
  and _50329_ (_18228_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _50330_ (_26942_, _18228_, _18227_);
  and _50331_ (_18229_, _17338_, _24051_);
  and _50332_ (_18230_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _50333_ (_26915_, _18230_, _18229_);
  and _50334_ (_18231_, _16773_, _23996_);
  and _50335_ (_18232_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or _50336_ (_27239_, _18232_, _18231_);
  and _50337_ (_18233_, _11419_, _23583_);
  and _50338_ (_18234_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _50339_ (_27086_, _18234_, _18233_);
  and _50340_ (_18235_, _17338_, _23996_);
  and _50341_ (_18236_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _50342_ (_26916_, _18236_, _18235_);
  and _50343_ (_18237_, _17036_, _24089_);
  and _50344_ (_18238_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or _50345_ (_27307_, _18238_, _18237_);
  and _50346_ (_18239_, _16468_, _23548_);
  and _50347_ (_18240_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _50348_ (_26943_, _18240_, _18239_);
  and _50349_ (_18241_, _16773_, _24134_);
  and _50350_ (_18242_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or _50351_ (_27238_, _18242_, _18241_);
  and _50352_ (_18243_, _17334_, _24219_);
  and _50353_ (_18244_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _50354_ (_26918_, _18244_, _18243_);
  and _50355_ (_18245_, _11419_, _23887_);
  and _50356_ (_18246_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _50357_ (_27085_, _18246_, _18245_);
  and _50358_ (_18247_, _17036_, _24051_);
  and _50359_ (_18248_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or _50360_ (_27308_, _18248_, _18247_);
  and _50361_ (_18249_, _16468_, _23583_);
  and _50362_ (_18250_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _50363_ (_26944_, _18250_, _18249_);
  and _50364_ (_18251_, _17334_, _23887_);
  and _50365_ (_18252_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _50366_ (_26919_, _18252_, _18251_);
  and _50367_ (_18253_, _16773_, _24051_);
  and _50368_ (_18254_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or _50369_ (_27237_, _18254_, _18253_);
  and _50370_ (_18255_, _10867_, _23583_);
  and _50371_ (_18256_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or _50372_ (_27261_, _18256_, _18255_);
  and _50373_ (_18257_, _08578_, _23887_);
  and _50374_ (_18258_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or _50375_ (_27077_, _18258_, _18257_);
  and _50376_ (_18259_, _16468_, _24051_);
  and _50377_ (_18260_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _50378_ (_26945_, _18260_, _18259_);
  and _50379_ (_18261_, _03275_, _23583_);
  and _50380_ (_18262_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _50381_ (_10810_, _18262_, _18261_);
  and _50382_ (_18263_, _17036_, _24134_);
  and _50383_ (_18264_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or _50384_ (_10812_, _18264_, _18263_);
  and _50385_ (_18265_, _17334_, _23583_);
  and _50386_ (_18266_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _50387_ (_26920_, _18266_, _18265_);
  and _50388_ (_18268_, _02996_, _23548_);
  and _50389_ (_18269_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  or _50390_ (_10818_, _18269_, _18268_);
  and _50391_ (_18270_, _10867_, _24134_);
  and _50392_ (_18271_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or _50393_ (_10820_, _18271_, _18270_);
  and _50394_ (_18272_, _16468_, _24134_);
  and _50395_ (_18273_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _50396_ (_26946_, _18273_, _18272_);
  and _50397_ (_18274_, _16468_, _23996_);
  and _50398_ (_18275_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _50399_ (_10826_, _18275_, _18274_);
  and _50400_ (_18276_, _16014_, _24089_);
  and _50401_ (_18277_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or _50402_ (_10828_, _18277_, _18276_);
  and _50403_ (_18278_, _16014_, _24134_);
  and _50404_ (_18279_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or _50405_ (_10831_, _18279_, _18278_);
  and _50406_ (_18280_, _16773_, _24089_);
  and _50407_ (_18281_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or _50408_ (_10833_, _18281_, _18280_);
  and _50409_ (_18282_, _24394_, _24219_);
  and _50410_ (_18283_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _50411_ (_10838_, _18283_, _18282_);
  and _50412_ (_18284_, _25018_, _25481_);
  nand _50413_ (_18285_, _18284_, _23504_);
  or _50414_ (_18286_, _18284_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _50415_ (_18287_, _18286_, _24539_);
  and _50416_ (_18288_, _18287_, _18285_);
  nand _50417_ (_18289_, _25026_, _23989_);
  or _50418_ (_18290_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _50419_ (_18291_, _18290_, _24179_);
  and _50420_ (_18292_, _18291_, _18289_);
  nor _50421_ (_18293_, _24178_, _04146_);
  or _50422_ (_18294_, _18293_, rst);
  or _50423_ (_18295_, _18294_, _18292_);
  or _50424_ (_10842_, _18295_, _18288_);
  and _50425_ (_18296_, _11311_, _24051_);
  and _50426_ (_18297_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or _50427_ (_10844_, _18297_, _18296_);
  and _50428_ (_18298_, _05465_, _23548_);
  and _50429_ (_18299_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or _50430_ (_27067_, _18299_, _18298_);
  and _50431_ (_18300_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _50432_ (_18301_, _26724_, _22737_);
  or _50433_ (_18302_, _18301_, _18300_);
  or _50434_ (_18303_, _18302_, _02359_);
  and _50435_ (_26848_[2], _18303_, _22731_);
  and _50436_ (_18304_, _23890_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _50437_ (_18305_, _23784_, _23824_);
  or _50438_ (_18306_, _04793_, _04795_);
  or _50439_ (_18307_, _18306_, _18305_);
  or _50440_ (_18308_, _26703_, _23828_);
  or _50441_ (_18309_, _18308_, _17182_);
  or _50442_ (_18310_, _18309_, _18307_);
  or _50443_ (_18311_, _18310_, _11472_);
  and _50444_ (_18312_, _18311_, _23855_);
  or _50445_ (_26847_[1], _18312_, _18304_);
  and _50446_ (_18313_, _17581_, _23548_);
  and _50447_ (_18314_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or _50448_ (_10853_, _18314_, _18313_);
  or _50449_ (_18315_, _23724_, _26679_);
  or _50450_ (_18316_, _22736_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _50451_ (_18317_, _18316_, _22731_);
  and _50452_ (_26844_[7], _18317_, _18315_);
  and _50453_ (_18318_, _25220_, _25481_);
  nand _50454_ (_18319_, _18318_, _23504_);
  or _50455_ (_18320_, _18318_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _50456_ (_18321_, _18320_, _24539_);
  and _50457_ (_18322_, _18321_, _18319_);
  nand _50458_ (_18323_, _25228_, _23989_);
  or _50459_ (_18324_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _50460_ (_18325_, _18324_, _24179_);
  and _50461_ (_18326_, _18325_, _18323_);
  nor _50462_ (_18327_, _24178_, _04001_);
  or _50463_ (_18328_, _18327_, rst);
  or _50464_ (_18329_, _18328_, _18326_);
  or _50465_ (_10857_, _18329_, _18322_);
  and _50466_ (_18330_, _16014_, _24051_);
  and _50467_ (_18331_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _50468_ (_10864_, _18331_, _18330_);
  and _50469_ (_18332_, _10867_, _23996_);
  and _50470_ (_18333_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or _50471_ (_10866_, _18333_, _18332_);
  and _50472_ (_18334_, _25319_, _25481_);
  nand _50473_ (_18335_, _18334_, _23504_);
  or _50474_ (_18336_, _18334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _50475_ (_18337_, _18336_, _24539_);
  and _50476_ (_18338_, _18337_, _18335_);
  nand _50477_ (_18339_, _25327_, _23989_);
  or _50478_ (_18340_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _50479_ (_18341_, _18340_, _24179_);
  and _50480_ (_18342_, _18341_, _18339_);
  nor _50481_ (_18343_, _24178_, _03944_);
  or _50482_ (_18344_, _18343_, rst);
  or _50483_ (_18345_, _18344_, _18342_);
  or _50484_ (_10870_, _18345_, _18338_);
  and _50485_ (_18346_, _16698_, _24219_);
  and _50486_ (_18347_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or _50487_ (_10881_, _18347_, _18346_);
  and _50488_ (_18348_, _16698_, _23887_);
  and _50489_ (_18349_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or _50490_ (_10883_, _18349_, _18348_);
  and _50491_ (_18350_, _17581_, _24219_);
  and _50492_ (_18351_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or _50493_ (_27218_, _18351_, _18350_);
  and _50494_ (_18352_, _11419_, _24134_);
  and _50495_ (_18353_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _50496_ (_10886_, _18353_, _18352_);
  and _50497_ (_18354_, _16698_, _23548_);
  and _50498_ (_18355_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or _50499_ (_27240_, _18355_, _18354_);
  and _50500_ (_18356_, _11419_, _23996_);
  and _50501_ (_18357_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _50502_ (_10891_, _18357_, _18356_);
  and _50503_ (_18358_, _03281_, _24051_);
  and _50504_ (_18359_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or _50505_ (_10893_, _18359_, _18358_);
  and _50506_ (_18360_, _16670_, _23996_);
  and _50507_ (_18361_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or _50508_ (_10897_, _18361_, _18360_);
  and _50509_ (_18362_, _03360_, _23887_);
  and _50510_ (_18363_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or _50511_ (_10899_, _18363_, _18362_);
  and _50512_ (_18364_, _10867_, _24219_);
  and _50513_ (_18365_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or _50514_ (_10901_, _18365_, _18364_);
  and _50515_ (_18366_, _25414_, _23996_);
  and _50516_ (_18367_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _50517_ (_10910_, _18367_, _18366_);
  and _50518_ (_18368_, _03281_, _24089_);
  and _50519_ (_18369_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or _50520_ (_10915_, _18369_, _18368_);
  and _50521_ (_18370_, _08578_, _24051_);
  and _50522_ (_18371_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or _50523_ (_10918_, _18371_, _18370_);
  and _50524_ (_18372_, _16034_, _24134_);
  and _50525_ (_18373_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or _50526_ (_10921_, _18373_, _18372_);
  and _50527_ (_18374_, _16066_, _24219_);
  and _50528_ (_18375_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or _50529_ (_10923_, _18375_, _18374_);
  and _50530_ (_18376_, _08578_, _24134_);
  and _50531_ (_18377_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or _50532_ (_10925_, _18377_, _18376_);
  and _50533_ (_18378_, _02996_, _23887_);
  and _50534_ (_18379_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or _50535_ (_10928_, _18379_, _18378_);
  and _50536_ (_18380_, _24142_, _24089_);
  and _50537_ (_18381_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or _50538_ (_10933_, _18381_, _18380_);
  and _50539_ (_18382_, _25414_, _24134_);
  and _50540_ (_18383_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _50541_ (_10936_, _18383_, _18382_);
  and _50542_ (_18384_, _24089_, _22983_);
  and _50543_ (_18385_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or _50544_ (_10938_, _18385_, _18384_);
  and _50545_ (_18386_, _16704_, _23996_);
  and _50546_ (_18387_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or _50547_ (_10941_, _18387_, _18386_);
  and _50548_ (_18388_, _24099_, _23548_);
  and _50549_ (_18389_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _50550_ (_10942_, _18389_, _18388_);
  and _50551_ (_18390_, _24160_, _24051_);
  and _50552_ (_18391_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or _50553_ (_10944_, _18391_, _18390_);
  and _50554_ (_18392_, _24160_, _23583_);
  and _50555_ (_18393_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or _50556_ (_26922_, _18393_, _18392_);
  and _50557_ (_18394_, _17032_, _23996_);
  and _50558_ (_18395_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or _50559_ (_10946_, _18395_, _18394_);
  and _50560_ (_18396_, _24219_, _22983_);
  and _50561_ (_18397_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or _50562_ (_10948_, _18397_, _18396_);
  and _50563_ (_18398_, _16014_, _23996_);
  and _50564_ (_18399_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _50565_ (_26958_, _18399_, _18398_);
  and _50566_ (_18400_, _24320_, _23887_);
  and _50567_ (_18401_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _50568_ (_10950_, _18401_, _18400_);
  and _50569_ (_18402_, _24160_, _24089_);
  and _50570_ (_18403_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or _50571_ (_10951_, _18403_, _18402_);
  and _50572_ (_18404_, _24219_, _24099_);
  and _50573_ (_18405_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _50574_ (_10953_, _18405_, _18404_);
  and _50575_ (_18406_, _23996_, _22983_);
  and _50576_ (_18407_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or _50577_ (_10955_, _18407_, _18406_);
  and _50578_ (_18408_, _16704_, _24134_);
  and _50579_ (_18409_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _50580_ (_10958_, _18409_, _18408_);
  and _50581_ (_18410_, _24219_, _24147_);
  and _50582_ (_18411_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _50583_ (_10964_, _18411_, _18410_);
  and _50584_ (_18412_, _24142_, _23996_);
  and _50585_ (_18413_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or _50586_ (_10967_, _18413_, _18412_);
  and _50587_ (_18414_, _24057_, _23583_);
  and _50588_ (_18415_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or _50589_ (_10968_, _18415_, _18414_);
  and _50590_ (_18416_, _03309_, _23887_);
  and _50591_ (_18417_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or _50592_ (_10970_, _18417_, _18416_);
  and _50593_ (_18418_, _16704_, _24051_);
  and _50594_ (_18419_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _50595_ (_27235_, _18419_, _18418_);
  and _50596_ (_18420_, _25637_, _23887_);
  and _50597_ (_18421_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _50598_ (_10974_, _18421_, _18420_);
  and _50599_ (_18422_, _24099_, _24051_);
  and _50600_ (_18423_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _50601_ (_10976_, _18423_, _18422_);
  and _50602_ (_18424_, _24219_, _24142_);
  and _50603_ (_18425_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or _50604_ (_10978_, _18425_, _18424_);
  and _50605_ (_18426_, _24160_, _24134_);
  and _50606_ (_18427_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or _50607_ (_10980_, _18427_, _18426_);
  and _50608_ (_18428_, _03281_, _24134_);
  and _50609_ (_18429_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or _50610_ (_10982_, _18429_, _18428_);
  and _50611_ (_18430_, _24099_, _23887_);
  and _50612_ (_18431_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _50613_ (_10984_, _18431_, _18430_);
  and _50614_ (_18432_, _24320_, _24051_);
  and _50615_ (_18433_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _50616_ (_27279_, _18433_, _18432_);
  and _50617_ (_18434_, _24160_, _23996_);
  and _50618_ (_18435_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or _50619_ (_10993_, _18435_, _18434_);
  and _50620_ (_18436_, _24099_, _23583_);
  and _50621_ (_18437_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _50622_ (_10995_, _18437_, _18436_);
  and _50623_ (_18438_, _24224_, _24089_);
  and _50624_ (_18439_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _50625_ (_27283_, _18439_, _18438_);
  and _50626_ (_18440_, _10867_, _23548_);
  and _50627_ (_18442_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or _50628_ (_10999_, _18442_, _18440_);
  and _50629_ (_18443_, _05465_, _23996_);
  and _50630_ (_18444_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or _50631_ (_11001_, _18444_, _18443_);
  and _50632_ (_18445_, _24099_, _24089_);
  and _50633_ (_18446_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _50634_ (_11005_, _18446_, _18445_);
  and _50635_ (_26840_[1], _23660_, _22731_);
  and _50636_ (_18447_, _24147_, _24134_);
  and _50637_ (_18448_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _50638_ (_11011_, _18448_, _18447_);
  and _50639_ (_18449_, _10867_, _23887_);
  and _50640_ (_18450_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or _50641_ (_11014_, _18450_, _18449_);
  and _50642_ (_18451_, _24373_, _23996_);
  and _50643_ (_18452_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _50644_ (_11017_, _18452_, _18451_);
  and _50645_ (_18453_, _16014_, _24219_);
  and _50646_ (_18454_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _50647_ (_11021_, _18454_, _18453_);
  and _50648_ (_18455_, _17032_, _24089_);
  and _50649_ (_18456_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or _50650_ (_11023_, _18456_, _18455_);
  and _50651_ (_18457_, _17032_, _24134_);
  and _50652_ (_18458_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or _50653_ (_11024_, _18458_, _18457_);
  nand _50654_ (_18459_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _50655_ (_18460_, _18459_, _16094_);
  not _50656_ (_18461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _50657_ (_18462_, _06162_, _18461_);
  and _50658_ (_18463_, _06162_, _18461_);
  or _50659_ (_18464_, _18463_, _18462_);
  or _50660_ (_18465_, _18464_, _02617_);
  nand _50661_ (_18466_, _02617_, _18461_);
  and _50662_ (_18467_, _18466_, _18465_);
  or _50663_ (_18468_, _18467_, _18460_);
  and _50664_ (_18469_, _18468_, _02295_);
  and _50665_ (_18470_, _02440_, _02689_);
  or _50666_ (_11027_, _18470_, _18469_);
  and _50667_ (_18471_, _24219_, _24160_);
  and _50668_ (_18472_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or _50669_ (_26921_, _18472_, _18471_);
  and _50670_ (_18473_, _24160_, _23548_);
  and _50671_ (_18474_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or _50672_ (_11030_, _18474_, _18473_);
  and _50673_ (_18475_, _24155_, _24089_);
  and _50674_ (_18476_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or _50675_ (_11036_, _18476_, _18475_);
  and _50676_ (_18477_, _17032_, _24051_);
  and _50677_ (_18478_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or _50678_ (_11039_, _18478_, _18477_);
  and _50679_ (_18479_, _17334_, _24134_);
  and _50680_ (_18480_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _50681_ (_11042_, _18480_, _18479_);
  and _50682_ (_18481_, _17032_, _23887_);
  and _50683_ (_18482_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or _50684_ (_11043_, _18482_, _18481_);
  and _50685_ (_18483_, _24373_, _24134_);
  and _50686_ (_18484_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _50687_ (_11048_, _18484_, _18483_);
  and _50688_ (_18485_, _17334_, _23996_);
  and _50689_ (_18486_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _50690_ (_11050_, _18486_, _18485_);
  and _50691_ (_18487_, _17032_, _23583_);
  and _50692_ (_18488_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or _50693_ (_27309_, _18488_, _18487_);
  and _50694_ (_18489_, _24147_, _23583_);
  and _50695_ (_18490_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _50696_ (_11056_, _18490_, _18489_);
  and _50697_ (_18491_, _16014_, _23887_);
  and _50698_ (_18492_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or _50699_ (_26957_, _18492_, _18491_);
  and _50700_ (_18493_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and _50701_ (_18494_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _50702_ (_18495_, _18494_, _18493_);
  and _50703_ (_18496_, _18495_, _09792_);
  and _50704_ (_18497_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and _50705_ (_18498_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _50706_ (_18499_, _18498_, _18497_);
  and _50707_ (_18500_, _18499_, _05549_);
  or _50708_ (_18501_, _18500_, _18496_);
  or _50709_ (_18502_, _18501_, _09791_);
  and _50710_ (_18503_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and _50711_ (_18504_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _50712_ (_18505_, _18504_, _18503_);
  and _50713_ (_18506_, _18505_, _09792_);
  and _50714_ (_18507_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and _50715_ (_18508_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _50716_ (_18509_, _18508_, _18507_);
  and _50717_ (_18510_, _18509_, _05549_);
  or _50718_ (_18511_, _18510_, _18506_);
  or _50719_ (_18512_, _18511_, _05535_);
  and _50720_ (_18513_, _18512_, _09805_);
  and _50721_ (_18514_, _18513_, _18502_);
  or _50722_ (_18515_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _50723_ (_18516_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and _50724_ (_18517_, _18516_, _18515_);
  and _50725_ (_18518_, _18517_, _09792_);
  or _50726_ (_18519_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _50727_ (_18520_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and _50728_ (_18521_, _18520_, _18519_);
  and _50729_ (_18522_, _18521_, _05549_);
  or _50730_ (_18523_, _18522_, _18518_);
  or _50731_ (_18524_, _18523_, _09791_);
  or _50732_ (_18525_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _50733_ (_18526_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and _50734_ (_18527_, _18526_, _18525_);
  and _50735_ (_18528_, _18527_, _09792_);
  or _50736_ (_18529_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _50737_ (_18530_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and _50738_ (_18531_, _18530_, _18529_);
  and _50739_ (_18532_, _18531_, _05549_);
  or _50740_ (_18533_, _18532_, _18528_);
  or _50741_ (_18534_, _18533_, _05535_);
  and _50742_ (_18535_, _18534_, _05542_);
  and _50743_ (_18536_, _18535_, _18524_);
  or _50744_ (_18537_, _18536_, _18514_);
  and _50745_ (_18538_, _18537_, _05518_);
  and _50746_ (_18539_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and _50747_ (_18540_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _50748_ (_18541_, _18540_, _18539_);
  and _50749_ (_18542_, _18541_, _09792_);
  and _50750_ (_18543_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and _50751_ (_18544_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _50752_ (_18545_, _18544_, _18543_);
  and _50753_ (_18546_, _18545_, _05549_);
  or _50754_ (_18547_, _18546_, _18542_);
  or _50755_ (_18548_, _18547_, _09791_);
  and _50756_ (_18549_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and _50757_ (_18550_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _50758_ (_18551_, _18550_, _18549_);
  and _50759_ (_18552_, _18551_, _09792_);
  and _50760_ (_18553_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and _50761_ (_18554_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _50762_ (_18555_, _18554_, _18553_);
  and _50763_ (_18556_, _18555_, _05549_);
  or _50764_ (_18557_, _18556_, _18552_);
  or _50765_ (_18558_, _18557_, _05535_);
  and _50766_ (_18559_, _18558_, _09805_);
  and _50767_ (_18560_, _18559_, _18548_);
  or _50768_ (_18561_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _50769_ (_18562_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and _50770_ (_18563_, _18562_, _05549_);
  and _50771_ (_18564_, _18563_, _18561_);
  or _50772_ (_18565_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _50773_ (_18566_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and _50774_ (_18567_, _18566_, _09792_);
  and _50775_ (_18568_, _18567_, _18565_);
  or _50776_ (_18569_, _18568_, _18564_);
  or _50777_ (_18570_, _18569_, _09791_);
  or _50778_ (_18571_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _50779_ (_18572_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and _50780_ (_18573_, _18572_, _05549_);
  and _50781_ (_18574_, _18573_, _18571_);
  or _50782_ (_18575_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _50783_ (_18576_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and _50784_ (_18577_, _18576_, _09792_);
  and _50785_ (_18578_, _18577_, _18575_);
  or _50786_ (_18579_, _18578_, _18574_);
  or _50787_ (_18580_, _18579_, _05535_);
  and _50788_ (_18581_, _18580_, _05542_);
  and _50789_ (_18582_, _18581_, _18570_);
  or _50790_ (_18583_, _18582_, _18560_);
  and _50791_ (_18584_, _18583_, _09850_);
  or _50792_ (_18585_, _18584_, _18538_);
  and _50793_ (_18586_, _18585_, _09790_);
  and _50794_ (_18587_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and _50795_ (_18588_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _50796_ (_18589_, _18588_, _18587_);
  and _50797_ (_18590_, _18589_, _09792_);
  and _50798_ (_18591_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _50799_ (_18592_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _50800_ (_18593_, _18592_, _18591_);
  and _50801_ (_18594_, _18593_, _05549_);
  or _50802_ (_18595_, _18594_, _18590_);
  and _50803_ (_18596_, _18595_, _05535_);
  and _50804_ (_18597_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and _50805_ (_18598_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _50806_ (_18599_, _18598_, _18597_);
  and _50807_ (_18600_, _18599_, _09792_);
  and _50808_ (_18601_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _50809_ (_18602_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _50810_ (_18603_, _18602_, _18601_);
  and _50811_ (_18604_, _18603_, _05549_);
  or _50812_ (_18605_, _18604_, _18600_);
  and _50813_ (_18606_, _18605_, _09791_);
  or _50814_ (_18607_, _18606_, _18596_);
  and _50815_ (_18608_, _18607_, _09805_);
  or _50816_ (_18609_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _50817_ (_18610_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _50818_ (_18611_, _18610_, _05549_);
  and _50819_ (_18612_, _18611_, _18609_);
  or _50820_ (_18613_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _50821_ (_18614_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _50822_ (_18615_, _18614_, _09792_);
  and _50823_ (_18616_, _18615_, _18613_);
  or _50824_ (_18617_, _18616_, _18612_);
  and _50825_ (_18618_, _18617_, _05535_);
  or _50826_ (_18619_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _50827_ (_18620_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _50828_ (_18621_, _18620_, _05549_);
  and _50829_ (_18622_, _18621_, _18619_);
  or _50830_ (_18623_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _50831_ (_18624_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and _50832_ (_18625_, _18624_, _09792_);
  and _50833_ (_18626_, _18625_, _18623_);
  or _50834_ (_18627_, _18626_, _18622_);
  and _50835_ (_18628_, _18627_, _09791_);
  or _50836_ (_18629_, _18628_, _18618_);
  and _50837_ (_18630_, _18629_, _05542_);
  or _50838_ (_18631_, _18630_, _18608_);
  and _50839_ (_18632_, _18631_, _09850_);
  and _50840_ (_18633_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and _50841_ (_18634_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _50842_ (_18635_, _18634_, _18633_);
  and _50843_ (_18636_, _18635_, _09792_);
  and _50844_ (_18637_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and _50845_ (_18638_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _50846_ (_18639_, _18638_, _18637_);
  and _50847_ (_18640_, _18639_, _05549_);
  or _50848_ (_18641_, _18640_, _18636_);
  and _50849_ (_18642_, _18641_, _05535_);
  and _50850_ (_18643_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and _50851_ (_18644_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _50852_ (_18645_, _18644_, _18643_);
  and _50853_ (_18646_, _18645_, _09792_);
  and _50854_ (_18647_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and _50855_ (_18648_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _50856_ (_18649_, _18648_, _18647_);
  and _50857_ (_18650_, _18649_, _05549_);
  or _50858_ (_18651_, _18650_, _18646_);
  and _50859_ (_18652_, _18651_, _09791_);
  or _50860_ (_18653_, _18652_, _18642_);
  and _50861_ (_18654_, _18653_, _09805_);
  or _50862_ (_18655_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _50863_ (_18656_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and _50864_ (_18657_, _18656_, _18655_);
  and _50865_ (_18658_, _18657_, _09792_);
  or _50866_ (_18659_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _50867_ (_18660_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and _50868_ (_18661_, _18660_, _18659_);
  and _50869_ (_18662_, _18661_, _05549_);
  or _50870_ (_18663_, _18662_, _18658_);
  and _50871_ (_18664_, _18663_, _05535_);
  or _50872_ (_18665_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _50873_ (_18666_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and _50874_ (_18667_, _18666_, _18665_);
  and _50875_ (_18668_, _18667_, _09792_);
  or _50876_ (_18669_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _50877_ (_18670_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and _50878_ (_18671_, _18670_, _18669_);
  and _50879_ (_18672_, _18671_, _05549_);
  or _50880_ (_18673_, _18672_, _18668_);
  and _50881_ (_18674_, _18673_, _09791_);
  or _50882_ (_18675_, _18674_, _18664_);
  and _50883_ (_18676_, _18675_, _05542_);
  or _50884_ (_18677_, _18676_, _18654_);
  and _50885_ (_18678_, _18677_, _05518_);
  or _50886_ (_18679_, _18678_, _18632_);
  and _50887_ (_18680_, _18679_, _05520_);
  or _50888_ (_18681_, _18680_, _18586_);
  or _50889_ (_18682_, _18681_, _05526_);
  and _50890_ (_18683_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and _50891_ (_18684_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _50892_ (_18685_, _18684_, _18683_);
  and _50893_ (_18686_, _18685_, _09792_);
  and _50894_ (_18687_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and _50895_ (_18688_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _50896_ (_18689_, _18688_, _18687_);
  and _50897_ (_18690_, _18689_, _05549_);
  or _50898_ (_18691_, _18690_, _18686_);
  or _50899_ (_18692_, _18691_, _09791_);
  and _50900_ (_18693_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and _50901_ (_18694_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _50902_ (_18695_, _18694_, _18693_);
  and _50903_ (_18696_, _18695_, _09792_);
  and _50904_ (_18697_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and _50905_ (_18698_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _50906_ (_18699_, _18698_, _18697_);
  and _50907_ (_18700_, _18699_, _05549_);
  or _50908_ (_18701_, _18700_, _18696_);
  or _50909_ (_18702_, _18701_, _05535_);
  and _50910_ (_18703_, _18702_, _09805_);
  and _50911_ (_18704_, _18703_, _18692_);
  or _50912_ (_18705_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _50913_ (_18706_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and _50914_ (_18707_, _18706_, _05549_);
  and _50915_ (_18708_, _18707_, _18705_);
  or _50916_ (_18709_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _50917_ (_18710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and _50918_ (_18711_, _18710_, _09792_);
  and _50919_ (_18712_, _18711_, _18709_);
  or _50920_ (_18713_, _18712_, _18708_);
  or _50921_ (_18714_, _18713_, _09791_);
  or _50922_ (_18715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _50923_ (_18716_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and _50924_ (_18717_, _18716_, _05549_);
  and _50925_ (_18718_, _18717_, _18715_);
  or _50926_ (_18719_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _50927_ (_18720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and _50928_ (_18721_, _18720_, _09792_);
  and _50929_ (_18722_, _18721_, _18719_);
  or _50930_ (_18723_, _18722_, _18718_);
  or _50931_ (_18724_, _18723_, _05535_);
  and _50932_ (_18725_, _18724_, _05542_);
  and _50933_ (_18726_, _18725_, _18714_);
  or _50934_ (_18727_, _18726_, _18704_);
  and _50935_ (_18728_, _18727_, _09850_);
  and _50936_ (_18729_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and _50937_ (_18730_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _50938_ (_18731_, _18730_, _18729_);
  and _50939_ (_18732_, _18731_, _09792_);
  and _50940_ (_18733_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _50941_ (_18734_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _50942_ (_18735_, _18734_, _18733_);
  and _50943_ (_18736_, _18735_, _05549_);
  or _50944_ (_18737_, _18736_, _18732_);
  or _50945_ (_18738_, _18737_, _09791_);
  and _50946_ (_18739_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and _50947_ (_18740_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _50948_ (_18741_, _18740_, _18739_);
  and _50949_ (_18742_, _18741_, _09792_);
  and _50950_ (_18743_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _50951_ (_18744_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _50952_ (_18745_, _18744_, _18743_);
  and _50953_ (_18746_, _18745_, _05549_);
  or _50954_ (_18747_, _18746_, _18742_);
  or _50955_ (_18748_, _18747_, _05535_);
  and _50956_ (_18749_, _18748_, _09805_);
  and _50957_ (_18750_, _18749_, _18738_);
  or _50958_ (_18751_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _50959_ (_18752_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _50960_ (_18753_, _18752_, _18751_);
  and _50961_ (_18754_, _18753_, _09792_);
  or _50962_ (_18755_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _50963_ (_18756_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and _50964_ (_18757_, _18756_, _18755_);
  and _50965_ (_18758_, _18757_, _05549_);
  or _50966_ (_18759_, _18758_, _18754_);
  or _50967_ (_18760_, _18759_, _09791_);
  or _50968_ (_18761_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _50969_ (_18762_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and _50970_ (_18763_, _18762_, _18761_);
  and _50971_ (_18764_, _18763_, _09792_);
  or _50972_ (_18765_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _50973_ (_18766_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _50974_ (_18767_, _18766_, _18765_);
  and _50975_ (_18768_, _18767_, _05549_);
  or _50976_ (_18769_, _18768_, _18764_);
  or _50977_ (_18770_, _18769_, _05535_);
  and _50978_ (_18771_, _18770_, _05542_);
  and _50979_ (_18772_, _18771_, _18760_);
  or _50980_ (_18773_, _18772_, _18750_);
  and _50981_ (_18774_, _18773_, _05518_);
  or _50982_ (_18775_, _18774_, _18728_);
  and _50983_ (_18776_, _18775_, _09790_);
  or _50984_ (_18777_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _50985_ (_18778_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and _50986_ (_18779_, _18778_, _18777_);
  and _50987_ (_18780_, _18779_, _09792_);
  or _50988_ (_18781_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _50989_ (_18782_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and _50990_ (_18783_, _18782_, _18781_);
  and _50991_ (_18784_, _18783_, _05549_);
  or _50992_ (_18785_, _18784_, _18780_);
  and _50993_ (_18786_, _18785_, _09791_);
  or _50994_ (_18787_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _50995_ (_18788_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and _50996_ (_18789_, _18788_, _18787_);
  and _50997_ (_18790_, _18789_, _09792_);
  or _50998_ (_18791_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _50999_ (_18792_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and _51000_ (_18793_, _18792_, _18791_);
  and _51001_ (_18794_, _18793_, _05549_);
  or _51002_ (_18795_, _18794_, _18790_);
  and _51003_ (_18796_, _18795_, _05535_);
  or _51004_ (_18797_, _18796_, _18786_);
  and _51005_ (_18798_, _18797_, _05542_);
  and _51006_ (_18799_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and _51007_ (_18800_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _51008_ (_18801_, _18800_, _18799_);
  and _51009_ (_18802_, _18801_, _09792_);
  and _51010_ (_18803_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and _51011_ (_18804_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _51012_ (_18805_, _18804_, _18803_);
  and _51013_ (_18806_, _18805_, _05549_);
  or _51014_ (_18807_, _18806_, _18802_);
  and _51015_ (_18808_, _18807_, _09791_);
  and _51016_ (_18809_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and _51017_ (_18810_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _51018_ (_18811_, _18810_, _18809_);
  and _51019_ (_18812_, _18811_, _09792_);
  and _51020_ (_18813_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and _51021_ (_18814_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _51022_ (_18815_, _18814_, _18813_);
  and _51023_ (_18816_, _18815_, _05549_);
  or _51024_ (_18817_, _18816_, _18812_);
  and _51025_ (_18818_, _18817_, _05535_);
  or _51026_ (_18819_, _18818_, _18808_);
  and _51027_ (_18820_, _18819_, _09805_);
  or _51028_ (_18821_, _18820_, _18798_);
  and _51029_ (_18822_, _18821_, _05518_);
  or _51030_ (_18823_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _51031_ (_18824_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and _51032_ (_18825_, _18824_, _05549_);
  and _51033_ (_18826_, _18825_, _18823_);
  or _51034_ (_18827_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _51035_ (_18828_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and _51036_ (_18829_, _18828_, _09792_);
  and _51037_ (_18830_, _18829_, _18827_);
  or _51038_ (_18831_, _18830_, _18826_);
  and _51039_ (_18832_, _18831_, _09791_);
  or _51040_ (_18833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _51041_ (_18834_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and _51042_ (_18835_, _18834_, _05549_);
  and _51043_ (_18836_, _18835_, _18833_);
  or _51044_ (_18837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _51045_ (_18838_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and _51046_ (_18839_, _18838_, _09792_);
  and _51047_ (_18840_, _18839_, _18837_);
  or _51048_ (_18841_, _18840_, _18836_);
  and _51049_ (_18842_, _18841_, _05535_);
  or _51050_ (_18843_, _18842_, _18832_);
  and _51051_ (_18844_, _18843_, _05542_);
  and _51052_ (_18845_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and _51053_ (_18846_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _51054_ (_18847_, _18846_, _18845_);
  and _51055_ (_18848_, _18847_, _09792_);
  and _51056_ (_18849_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and _51057_ (_18850_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _51058_ (_18851_, _18850_, _18849_);
  and _51059_ (_18852_, _18851_, _05549_);
  or _51060_ (_18853_, _18852_, _18848_);
  and _51061_ (_18854_, _18853_, _09791_);
  and _51062_ (_18855_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and _51063_ (_18856_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _51064_ (_18857_, _18856_, _18855_);
  and _51065_ (_18858_, _18857_, _09792_);
  and _51066_ (_18859_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _51067_ (_18860_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _51068_ (_18861_, _18860_, _18859_);
  and _51069_ (_18862_, _18861_, _05549_);
  or _51070_ (_18863_, _18862_, _18858_);
  and _51071_ (_18864_, _18863_, _05535_);
  or _51072_ (_18865_, _18864_, _18854_);
  and _51073_ (_18866_, _18865_, _09805_);
  or _51074_ (_18867_, _18866_, _18844_);
  and _51075_ (_18868_, _18867_, _09850_);
  or _51076_ (_18869_, _18868_, _18822_);
  and _51077_ (_18870_, _18869_, _05520_);
  or _51078_ (_18871_, _18870_, _18776_);
  or _51079_ (_18872_, _18871_, _10033_);
  and _51080_ (_18873_, _18872_, _18682_);
  or _51081_ (_18874_, _18873_, _00143_);
  and _51082_ (_18875_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and _51083_ (_18876_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _51084_ (_18877_, _18876_, _18875_);
  and _51085_ (_18878_, _18877_, _09792_);
  and _51086_ (_18879_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and _51087_ (_18880_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _51088_ (_18881_, _18880_, _18879_);
  and _51089_ (_18882_, _18881_, _05549_);
  or _51090_ (_18883_, _18882_, _18878_);
  or _51091_ (_18884_, _18883_, _09791_);
  and _51092_ (_18885_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and _51093_ (_18886_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _51094_ (_18887_, _18886_, _18885_);
  and _51095_ (_18888_, _18887_, _09792_);
  and _51096_ (_18889_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and _51097_ (_18890_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _51098_ (_18891_, _18890_, _18889_);
  and _51099_ (_18892_, _18891_, _05549_);
  or _51100_ (_18893_, _18892_, _18888_);
  or _51101_ (_18894_, _18893_, _05535_);
  and _51102_ (_18895_, _18894_, _09805_);
  and _51103_ (_18896_, _18895_, _18884_);
  or _51104_ (_18897_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _51105_ (_18898_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and _51106_ (_18899_, _18898_, _18897_);
  and _51107_ (_18900_, _18899_, _09792_);
  or _51108_ (_18901_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _51109_ (_18902_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and _51110_ (_18903_, _18902_, _18901_);
  and _51111_ (_18904_, _18903_, _05549_);
  or _51112_ (_18905_, _18904_, _18900_);
  or _51113_ (_18906_, _18905_, _09791_);
  or _51114_ (_18907_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _51115_ (_18908_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and _51116_ (_18909_, _18908_, _18907_);
  and _51117_ (_18910_, _18909_, _09792_);
  or _51118_ (_18911_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _51119_ (_18912_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and _51120_ (_18913_, _18912_, _18911_);
  and _51121_ (_18914_, _18913_, _05549_);
  or _51122_ (_18915_, _18914_, _18910_);
  or _51123_ (_18916_, _18915_, _05535_);
  and _51124_ (_18917_, _18916_, _05542_);
  and _51125_ (_18918_, _18917_, _18906_);
  or _51126_ (_18919_, _18918_, _18896_);
  and _51127_ (_18920_, _18919_, _05518_);
  and _51128_ (_18921_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _51129_ (_18922_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _51130_ (_18923_, _18922_, _18921_);
  and _51131_ (_18924_, _18923_, _09792_);
  and _51132_ (_18925_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _51133_ (_18926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _51134_ (_18927_, _18926_, _18925_);
  and _51135_ (_18928_, _18927_, _05549_);
  or _51136_ (_18929_, _18928_, _18924_);
  or _51137_ (_18930_, _18929_, _09791_);
  and _51138_ (_18931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _51139_ (_18932_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or _51140_ (_18933_, _18932_, _18931_);
  and _51141_ (_18934_, _18933_, _09792_);
  and _51142_ (_18935_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _51143_ (_18936_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _51144_ (_18937_, _18936_, _18935_);
  and _51145_ (_18938_, _18937_, _05549_);
  or _51146_ (_18939_, _18938_, _18934_);
  or _51147_ (_18940_, _18939_, _05535_);
  and _51148_ (_18941_, _18940_, _09805_);
  and _51149_ (_18942_, _18941_, _18930_);
  or _51150_ (_18943_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or _51151_ (_18944_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _51152_ (_18945_, _18944_, _05549_);
  and _51153_ (_18946_, _18945_, _18943_);
  or _51154_ (_18947_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _51155_ (_18948_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _51156_ (_18949_, _18948_, _09792_);
  and _51157_ (_18951_, _18949_, _18947_);
  or _51158_ (_18952_, _18951_, _18946_);
  or _51159_ (_18953_, _18952_, _09791_);
  or _51160_ (_18954_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _51161_ (_18955_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _51162_ (_18956_, _18955_, _05549_);
  and _51163_ (_18957_, _18956_, _18954_);
  or _51164_ (_18958_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or _51165_ (_18959_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _51166_ (_18960_, _18959_, _09792_);
  and _51167_ (_18961_, _18960_, _18958_);
  or _51168_ (_18962_, _18961_, _18957_);
  or _51169_ (_18963_, _18962_, _05535_);
  and _51170_ (_18964_, _18963_, _05542_);
  and _51171_ (_18965_, _18964_, _18953_);
  or _51172_ (_18966_, _18965_, _18942_);
  and _51173_ (_18967_, _18966_, _09850_);
  or _51174_ (_18968_, _18967_, _18920_);
  and _51175_ (_18969_, _18968_, _09790_);
  and _51176_ (_18970_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _51177_ (_18971_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or _51178_ (_18972_, _18971_, _18970_);
  and _51179_ (_18973_, _18972_, _09792_);
  and _51180_ (_18974_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _51181_ (_18975_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _51182_ (_18976_, _18975_, _18974_);
  and _51183_ (_18977_, _18976_, _05549_);
  or _51184_ (_18978_, _18977_, _18973_);
  and _51185_ (_18979_, _18978_, _05535_);
  and _51186_ (_18980_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _51187_ (_18981_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or _51188_ (_18982_, _18981_, _18980_);
  and _51189_ (_18983_, _18982_, _09792_);
  and _51190_ (_18984_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _51191_ (_18985_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _51192_ (_18986_, _18985_, _18984_);
  and _51193_ (_18987_, _18986_, _05549_);
  or _51194_ (_18988_, _18987_, _18983_);
  and _51195_ (_18989_, _18988_, _09791_);
  or _51196_ (_18990_, _18989_, _18979_);
  and _51197_ (_18991_, _18990_, _09805_);
  or _51198_ (_18992_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _51199_ (_18993_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _51200_ (_18994_, _18993_, _05549_);
  and _51201_ (_18995_, _18994_, _18992_);
  or _51202_ (_18996_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or _51203_ (_18997_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _51204_ (_18998_, _18997_, _09792_);
  and _51205_ (_18999_, _18998_, _18996_);
  or _51206_ (_19000_, _18999_, _18995_);
  and _51207_ (_19001_, _19000_, _05535_);
  or _51208_ (_19002_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _51209_ (_19003_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _51210_ (_19004_, _19003_, _05549_);
  and _51211_ (_19005_, _19004_, _19002_);
  or _51212_ (_19006_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or _51213_ (_19007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _51214_ (_19008_, _19007_, _09792_);
  and _51215_ (_19009_, _19008_, _19006_);
  or _51216_ (_19010_, _19009_, _19005_);
  and _51217_ (_19011_, _19010_, _09791_);
  or _51218_ (_19012_, _19011_, _19001_);
  and _51219_ (_19013_, _19012_, _05542_);
  or _51220_ (_19014_, _19013_, _18991_);
  and _51221_ (_19015_, _19014_, _09850_);
  and _51222_ (_19016_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and _51223_ (_19017_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _51224_ (_19018_, _19017_, _19016_);
  and _51225_ (_19019_, _19018_, _09792_);
  and _51226_ (_19020_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and _51227_ (_19021_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _51228_ (_19022_, _19021_, _19020_);
  and _51229_ (_19023_, _19022_, _05549_);
  or _51230_ (_19024_, _19023_, _19019_);
  and _51231_ (_19025_, _19024_, _05535_);
  and _51232_ (_19026_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _51233_ (_19027_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _51234_ (_19028_, _19027_, _19026_);
  and _51235_ (_19029_, _19028_, _09792_);
  and _51236_ (_19030_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and _51237_ (_19031_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _51238_ (_19032_, _19031_, _19030_);
  and _51239_ (_19033_, _19032_, _05549_);
  or _51240_ (_19034_, _19033_, _19029_);
  and _51241_ (_19035_, _19034_, _09791_);
  or _51242_ (_19036_, _19035_, _19025_);
  and _51243_ (_19037_, _19036_, _09805_);
  or _51244_ (_19038_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _51245_ (_19039_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and _51246_ (_19040_, _19039_, _19038_);
  and _51247_ (_19041_, _19040_, _09792_);
  or _51248_ (_19042_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _51249_ (_19043_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and _51250_ (_19044_, _19043_, _19042_);
  and _51251_ (_19045_, _19044_, _05549_);
  or _51252_ (_19046_, _19045_, _19041_);
  and _51253_ (_19047_, _19046_, _05535_);
  or _51254_ (_19048_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _51255_ (_19049_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and _51256_ (_19050_, _19049_, _19048_);
  and _51257_ (_19051_, _19050_, _09792_);
  or _51258_ (_19052_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _51259_ (_19053_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _51260_ (_19054_, _19053_, _19052_);
  and _51261_ (_19055_, _19054_, _05549_);
  or _51262_ (_19056_, _19055_, _19051_);
  and _51263_ (_19057_, _19056_, _09791_);
  or _51264_ (_19058_, _19057_, _19047_);
  and _51265_ (_19059_, _19058_, _05542_);
  or _51266_ (_19060_, _19059_, _19037_);
  and _51267_ (_19061_, _19060_, _05518_);
  or _51268_ (_19062_, _19061_, _19015_);
  and _51269_ (_19063_, _19062_, _05520_);
  or _51270_ (_19064_, _19063_, _18969_);
  or _51271_ (_19065_, _19064_, _05526_);
  and _51272_ (_19066_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and _51273_ (_19067_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _51274_ (_19068_, _19067_, _19066_);
  and _51275_ (_19069_, _19068_, _09792_);
  and _51276_ (_19070_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and _51277_ (_19071_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _51278_ (_19072_, _19071_, _19070_);
  and _51279_ (_19073_, _19072_, _05549_);
  or _51280_ (_19074_, _19073_, _19069_);
  or _51281_ (_19075_, _19074_, _09791_);
  and _51282_ (_19076_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and _51283_ (_19077_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _51284_ (_19078_, _19077_, _19076_);
  and _51285_ (_19079_, _19078_, _09792_);
  and _51286_ (_19080_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and _51287_ (_19081_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _51288_ (_19082_, _19081_, _19080_);
  and _51289_ (_19083_, _19082_, _05549_);
  or _51290_ (_19084_, _19083_, _19079_);
  or _51291_ (_19085_, _19084_, _05535_);
  and _51292_ (_19086_, _19085_, _09805_);
  and _51293_ (_19087_, _19086_, _19075_);
  or _51294_ (_19088_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _51295_ (_19089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and _51296_ (_19090_, _19089_, _05549_);
  and _51297_ (_19091_, _19090_, _19088_);
  or _51298_ (_19092_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _51299_ (_19093_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and _51300_ (_19094_, _19093_, _09792_);
  and _51301_ (_19095_, _19094_, _19092_);
  or _51302_ (_19096_, _19095_, _19091_);
  or _51303_ (_19097_, _19096_, _09791_);
  or _51304_ (_19098_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _51305_ (_19099_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and _51306_ (_19100_, _19099_, _05549_);
  and _51307_ (_19101_, _19100_, _19098_);
  or _51308_ (_19102_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _51309_ (_19103_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and _51310_ (_19104_, _19103_, _09792_);
  and _51311_ (_19105_, _19104_, _19102_);
  or _51312_ (_19106_, _19105_, _19101_);
  or _51313_ (_19107_, _19106_, _05535_);
  and _51314_ (_19108_, _19107_, _05542_);
  and _51315_ (_19109_, _19108_, _19097_);
  or _51316_ (_19110_, _19109_, _19087_);
  and _51317_ (_19111_, _19110_, _09850_);
  and _51318_ (_19112_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _51319_ (_19113_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or _51320_ (_19114_, _19113_, _19112_);
  and _51321_ (_19115_, _19114_, _09792_);
  and _51322_ (_19116_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _51323_ (_19117_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _51324_ (_19118_, _19117_, _19116_);
  and _51325_ (_19119_, _19118_, _05549_);
  or _51326_ (_19120_, _19119_, _19115_);
  or _51327_ (_19121_, _19120_, _09791_);
  and _51328_ (_19122_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _51329_ (_19123_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or _51330_ (_19124_, _19123_, _19122_);
  and _51331_ (_19125_, _19124_, _09792_);
  and _51332_ (_19126_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _51333_ (_19127_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _51334_ (_19128_, _19127_, _19126_);
  and _51335_ (_19129_, _19128_, _05549_);
  or _51336_ (_19130_, _19129_, _19125_);
  or _51337_ (_19131_, _19130_, _05535_);
  and _51338_ (_19132_, _19131_, _09805_);
  and _51339_ (_19133_, _19132_, _19121_);
  or _51340_ (_19134_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or _51341_ (_19135_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _51342_ (_19136_, _19135_, _19134_);
  and _51343_ (_19137_, _19136_, _09792_);
  or _51344_ (_19138_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _51345_ (_19139_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _51346_ (_19140_, _19139_, _19138_);
  and _51347_ (_19141_, _19140_, _05549_);
  or _51348_ (_19142_, _19141_, _19137_);
  or _51349_ (_19143_, _19142_, _09791_);
  or _51350_ (_19144_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or _51351_ (_19145_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _51352_ (_19146_, _19145_, _19144_);
  and _51353_ (_19147_, _19146_, _09792_);
  or _51354_ (_19148_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _51355_ (_19149_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and _51356_ (_19150_, _19149_, _19148_);
  and _51357_ (_19151_, _19150_, _05549_);
  or _51358_ (_19152_, _19151_, _19147_);
  or _51359_ (_19153_, _19152_, _05535_);
  and _51360_ (_19154_, _19153_, _05542_);
  and _51361_ (_19155_, _19154_, _19143_);
  or _51362_ (_19156_, _19155_, _19133_);
  and _51363_ (_19157_, _19156_, _05518_);
  or _51364_ (_19158_, _19157_, _19111_);
  and _51365_ (_19159_, _19158_, _09790_);
  or _51366_ (_19160_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _51367_ (_19161_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _51368_ (_19162_, _19161_, _19160_);
  and _51369_ (_19163_, _19162_, _09792_);
  or _51370_ (_19164_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or _51371_ (_19165_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _51372_ (_19166_, _19165_, _19164_);
  and _51373_ (_19167_, _19166_, _05549_);
  or _51374_ (_19168_, _19167_, _19163_);
  and _51375_ (_19169_, _19168_, _09791_);
  or _51376_ (_19170_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _51377_ (_19171_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _51378_ (_19172_, _19171_, _19170_);
  and _51379_ (_19173_, _19172_, _09792_);
  or _51380_ (_19174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or _51381_ (_19175_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _51382_ (_19176_, _19175_, _19174_);
  and _51383_ (_19177_, _19176_, _05549_);
  or _51384_ (_19178_, _19177_, _19173_);
  and _51385_ (_19179_, _19178_, _05535_);
  or _51386_ (_19180_, _19179_, _19169_);
  and _51387_ (_19181_, _19180_, _05542_);
  and _51388_ (_19182_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _51389_ (_19183_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or _51390_ (_19184_, _19183_, _19182_);
  and _51391_ (_19185_, _19184_, _09792_);
  and _51392_ (_19186_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _51393_ (_19187_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _51394_ (_19188_, _19187_, _19186_);
  and _51395_ (_19189_, _19188_, _05549_);
  or _51396_ (_19190_, _19189_, _19185_);
  and _51397_ (_19191_, _19190_, _09791_);
  and _51398_ (_19192_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _51399_ (_19193_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _51400_ (_19194_, _19193_, _19192_);
  and _51401_ (_19195_, _19194_, _09792_);
  and _51402_ (_19196_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _51403_ (_19197_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or _51404_ (_19198_, _19197_, _19196_);
  and _51405_ (_19199_, _19198_, _05549_);
  or _51406_ (_19200_, _19199_, _19195_);
  and _51407_ (_19202_, _19200_, _05535_);
  or _51408_ (_19203_, _19202_, _19191_);
  and _51409_ (_19204_, _19203_, _09805_);
  or _51410_ (_19205_, _19204_, _19181_);
  and _51411_ (_19206_, _19205_, _05518_);
  or _51412_ (_19207_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or _51413_ (_19208_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and _51414_ (_19209_, _19208_, _05549_);
  and _51415_ (_19210_, _19209_, _19207_);
  or _51416_ (_19211_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or _51417_ (_19212_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and _51418_ (_19213_, _19212_, _09792_);
  and _51419_ (_19214_, _19213_, _19211_);
  or _51420_ (_19215_, _19214_, _19210_);
  and _51421_ (_19216_, _19215_, _09791_);
  or _51422_ (_19217_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or _51423_ (_19218_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and _51424_ (_19219_, _19218_, _05549_);
  and _51425_ (_19220_, _19219_, _19217_);
  or _51426_ (_19221_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or _51427_ (_19222_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and _51428_ (_19223_, _19222_, _09792_);
  and _51429_ (_19224_, _19223_, _19221_);
  or _51430_ (_19225_, _19224_, _19220_);
  and _51431_ (_19226_, _19225_, _05535_);
  or _51432_ (_19227_, _19226_, _19216_);
  and _51433_ (_19228_, _19227_, _05542_);
  and _51434_ (_19229_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and _51435_ (_19230_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or _51436_ (_19231_, _19230_, _19229_);
  and _51437_ (_19232_, _19231_, _09792_);
  and _51438_ (_19233_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and _51439_ (_19234_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or _51440_ (_19235_, _19234_, _19233_);
  and _51441_ (_19236_, _19235_, _05549_);
  or _51442_ (_19237_, _19236_, _19232_);
  and _51443_ (_19238_, _19237_, _09791_);
  and _51444_ (_19239_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and _51445_ (_19240_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or _51446_ (_19241_, _19240_, _19239_);
  and _51447_ (_19242_, _19241_, _09792_);
  and _51448_ (_19243_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and _51449_ (_19244_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or _51450_ (_19245_, _19244_, _19243_);
  and _51451_ (_19246_, _19245_, _05549_);
  or _51452_ (_19247_, _19246_, _19242_);
  and _51453_ (_19248_, _19247_, _05535_);
  or _51454_ (_19249_, _19248_, _19238_);
  and _51455_ (_19250_, _19249_, _09805_);
  or _51456_ (_19251_, _19250_, _19228_);
  and _51457_ (_19252_, _19251_, _09850_);
  or _51458_ (_19253_, _19252_, _19206_);
  and _51459_ (_19254_, _19253_, _05520_);
  or _51460_ (_19255_, _19254_, _19159_);
  or _51461_ (_19256_, _19255_, _10033_);
  and _51462_ (_19257_, _19256_, _19065_);
  or _51463_ (_19258_, _19257_, _04413_);
  and _51464_ (_19259_, _19258_, _18874_);
  or _51465_ (_19260_, _19259_, _05563_);
  or _51466_ (_19261_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _51467_ (_19262_, _19261_, _22731_);
  and _51468_ (_11068_, _19262_, _19260_);
  and _51469_ (_19263_, _16670_, _23887_);
  and _51470_ (_19264_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or _51471_ (_11071_, _19264_, _19263_);
  and _51472_ (_19265_, _03281_, _23887_);
  and _51473_ (_19266_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _51474_ (_27164_, _19266_, _19265_);
  and _51475_ (_19267_, _15996_, _23996_);
  and _51476_ (_19268_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or _51477_ (_11074_, _19268_, _19267_);
  and _51478_ (_19269_, _02065_, _24134_);
  and _51479_ (_19270_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or _51480_ (_11076_, _19270_, _19269_);
  and _51481_ (_19271_, _24367_, _24089_);
  and _51482_ (_19272_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or _51483_ (_11077_, _19272_, _19271_);
  and _51484_ (_19273_, _24367_, _23887_);
  and _51485_ (_19274_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or _51486_ (_11081_, _19274_, _19273_);
  and _51487_ (_19275_, _24952_, _24051_);
  and _51488_ (_19276_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _51489_ (_11085_, _19276_, _19275_);
  and _51490_ (_19277_, _24952_, _23583_);
  and _51491_ (_19278_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _51492_ (_11088_, _19278_, _19277_);
  and _51493_ (_19279_, _24900_, _23996_);
  and _51494_ (_19280_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _51495_ (_11091_, _19280_, _19279_);
  and _51496_ (_19281_, _16670_, _23548_);
  and _51497_ (_19282_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or _51498_ (_27257_, _19282_, _19281_);
  and _51499_ (_19283_, _24900_, _23887_);
  and _51500_ (_19284_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _51501_ (_11103_, _19284_, _19283_);
  and _51502_ (_19285_, _02065_, _24051_);
  and _51503_ (_19286_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or _51504_ (_27084_, _19286_, _19285_);
  and _51505_ (_19287_, _24832_, _23583_);
  and _51506_ (_19288_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or _51507_ (_11106_, _19288_, _19287_);
  and _51508_ (_19289_, _24813_, _23583_);
  and _51509_ (_19290_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _51510_ (_11109_, _19290_, _19289_);
  and _51511_ (_19291_, _03281_, _23548_);
  and _51512_ (_19292_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or _51513_ (_11111_, _19292_, _19291_);
  and _51514_ (_19293_, _24735_, _24089_);
  and _51515_ (_19294_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or _51516_ (_11113_, _19294_, _19293_);
  and _51517_ (_19295_, _24735_, _23548_);
  and _51518_ (_19296_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or _51519_ (_11115_, _19296_, _19295_);
  and _51520_ (_19297_, _24694_, _24134_);
  and _51521_ (_19298_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or _51522_ (_11117_, _19298_, _19297_);
  and _51523_ (_19299_, _24694_, _23887_);
  and _51524_ (_19300_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or _51525_ (_11121_, _19300_, _19299_);
  and _51526_ (_19301_, _24503_, _23996_);
  and _51527_ (_19302_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _51528_ (_27195_, _19302_, _19301_);
  and _51529_ (_19303_, _05431_, _24134_);
  and _51530_ (_19304_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or _51531_ (_27131_, _19304_, _19303_);
  and _51532_ (_19305_, _16773_, _23548_);
  and _51533_ (_19306_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or _51534_ (_27236_, _19306_, _19305_);
  and _51535_ (_19307_, _16670_, _24051_);
  and _51536_ (_19308_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or _51537_ (_11124_, _19308_, _19307_);
  and _51538_ (_19309_, _24490_, _23548_);
  and _51539_ (_19310_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _51540_ (_11126_, _19310_, _19309_);
  and _51541_ (_19311_, _24602_, _23996_);
  and _51542_ (_19312_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or _51543_ (_11128_, _19312_, _19311_);
  and _51544_ (_19313_, _02065_, _24089_);
  and _51545_ (_19314_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or _51546_ (_11133_, _19314_, _19313_);
  and _51547_ (_19315_, _24602_, _23887_);
  and _51548_ (_19316_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or _51549_ (_11135_, _19316_, _19315_);
  and _51550_ (_19317_, _16072_, _24089_);
  and _51551_ (_19318_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or _51552_ (_11142_, _19318_, _19317_);
  and _51553_ (_19319_, _16670_, _24089_);
  and _51554_ (_19320_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or _51555_ (_11144_, _19320_, _19319_);
  and _51556_ (_19321_, _24525_, _23548_);
  and _51557_ (_19322_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or _51558_ (_11146_, _19322_, _19321_);
  and _51559_ (_19323_, _24510_, _24134_);
  and _51560_ (_19324_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _51561_ (_27192_, _19324_, _19323_);
  and _51562_ (_19325_, _16670_, _23583_);
  and _51563_ (_19326_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or _51564_ (_11156_, _19326_, _19325_);
  and _51565_ (_19327_, _16072_, _23583_);
  and _51566_ (_19328_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or _51567_ (_11162_, _19328_, _19327_);
  and _51568_ (_19329_, _24503_, _23583_);
  and _51569_ (_19330_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _51570_ (_11167_, _19330_, _19329_);
  and _51571_ (_19331_, _17581_, _23887_);
  and _51572_ (_19332_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or _51573_ (_11170_, _19332_, _19331_);
  and _51574_ (_19333_, _24490_, _23996_);
  and _51575_ (_19334_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _51576_ (_11172_, _19334_, _19333_);
  and _51577_ (_19335_, _24155_, _24134_);
  and _51578_ (_19336_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or _51579_ (_11173_, _19336_, _19335_);
  and _51580_ (_19337_, _24952_, _23996_);
  and _51581_ (_19338_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _51582_ (_11176_, _19338_, _19337_);
  and _51583_ (_19339_, _24900_, _24089_);
  and _51584_ (_19340_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _51585_ (_11178_, _19340_, _19339_);
  and _51586_ (_19341_, _24900_, _24219_);
  and _51587_ (_19342_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _51588_ (_11180_, _19342_, _19341_);
  and _51589_ (_19343_, _24302_, _24219_);
  and _51590_ (_19344_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or _51591_ (_27230_, _19344_, _19343_);
  and _51592_ (_19345_, _24832_, _24051_);
  and _51593_ (_19346_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or _51594_ (_27199_, _19346_, _19345_);
  and _51595_ (_19347_, _24832_, _24219_);
  and _51596_ (_19348_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or _51597_ (_27197_, _19348_, _19347_);
  and _51598_ (_19349_, _24813_, _24051_);
  and _51599_ (_19350_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _51600_ (_11188_, _19350_, _19349_);
  and _51601_ (_19351_, _24813_, _23548_);
  and _51602_ (_19352_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _51603_ (_11190_, _19352_, _19351_);
  and _51604_ (_19353_, _24735_, _24134_);
  and _51605_ (_19354_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or _51606_ (_11192_, _19354_, _19353_);
  and _51607_ (_19355_, _17581_, _24089_);
  and _51608_ (_19356_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or _51609_ (_11197_, _19356_, _19355_);
  and _51610_ (_19357_, _03281_, _23583_);
  and _51611_ (_19358_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or _51612_ (_11199_, _19358_, _19357_);
  and _51613_ (_19359_, _24490_, _23583_);
  and _51614_ (_19360_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _51615_ (_11200_, _19360_, _19359_);
  and _51616_ (_19361_, _24602_, _24089_);
  and _51617_ (_19362_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or _51618_ (_11202_, _19362_, _19361_);
  and _51619_ (_19363_, _24602_, _24219_);
  and _51620_ (_19364_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or _51621_ (_11204_, _19364_, _19363_);
  and _51622_ (_19365_, _24525_, _24051_);
  and _51623_ (_19366_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or _51624_ (_27193_, _19366_, _19365_);
  and _51625_ (_19367_, _24503_, _24219_);
  and _51626_ (_19368_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _51627_ (_11213_, _19368_, _19367_);
  and _51628_ (_19369_, _24367_, _24134_);
  and _51629_ (_19370_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or _51630_ (_11215_, _19370_, _19369_);
  and _51631_ (_19371_, _16678_, _24051_);
  and _51632_ (_19372_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or _51633_ (_11220_, _19372_, _19371_);
  and _51634_ (_19373_, _24735_, _23887_);
  and _51635_ (_19374_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or _51636_ (_11222_, _19374_, _19373_);
  and _51637_ (_19375_, _24694_, _23583_);
  and _51638_ (_19376_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or _51639_ (_11224_, _19376_, _19375_);
  and _51640_ (_19377_, _16773_, _24219_);
  and _51641_ (_19378_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or _51642_ (_11228_, _19378_, _19377_);
  and _51643_ (_19379_, _24525_, _23887_);
  and _51644_ (_19380_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or _51645_ (_11232_, _19380_, _19379_);
  and _51646_ (_19381_, _24503_, _24089_);
  and _51647_ (_19382_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _51648_ (_11234_, _19382_, _19381_);
  and _51649_ (_19383_, _24952_, _24219_);
  and _51650_ (_19384_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _51651_ (_11237_, _19384_, _19383_);
  and _51652_ (_19385_, _24832_, _23548_);
  and _51653_ (_19386_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or _51654_ (_11240_, _19386_, _19385_);
  and _51655_ (_19387_, _16678_, _24089_);
  and _51656_ (_19388_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _51657_ (_11242_, _19388_, _19387_);
  and _51658_ (_19389_, _16678_, _23583_);
  and _51659_ (_19390_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or _51660_ (_27256_, _19390_, _19389_);
  and _51661_ (_19391_, _25210_, _23996_);
  and _51662_ (_19392_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or _51663_ (_27156_, _19392_, _19391_);
  and _51664_ (_19393_, _16072_, _24134_);
  and _51665_ (_19394_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or _51666_ (_11249_, _19394_, _19393_);
  and _51667_ (_19395_, _24840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _51668_ (_19396_, _24750_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _51669_ (_19397_, _24750_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _51670_ (_19398_, _19397_, _19396_);
  nor _51671_ (_19399_, _19398_, _24781_);
  or _51672_ (_19400_, _19399_, _24747_);
  or _51673_ (_19401_, _19400_, _19395_);
  or _51674_ (_19402_, _19398_, _24844_);
  and _51675_ (_19403_, _19402_, _22731_);
  and _51676_ (_11258_, _19403_, _19401_);
  and _51677_ (_19404_, _16072_, _24051_);
  and _51678_ (_19405_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  or _51679_ (_11262_, _19405_, _19404_);
  or _51680_ (_19406_, _24913_, _24851_);
  and _51681_ (_19407_, _19406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _51682_ (_19408_, _19407_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor _51683_ (_19409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _24750_);
  not _51684_ (_19410_, _19409_);
  nor _51685_ (_19411_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _51686_ (_19412_, _19411_, _24749_);
  and _51687_ (_19413_, _19412_, _19410_);
  nor _51688_ (_19414_, _02137_, _02113_);
  nor _51689_ (_19415_, _19414_, _24749_);
  nor _51690_ (_19416_, _19415_, _19413_);
  and _51691_ (_19417_, _19416_, _19408_);
  or _51692_ (_19418_, _19417_, _04091_);
  and _51693_ (_19419_, _19418_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _51694_ (_19420_, _24174_, _24187_);
  nor _51695_ (_19421_, _24540_, _19420_);
  or _51696_ (_19422_, _19421_, _19419_);
  nand _51697_ (_19423_, _19421_, _24531_);
  and _51698_ (_19424_, _19423_, _19422_);
  nand _51699_ (_19425_, _19424_, _24704_);
  nand _51700_ (_19426_, _24703_, _23542_);
  and _51701_ (_19427_, _19426_, _22731_);
  and _51702_ (_11268_, _19427_, _19425_);
  and _51703_ (_11283_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _22731_);
  and _51704_ (_19428_, _02232_, _24089_);
  and _51705_ (_19429_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or _51706_ (_11285_, _19429_, _19428_);
  and _51707_ (_19430_, _02498_, _23548_);
  and _51708_ (_19431_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _51709_ (_11287_, _19431_, _19430_);
  and _51710_ (_19432_, _02882_, _23583_);
  and _51711_ (_19433_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _51712_ (_11289_, _19433_, _19432_);
  and _51713_ (_19434_, _02980_, _24134_);
  and _51714_ (_19435_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _51715_ (_26972_, _19435_, _19434_);
  and _51716_ (_19436_, _02980_, _23548_);
  and _51717_ (_19437_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _51718_ (_26970_, _19437_, _19436_);
  and _51719_ (_19438_, _03020_, _23583_);
  and _51720_ (_19439_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or _51721_ (_11292_, _19439_, _19438_);
  and _51722_ (_19440_, _03180_, _24134_);
  and _51723_ (_19441_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _51724_ (_11294_, _19441_, _19440_);
  and _51725_ (_19442_, _03217_, _24219_);
  and _51726_ (_19443_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _51727_ (_11296_, _19443_, _19442_);
  and _51728_ (_19444_, _03343_, _24134_);
  and _51729_ (_19445_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _51730_ (_11298_, _19445_, _19444_);
  and _51731_ (_19446_, _04608_, _24051_);
  and _51732_ (_19447_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _51733_ (_11300_, _19447_, _19446_);
  and _51734_ (_19448_, _16678_, _23996_);
  and _51735_ (_19449_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _51736_ (_11303_, _19449_, _19448_);
  and _51737_ (_19450_, _17581_, _23583_);
  and _51738_ (_19451_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or _51739_ (_11305_, _19451_, _19450_);
  not _51740_ (_19452_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _51741_ (_19453_, _19407_, _19452_);
  nand _51742_ (_19454_, _19414_, _19413_);
  or _51743_ (_19455_, _19454_, _19453_);
  and _51744_ (_19456_, _19455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _51745_ (_19457_, _19456_, _04687_);
  and _51746_ (_19458_, _24541_, _24174_);
  and _51747_ (_19459_, _19458_, _25481_);
  or _51748_ (_19460_, _19459_, _19457_);
  nand _51749_ (_19461_, _19459_, _23504_);
  and _51750_ (_19462_, _19461_, _19460_);
  or _51751_ (_19463_, _19462_, _24703_);
  nand _51752_ (_19464_, _24703_, _23989_);
  and _51753_ (_19465_, _19464_, _22731_);
  and _51754_ (_11310_, _19465_, _19463_);
  and _51755_ (_19466_, _04950_, _24134_);
  and _51756_ (_19467_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  or _51757_ (_27163_, _19467_, _19466_);
  and _51758_ (_11315_, _26285_, _22731_);
  and _51759_ (_19468_, _16072_, _24219_);
  and _51760_ (_19469_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or _51761_ (_26953_, _19469_, _19468_);
  nand _51762_ (_19470_, _22886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _51763_ (_19471_, _19470_, _24593_);
  or _51764_ (_19472_, _19471_, _03798_);
  and _51765_ (_19473_, _19472_, _24699_);
  nand _51766_ (_19474_, _24699_, _22886_);
  and _51767_ (_19475_, _19474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _51768_ (_19476_, _19475_, _24703_);
  or _51769_ (_19477_, _19476_, _19473_);
  nand _51770_ (_19478_, _24703_, _24126_);
  and _51771_ (_19479_, _19478_, _22731_);
  and _51772_ (_11322_, _19479_, _19477_);
  and _51773_ (_19480_, _24089_, _23946_);
  and _51774_ (_19481_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or _51775_ (_11326_, _19481_, _19480_);
  and _51776_ (_19482_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nand _51777_ (_19483_, _24779_, _24765_);
  and _51778_ (_19484_, _19483_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _51779_ (_19485_, _24793_, _24809_);
  and _51780_ (_19486_, _19485_, _19484_);
  or _51781_ (_19487_, _19486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor _51782_ (_19488_, _24803_, _24750_);
  nand _51783_ (_19489_, _19488_, _24807_);
  nor _51784_ (_19490_, _24765_, _24747_);
  or _51785_ (_19491_, _19490_, _24748_);
  and _51786_ (_19492_, _19491_, _19489_);
  and _51787_ (_19493_, _19492_, _19487_);
  or _51788_ (_19494_, _19493_, _19482_);
  and _51789_ (_11328_, _19494_, _22731_);
  and _51790_ (_19495_, _04950_, _24051_);
  and _51791_ (_19496_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or _51792_ (_11331_, _19496_, _19495_);
  and _51793_ (_11332_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _22731_);
  and _51794_ (_19497_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _51795_ (_19498_, _19490_, _24827_);
  and _51796_ (_19499_, _24804_, _24750_);
  nand _51797_ (_19500_, _19499_, _24781_);
  and _51798_ (_19501_, _19500_, _19498_);
  or _51799_ (_19502_, _19501_, _19497_);
  and _51800_ (_19503_, _19485_, _19483_);
  or _51801_ (_19504_, _19503_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _51802_ (_19505_, _19409_, rst);
  and _51803_ (_19506_, _19505_, _19504_);
  and _51804_ (_11334_, _19506_, _19502_);
  and _51805_ (_11336_, _26377_, _22731_);
  nor _51806_ (_19507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _17565_);
  not _51807_ (_19508_, _19413_);
  and _51808_ (_19509_, _19415_, _19508_);
  not _51809_ (_19510_, _19509_);
  or _51810_ (_19511_, _19510_, _19453_);
  and _51811_ (_19512_, _19511_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _51812_ (_19513_, _19512_, _19507_);
  and _51813_ (_19514_, _19458_, _24607_);
  or _51814_ (_19515_, _19514_, _19513_);
  nand _51815_ (_19516_, _19514_, _23504_);
  and _51816_ (_19517_, _19516_, _19515_);
  or _51817_ (_19518_, _19517_, _24703_);
  nand _51818_ (_19519_, _24703_, _24043_);
  and _51819_ (_19520_, _19519_, _22731_);
  and _51820_ (_11347_, _19520_, _19518_);
  and _51821_ (_19521_, _19458_, _24533_);
  and _51822_ (_19522_, _19521_, _24531_);
  nand _51823_ (_19523_, _24627_, _24188_);
  nand _51824_ (_19524_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _51825_ (_19525_, _19509_, _19408_);
  or _51826_ (_19526_, _19525_, _19524_);
  or _51827_ (_19527_, _19526_, _19521_);
  nand _51828_ (_19528_, _19527_, _19523_);
  or _51829_ (_19529_, _19528_, _19522_);
  or _51830_ (_19530_, _24704_, _23577_);
  and _51831_ (_19531_, _19530_, _22731_);
  and _51832_ (_11352_, _19531_, _19529_);
  and _51833_ (_19532_, _25481_, _24544_);
  nand _51834_ (_19533_, _19532_, _23504_);
  or _51835_ (_19534_, _19532_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _51836_ (_19535_, _19534_, _24557_);
  and _51837_ (_19536_, _19535_, _19533_);
  nor _51838_ (_19537_, _24557_, _23989_);
  or _51839_ (_19538_, _19537_, _19536_);
  and _51840_ (_11355_, _19538_, _22731_);
  and _51841_ (_19539_, _16020_, _23996_);
  and _51842_ (_19540_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or _51843_ (_11357_, _19540_, _19539_);
  and _51844_ (_26840_[5], _23765_, _22731_);
  nand _51845_ (_19541_, _24840_, _24749_);
  nand _51846_ (_19542_, _19396_, _24747_);
  and _51847_ (_19543_, _19542_, _22731_);
  and _51848_ (_11366_, _19543_, _19541_);
  and _51849_ (_19544_, _16678_, _24134_);
  and _51850_ (_19545_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _51851_ (_11369_, _19545_, _19544_);
  and _51852_ (_19546_, _24621_, _25481_);
  nand _51853_ (_19547_, _19546_, _23504_);
  or _51854_ (_19548_, _19546_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _51855_ (_19549_, _19548_, _24630_);
  and _51856_ (_19550_, _19549_, _19547_);
  nor _51857_ (_19551_, _24630_, _23989_);
  or _51858_ (_19552_, _19551_, _19550_);
  and _51859_ (_11372_, _19552_, _22731_);
  and _51860_ (_19553_, _25432_, _24051_);
  and _51861_ (_19554_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _51862_ (_11375_, _19554_, _19553_);
  and _51863_ (_19555_, _01832_, _23887_);
  and _51864_ (_19556_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _51865_ (_11380_, _19556_, _19555_);
  and _51866_ (_19557_, _25672_, _23887_);
  and _51867_ (_19558_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _51868_ (_11383_, _19558_, _19557_);
  and _51869_ (_19559_, _03324_, _24089_);
  and _51870_ (_19560_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _51871_ (_27260_, _19560_, _19559_);
  and _51872_ (_19561_, _04709_, _23887_);
  and _51873_ (_19562_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _51874_ (_11390_, _19562_, _19561_);
  and _51875_ (_19563_, _16072_, _23548_);
  and _51876_ (_19564_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or _51877_ (_26954_, _19564_, _19563_);
  or _51878_ (_19565_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand _51879_ (_19566_, _22740_, _04912_);
  and _51880_ (_19567_, _19566_, _22731_);
  and _51881_ (_26863_[15], _19567_, _19565_);
  nor _51882_ (_11407_, _00780_, rst);
  and _51883_ (_11408_, _00352_, _22731_);
  and _51884_ (_11411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _22731_);
  and _51885_ (_19568_, _17545_, _23996_);
  and _51886_ (_19569_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or _51887_ (_11425_, _19569_, _19568_);
  and _51888_ (_19570_, _04950_, _23996_);
  and _51889_ (_19571_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or _51890_ (_11436_, _19571_, _19570_);
  and _51891_ (_19572_, _02498_, _23887_);
  and _51892_ (_19573_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or _51893_ (_11439_, _19573_, _19572_);
  and _51894_ (_19574_, _03020_, _24089_);
  and _51895_ (_19575_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _51896_ (_11440_, _19575_, _19574_);
  and _51897_ (_19576_, _02767_, _24134_);
  and _51898_ (_19577_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _51899_ (_11442_, _19577_, _19576_);
  and _51900_ (_19578_, _03217_, _23548_);
  and _51901_ (_19579_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _51902_ (_27311_, _19579_, _19578_);
  and _51903_ (_19580_, _04647_, _24089_);
  and _51904_ (_19581_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _51905_ (_11446_, _19581_, _19580_);
  and _51906_ (_19582_, _01832_, _23583_);
  and _51907_ (_19583_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _51908_ (_11450_, _19583_, _19582_);
  and _51909_ (_19584_, _17545_, _24134_);
  and _51910_ (_19585_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _51911_ (_11452_, _19585_, _19584_);
  and _51912_ (_19586_, _03020_, _24051_);
  and _51913_ (_19587_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _51914_ (_11455_, _19587_, _19586_);
  or _51915_ (_19588_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _51916_ (_11462_, _19588_, _03411_);
  and _51917_ (_19589_, _03404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _51918_ (_11463_, _19589_, _03406_);
  or _51919_ (_19590_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _51920_ (_11466_, _19590_, _03423_);
  and _51921_ (_11475_, _00540_, _22731_);
  and _51922_ (_11486_, _16453_, _24747_);
  and _51923_ (_11487_, _00437_, _22731_);
  and _51924_ (_19591_, _15581_, _24134_);
  and _51925_ (_19592_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or _51926_ (_27210_, _19592_, _19591_);
  and _51927_ (_19593_, _02045_, _23996_);
  and _51928_ (_19594_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _51929_ (_27233_, _19594_, _19593_);
  and _51930_ (_19595_, _24051_, _23946_);
  and _51931_ (_19596_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or _51932_ (_11496_, _19596_, _19595_);
  and _51933_ (_11510_, _00708_, _22731_);
  and _51934_ (_19597_, _16020_, _23583_);
  and _51935_ (_19598_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  or _51936_ (_11512_, _19598_, _19597_);
  and _51937_ (_11514_, _26381_, _22731_);
  and _51938_ (_11517_, _00621_, _22731_);
  and _51939_ (_19599_, _05491_, _23583_);
  and _51940_ (_19600_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or _51941_ (_11519_, _19600_, _19599_);
  and _51942_ (_19601_, _15581_, _23996_);
  and _51943_ (_19602_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or _51944_ (_11526_, _19602_, _19601_);
  and _51945_ (_19603_, _24442_, _23996_);
  and _51946_ (_19604_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or _51947_ (_11528_, _19604_, _19603_);
  and _51948_ (_19606_, _04950_, _24219_);
  and _51949_ (_19607_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  or _51950_ (_11539_, _19607_, _19606_);
  and _51951_ (_19608_, _01810_, _23887_);
  and _51952_ (_19609_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or _51953_ (_11550_, _19609_, _19608_);
  and _51954_ (_19610_, _04768_, _24051_);
  and _51955_ (_19611_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _51956_ (_11553_, _19611_, _19610_);
  and _51957_ (_19612_, _01810_, _24089_);
  and _51958_ (_19613_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or _51959_ (_27217_, _19613_, _19612_);
  and _51960_ (_19614_, _17545_, _24051_);
  and _51961_ (_19615_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _51962_ (_27255_, _19615_, _19614_);
  and _51963_ (_19616_, _04709_, _23548_);
  and _51964_ (_19617_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _51965_ (_11563_, _19617_, _19616_);
  and _51966_ (_19618_, _04709_, _24051_);
  and _51967_ (_19619_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _51968_ (_11592_, _19619_, _19618_);
  and _51969_ (_19620_, _01810_, _23583_);
  and _51970_ (_19621_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or _51971_ (_11594_, _19621_, _19620_);
  and _51972_ (_19622_, _24889_, _23996_);
  and _51973_ (_19623_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _51974_ (_11596_, _19623_, _19622_);
  and _51975_ (_19624_, _17545_, _24089_);
  and _51976_ (_19625_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or _51977_ (_11601_, _19625_, _19624_);
  and _51978_ (_19626_, _03667_, _23548_);
  and _51979_ (_19627_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _51980_ (_11603_, _19627_, _19626_);
  and _51981_ (_19628_, _04950_, _23548_);
  and _51982_ (_19629_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  or _51983_ (_11605_, _19629_, _19628_);
  and _51984_ (_19630_, _03667_, _24051_);
  and _51985_ (_19631_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or _51986_ (_11611_, _19631_, _19630_);
  and _51987_ (_19632_, _24889_, _24134_);
  and _51988_ (_19633_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _51989_ (_11614_, _19633_, _19632_);
  and _51990_ (_19634_, _03313_, _23548_);
  and _51991_ (_19635_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or _51992_ (_27176_, _19635_, _19634_);
  and _51993_ (_19636_, _16034_, _24219_);
  and _51994_ (_19637_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or _51995_ (_11627_, _19637_, _19636_);
  and _51996_ (_19638_, _03324_, _23583_);
  and _51997_ (_19640_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _51998_ (_27259_, _19640_, _19638_);
  and _51999_ (_19641_, _03324_, _23548_);
  and _52000_ (_19642_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _52001_ (_11630_, _19642_, _19641_);
  and _52002_ (_19643_, _03251_, _24219_);
  and _52003_ (_19644_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _52004_ (_11632_, _19644_, _19643_);
  and _52005_ (_19645_, _03217_, _23996_);
  and _52006_ (_19646_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _52007_ (_11638_, _19646_, _19645_);
  and _52008_ (_19647_, _16020_, _24051_);
  and _52009_ (_19648_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or _52010_ (_11641_, _19648_, _19647_);
  and _52011_ (_19649_, _15996_, _23583_);
  and _52012_ (_19650_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or _52013_ (_11654_, _19650_, _19649_);
  and _52014_ (_19651_, _03217_, _23583_);
  and _52015_ (_19652_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _52016_ (_11656_, _19652_, _19651_);
  and _52017_ (_19653_, _01810_, _24051_);
  and _52018_ (_19654_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or _52019_ (_11658_, _19654_, _19653_);
  and _52020_ (_19655_, _03180_, _23887_);
  and _52021_ (_19656_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _52022_ (_26917_, _19656_, _19655_);
  and _52023_ (_19657_, _03048_, _24089_);
  and _52024_ (_19658_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or _52025_ (_11661_, _19658_, _19657_);
  and _52026_ (_19659_, _03048_, _23548_);
  and _52027_ (_19660_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _52028_ (_26932_, _19660_, _19659_);
  and _52029_ (_19661_, _04950_, _23583_);
  and _52030_ (_19662_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or _52031_ (_11685_, _19662_, _19661_);
  and _52032_ (_19663_, _02980_, _24089_);
  and _52033_ (_19664_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _52034_ (_11688_, _19664_, _19663_);
  and _52035_ (_19665_, _02498_, _24051_);
  and _52036_ (_19666_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _52037_ (_11691_, _19666_, _19665_);
  and _52038_ (_19667_, _16678_, _23548_);
  and _52039_ (_19668_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or _52040_ (_11694_, _19668_, _19667_);
  and _52041_ (_19669_, _02093_, _23887_);
  and _52042_ (_19670_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _52043_ (_11696_, _19670_, _19669_);
  and _52044_ (_19671_, _01832_, _23548_);
  and _52045_ (_19672_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _52046_ (_11699_, _19672_, _19671_);
  nor _52047_ (_19673_, _23531_, _26401_);
  and _52048_ (_19674_, _23531_, _26401_);
  or _52049_ (_19675_, _19674_, _19673_);
  and _52050_ (_11708_, _19675_, _22731_);
  and _52051_ (_19676_, _04950_, _23887_);
  and _52052_ (_19677_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  or _52053_ (_11711_, _19677_, _19676_);
  and _52054_ (_19678_, _02093_, _24134_);
  and _52055_ (_19679_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _52056_ (_27038_, _19679_, _19678_);
  and _52057_ (_19680_, _26020_, _24219_);
  and _52058_ (_19681_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or _52059_ (_11714_, _19681_, _19680_);
  and _52060_ (_11716_, _01167_, _22731_);
  and _52061_ (_11721_, _26457_, _22731_);
  and _52062_ (_11723_, _00449_, _22731_);
  and _52063_ (_11726_, _01042_, _22731_);
  and _52064_ (_11728_, _01253_, _22731_);
  and _52065_ (_11730_, _00364_, _22731_);
  and _52066_ (_11734_, _01325_, _22731_);
  and _52067_ (_11736_, _26560_, _22731_);
  and _52068_ (_11738_, _01099_, _22731_);
  and _52069_ (_11740_, _03830_, _22731_);
  and _52070_ (_11742_, _00627_, _22731_);
  and _52071_ (_11746_, _00530_, _22731_);
  and _52072_ (_19682_, _26020_, _23996_);
  and _52073_ (_19683_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or _52074_ (_11750_, _19683_, _19682_);
  and _52075_ (_19684_, _16678_, _24219_);
  and _52076_ (_19685_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _52077_ (_11752_, _19685_, _19684_);
  and _52078_ (_19686_, _25627_, _24134_);
  and _52079_ (_19687_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or _52080_ (_11754_, _19687_, _19686_);
  and _52081_ (_19688_, _25432_, _24089_);
  and _52082_ (_19689_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _52083_ (_11757_, _19689_, _19688_);
  and _52084_ (_19690_, _25432_, _23548_);
  and _52085_ (_19691_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _52086_ (_11759_, _19691_, _19690_);
  and _52087_ (_19692_, _25314_, _23583_);
  and _52088_ (_19693_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _52089_ (_11761_, _19693_, _19692_);
  and _52090_ (_19694_, _25210_, _24219_);
  and _52091_ (_19695_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or _52092_ (_27154_, _19695_, _19694_);
  and _52093_ (_11776_, _00715_, _22731_);
  and _52094_ (_19696_, _25210_, _24089_);
  and _52095_ (_19697_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or _52096_ (_11778_, _19697_, _19696_);
  and _52097_ (_19698_, _24478_, _24089_);
  and _52098_ (_19699_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _52099_ (_11792_, _19699_, _19698_);
  and _52100_ (_19700_, _16020_, _24219_);
  and _52101_ (_19701_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  or _52102_ (_11795_, _19701_, _19700_);
  and _52103_ (_19702_, _01810_, _24134_);
  and _52104_ (_19703_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or _52105_ (_11902_, _19703_, _19702_);
  and _52106_ (_19704_, _03287_, _23583_);
  and _52107_ (_19705_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  or _52108_ (_11906_, _19705_, _19704_);
  and _52109_ (_19706_, _16020_, _23548_);
  and _52110_ (_19707_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or _52111_ (_11909_, _19707_, _19706_);
  and _52112_ (_19708_, _03309_, _23583_);
  and _52113_ (_19709_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  or _52114_ (_11914_, _19709_, _19708_);
  and _52115_ (_19710_, _11419_, _24219_);
  and _52116_ (_19711_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or _52117_ (_11916_, _19711_, _19710_);
  and _52118_ (_19712_, _07779_, _24134_);
  and _52119_ (_19713_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  or _52120_ (_11920_, _19713_, _19712_);
  and _52121_ (_19714_, _02065_, _23996_);
  and _52122_ (_19715_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or _52123_ (_11925_, _19715_, _19714_);
  and _52124_ (_19716_, _08578_, _24219_);
  and _52125_ (_19717_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or _52126_ (_11927_, _19717_, _19716_);
  and _52127_ (_19718_, _15605_, _23548_);
  and _52128_ (_19719_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or _52129_ (_27179_, _19719_, _19718_);
  and _52130_ (_19720_, _16026_, _24089_);
  and _52131_ (_19721_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or _52132_ (_26949_, _19721_, _19720_);
  and _52133_ (_19722_, _16026_, _23583_);
  and _52134_ (_19723_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or _52135_ (_11932_, _19723_, _19722_);
  and _52136_ (_11934_, _01000_, _22731_);
  and _52137_ (_19724_, _03287_, _24051_);
  and _52138_ (_19725_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or _52139_ (_11937_, _19725_, _19724_);
  and _52140_ (_19726_, _03287_, _24089_);
  and _52141_ (_19727_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  or _52142_ (_12092_, _19727_, _19726_);
  and _52143_ (_26840_[0], _23681_, _22731_);
  and _52144_ (_19728_, _16704_, _23548_);
  and _52145_ (_19729_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or _52146_ (_12140_, _19729_, _19728_);
  and _52147_ (_19730_, _16704_, _23583_);
  and _52148_ (_19731_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or _52149_ (_12142_, _19731_, _19730_);
  and _52150_ (_19732_, _03043_, _24089_);
  and _52151_ (_19733_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or _52152_ (_12148_, _19733_, _19732_);
  and _52153_ (_19734_, _16704_, _23887_);
  and _52154_ (_19735_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or _52155_ (_12154_, _19735_, _19734_);
  nor _52156_ (_19736_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _52157_ (_19737_, _19736_);
  and _52158_ (_19738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _52159_ (_19739_, _19738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _52160_ (_19740_, _19738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _52161_ (_19741_, _19740_, _19739_);
  not _52162_ (_19742_, _19741_);
  and _52163_ (_19743_, _19739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52164_ (_19744_, _19739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52165_ (_19745_, _19744_, _19743_);
  nor _52166_ (_19746_, _19745_, _05614_);
  and _52167_ (_19747_, _19745_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _52168_ (_19748_, _19747_, _19746_);
  nor _52169_ (_19749_, _19748_, _19742_);
  nor _52170_ (_19750_, _19745_, _05653_);
  and _52171_ (_19751_, _19745_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _52172_ (_19752_, _19751_, _19750_);
  nor _52173_ (_19753_, _19752_, _19741_);
  nor _52174_ (_19754_, _19753_, _19749_);
  nor _52175_ (_19755_, _19754_, _19737_);
  and _52176_ (_19756_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _22742_);
  not _52177_ (_19757_, _19756_);
  and _52178_ (_19758_, _19745_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _52179_ (_19759_, _19745_, _05641_);
  nor _52180_ (_19760_, _19759_, _19758_);
  nor _52181_ (_19761_, _19760_, _19742_);
  nor _52182_ (_19762_, _19745_, _05634_);
  and _52183_ (_19763_, _19745_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _52184_ (_19764_, _19763_, _19762_);
  nor _52185_ (_19765_, _19764_, _19741_);
  nor _52186_ (_19766_, _19765_, _19761_);
  nor _52187_ (_19767_, _19766_, _19757_);
  nor _52188_ (_19768_, _19767_, _19755_);
  not _52189_ (_19769_, _19738_);
  nor _52190_ (_19770_, _19745_, _05660_);
  and _52191_ (_19771_, _19745_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _52192_ (_19772_, _19771_, _19770_);
  nor _52193_ (_19773_, _19772_, _19742_);
  not _52194_ (_19774_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _52195_ (_19775_, _19745_, _19774_);
  and _52196_ (_19776_, _19745_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _52197_ (_19777_, _19776_, _19775_);
  nor _52198_ (_19778_, _19777_, _19741_);
  nor _52199_ (_19779_, _19778_, _19773_);
  nor _52200_ (_19780_, _19779_, _19769_);
  and _52201_ (_19781_, _22747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _52202_ (_19782_, _19781_);
  and _52203_ (_19783_, _19745_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _52204_ (_19784_, _19745_, _06106_);
  nor _52205_ (_19785_, _19784_, _19783_);
  nor _52206_ (_19786_, _19785_, _19742_);
  not _52207_ (_19787_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _52208_ (_19788_, _19745_, _19787_);
  and _52209_ (_19789_, _19745_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _52210_ (_19790_, _19789_, _19788_);
  nor _52211_ (_19791_, _19790_, _19741_);
  nor _52212_ (_19792_, _19791_, _19786_);
  nor _52213_ (_19793_, _19792_, _19782_);
  nor _52214_ (_19794_, _19793_, _19780_);
  and _52215_ (_19795_, _19794_, _19768_);
  and _52216_ (_19796_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _52217_ (_19797_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor _52218_ (_19798_, _19797_, _19796_);
  and _52219_ (_19799_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _52220_ (_19800_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _52221_ (_19801_, _19800_, _19799_);
  and _52222_ (_19802_, _19801_, _19798_);
  and _52223_ (_19803_, _19802_, _19742_);
  and _52224_ (_19804_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _52225_ (_19805_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _52226_ (_19806_, _19805_, _19804_);
  and _52227_ (_19807_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _52228_ (_19808_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _52229_ (_19809_, _19808_, _19807_);
  and _52230_ (_19810_, _19809_, _19806_);
  and _52231_ (_19811_, _19810_, _19741_);
  or _52232_ (_19812_, _19811_, _19745_);
  nor _52233_ (_19813_, _19812_, _19803_);
  and _52234_ (_19814_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _52235_ (_19815_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor _52236_ (_19816_, _19815_, _19814_);
  and _52237_ (_19817_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _52238_ (_19818_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _52239_ (_19819_, _19818_, _19817_);
  and _52240_ (_19820_, _19819_, _19816_);
  nor _52241_ (_19821_, _19820_, _19741_);
  and _52242_ (_19822_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _52243_ (_19823_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _52244_ (_19824_, _19823_, _19822_);
  and _52245_ (_19825_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _52246_ (_19826_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _52247_ (_19827_, _19826_, _19825_);
  and _52248_ (_19828_, _19827_, _19824_);
  nor _52249_ (_19829_, _19828_, _19742_);
  or _52250_ (_19830_, _19829_, _19821_);
  and _52251_ (_19831_, _19830_, _19745_);
  nor _52252_ (_19832_, _19831_, _19813_);
  nor _52253_ (_19833_, _19832_, _19795_);
  and _52254_ (_19834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _52255_ (_19835_, _19834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _52256_ (_19836_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _52257_ (_19837_, _19836_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _52258_ (_19838_, _19837_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _52259_ (_19839_, _19838_, _19835_);
  and _52260_ (_19840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _52261_ (_19841_, _19840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _52262_ (_19842_, _19841_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _52263_ (_19843_, _19842_, _19839_);
  and _52264_ (_19844_, _19843_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _52265_ (_19845_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _52266_ (_19846_, _19845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and _52267_ (_19847_, _19845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _52268_ (_19848_, _19847_, _19846_);
  and _52269_ (_19849_, _19848_, _19833_);
  nor _52270_ (_19850_, _19844_, _22802_);
  and _52271_ (_19851_, _19841_, _19839_);
  and _52272_ (_19852_, _19851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _52273_ (_19853_, _19852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _52274_ (_19854_, _19853_, _22802_);
  nor _52275_ (_19855_, _19854_, _19850_);
  not _52276_ (_19856_, _19855_);
  and _52277_ (_19857_, _19856_, _19833_);
  nor _52278_ (_19858_, _19843_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _52279_ (_19859_, _19858_, _19844_);
  and _52280_ (_19860_, _19859_, _19833_);
  nor _52281_ (_19861_, _19856_, _19833_);
  nor _52282_ (_19862_, _19861_, _19857_);
  nor _52283_ (_19863_, _19851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _52284_ (_19864_, _19863_, _19852_);
  and _52285_ (_19865_, _19864_, _19833_);
  and _52286_ (_19866_, _19840_, _19839_);
  nor _52287_ (_19867_, _19866_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _52288_ (_19868_, _19867_, _19851_);
  and _52289_ (_19869_, _19868_, _19833_);
  nor _52290_ (_19870_, _19864_, _19833_);
  nor _52291_ (_19871_, _19870_, _19865_);
  nor _52292_ (_19872_, _19868_, _19833_);
  nor _52293_ (_19873_, _19872_, _19869_);
  not _52294_ (_19874_, _19873_);
  and _52295_ (_19875_, _19839_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _52296_ (_19876_, _19875_, _22784_);
  nor _52297_ (_19877_, _19875_, _22784_);
  nor _52298_ (_19878_, _19877_, _19876_);
  not _52299_ (_19879_, _19878_);
  and _52300_ (_19880_, _19879_, _19833_);
  nor _52301_ (_19881_, _19839_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _52302_ (_19882_, _19881_, _19875_);
  and _52303_ (_19883_, _19882_, _19833_);
  nor _52304_ (_19884_, _19879_, _19833_);
  nor _52305_ (_19885_, _19884_, _19880_);
  and _52306_ (_19886_, _19837_, _19835_);
  nor _52307_ (_19887_, _19886_, _22776_);
  and _52308_ (_19888_, _19886_, _22776_);
  nor _52309_ (_19889_, _19888_, _19887_);
  not _52310_ (_19890_, _19889_);
  and _52311_ (_19891_, _19890_, _19833_);
  nor _52312_ (_19892_, _19890_, _19833_);
  nor _52313_ (_19893_, _19892_, _19891_);
  not _52314_ (_19894_, _19893_);
  not _52315_ (_19895_, _19795_);
  not _52316_ (_19896_, _19745_);
  and _52317_ (_19897_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _52318_ (_19898_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _52319_ (_19899_, _19898_, _19897_);
  and _52320_ (_19900_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _52321_ (_19901_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _52322_ (_19902_, _19901_, _19900_);
  and _52323_ (_19903_, _19902_, _19899_);
  and _52324_ (_19904_, _19903_, _19742_);
  and _52325_ (_19905_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _52326_ (_19906_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _52327_ (_19908_, _19906_, _19905_);
  and _52328_ (_19909_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _52329_ (_19910_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _52330_ (_19911_, _19910_, _19909_);
  and _52331_ (_19912_, _19911_, _19908_);
  and _52332_ (_19913_, _19912_, _19741_);
  nor _52333_ (_19914_, _19913_, _19904_);
  nor _52334_ (_19915_, _19914_, _19896_);
  and _52335_ (_19916_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _52336_ (_19917_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _52337_ (_19918_, _19917_, _19916_);
  and _52338_ (_19919_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _52339_ (_19920_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _52340_ (_19921_, _19920_, _19919_);
  and _52341_ (_19922_, _19921_, _19918_);
  and _52342_ (_19923_, _19922_, _19742_);
  and _52343_ (_19924_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _52344_ (_19925_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _52345_ (_19926_, _19925_, _19924_);
  and _52346_ (_19927_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _52347_ (_19928_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _52348_ (_19929_, _19928_, _19927_);
  and _52349_ (_19930_, _19929_, _19926_);
  and _52350_ (_19931_, _19930_, _19741_);
  nor _52351_ (_19932_, _19931_, _19923_);
  nor _52352_ (_19933_, _19932_, _19745_);
  nor _52353_ (_19934_, _19933_, _19915_);
  and _52354_ (_19935_, _19934_, _19895_);
  and _52355_ (_19936_, _19836_, _19835_);
  nor _52356_ (_19937_, _19936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _52357_ (_19938_, _19937_, _19886_);
  and _52358_ (_19939_, _19938_, _19935_);
  nor _52359_ (_19940_, _19938_, _19935_);
  nor _52360_ (_19941_, _19940_, _19939_);
  and _52361_ (_19942_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _52362_ (_19943_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _52363_ (_19944_, _19943_, _19942_);
  and _52364_ (_19945_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _52365_ (_19946_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _52366_ (_19947_, _19946_, _19945_);
  and _52367_ (_19948_, _19947_, _19944_);
  and _52368_ (_19949_, _19948_, _19741_);
  and _52369_ (_19950_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _52370_ (_19951_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _52371_ (_19952_, _19951_, _19950_);
  and _52372_ (_19953_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _52373_ (_19954_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _52374_ (_19955_, _19954_, _19953_);
  and _52375_ (_19956_, _19955_, _19952_);
  and _52376_ (_19957_, _19956_, _19742_);
  nor _52377_ (_19958_, _19957_, _19949_);
  nor _52378_ (_19959_, _19958_, _19896_);
  and _52379_ (_19960_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _52380_ (_19961_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _52381_ (_19962_, _19961_, _19960_);
  and _52382_ (_19963_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _52383_ (_19964_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _52384_ (_19965_, _19964_, _19963_);
  and _52385_ (_19966_, _19965_, _19962_);
  and _52386_ (_19967_, _19966_, _19742_);
  and _52387_ (_19968_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _52388_ (_19969_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _52389_ (_19970_, _19969_, _19968_);
  and _52390_ (_19971_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _52391_ (_19972_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _52392_ (_19973_, _19972_, _19971_);
  and _52393_ (_19974_, _19973_, _19970_);
  and _52394_ (_19975_, _19974_, _19741_);
  nor _52395_ (_19976_, _19975_, _19967_);
  nor _52396_ (_19977_, _19976_, _19745_);
  nor _52397_ (_19978_, _19977_, _19959_);
  and _52398_ (_19979_, _19978_, _19895_);
  and _52399_ (_19980_, _19835_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _52400_ (_19981_, _19980_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _52401_ (_19982_, _19981_, _19936_);
  and _52402_ (_19983_, _19982_, _19979_);
  nor _52403_ (_19984_, _19982_, _19979_);
  and _52404_ (_19985_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _52405_ (_19986_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _52406_ (_19987_, _19986_, _19985_);
  and _52407_ (_19988_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _52408_ (_19989_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _52409_ (_19990_, _19989_, _19988_);
  and _52410_ (_19991_, _19990_, _19987_);
  and _52411_ (_19992_, _19991_, _19742_);
  and _52412_ (_19993_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _52413_ (_19994_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _52414_ (_19995_, _19994_, _19993_);
  and _52415_ (_19996_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _52416_ (_19997_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _52417_ (_19998_, _19997_, _19996_);
  and _52418_ (_19999_, _19998_, _19995_);
  and _52419_ (_20000_, _19999_, _19741_);
  or _52420_ (_20001_, _20000_, _19745_);
  nor _52421_ (_20002_, _20001_, _19992_);
  and _52422_ (_20003_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _52423_ (_20004_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _52424_ (_20005_, _20004_, _20003_);
  and _52425_ (_20006_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _52426_ (_20007_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _52427_ (_20008_, _20007_, _20006_);
  and _52428_ (_20009_, _20008_, _20005_);
  nor _52429_ (_20010_, _20009_, _19741_);
  and _52430_ (_20011_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _52431_ (_20012_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _52432_ (_20013_, _20012_, _20011_);
  and _52433_ (_20014_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _52434_ (_20015_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _52435_ (_20016_, _20015_, _20014_);
  and _52436_ (_20017_, _20016_, _20013_);
  nor _52437_ (_20018_, _20017_, _19742_);
  or _52438_ (_20019_, _20018_, _20010_);
  and _52439_ (_20020_, _20019_, _19745_);
  nor _52440_ (_20021_, _20020_, _20002_);
  nor _52441_ (_20022_, _20021_, _19795_);
  nor _52442_ (_20023_, _19835_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _52443_ (_20024_, _20023_, _19980_);
  and _52444_ (_20025_, _20024_, _20022_);
  and _52445_ (_20026_, _19834_, _22758_);
  nor _52446_ (_20027_, _19834_, _22758_);
  nor _52447_ (_20028_, _20027_, _20026_);
  not _52448_ (_20029_, _20028_);
  and _52449_ (_20030_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _52450_ (_20031_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _52451_ (_20032_, _20031_, _20030_);
  and _52452_ (_20033_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _52453_ (_20034_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _52454_ (_20035_, _20034_, _20033_);
  and _52455_ (_20036_, _20035_, _20032_);
  and _52456_ (_20037_, _20036_, _19742_);
  and _52457_ (_20038_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _52458_ (_20039_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _52459_ (_20040_, _20039_, _20038_);
  and _52460_ (_20041_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _52461_ (_20042_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _52462_ (_20043_, _20042_, _20041_);
  and _52463_ (_20044_, _20043_, _20040_);
  and _52464_ (_20045_, _20044_, _19741_);
  or _52465_ (_20046_, _20045_, _19745_);
  nor _52466_ (_20047_, _20046_, _20037_);
  and _52467_ (_20048_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _52468_ (_20049_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _52469_ (_20050_, _20049_, _20048_);
  and _52470_ (_20051_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _52471_ (_20052_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _52472_ (_20053_, _20052_, _20051_);
  and _52473_ (_20054_, _20053_, _20050_);
  nor _52474_ (_20055_, _20054_, _19741_);
  and _52475_ (_20056_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _52476_ (_20057_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _52477_ (_20058_, _20057_, _20056_);
  and _52478_ (_20059_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _52479_ (_20060_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _52480_ (_20061_, _20060_, _20059_);
  and _52481_ (_20062_, _20061_, _20058_);
  nor _52482_ (_20063_, _20062_, _19742_);
  or _52483_ (_20064_, _20063_, _20055_);
  and _52484_ (_20065_, _20064_, _19745_);
  nor _52485_ (_20066_, _20065_, _20047_);
  nor _52486_ (_20067_, _20066_, _19795_);
  and _52487_ (_20068_, _20067_, _20029_);
  nor _52488_ (_20069_, _20067_, _20029_);
  nor _52489_ (_20070_, _20069_, _20068_);
  not _52490_ (_20071_, _20070_);
  and _52491_ (_20072_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _52492_ (_20073_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _52493_ (_20074_, _20073_, _20072_);
  and _52494_ (_20075_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _52495_ (_20076_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _52496_ (_20077_, _20076_, _20075_);
  and _52497_ (_20078_, _20077_, _20074_);
  and _52498_ (_20079_, _20078_, _19742_);
  and _52499_ (_20080_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _52500_ (_20081_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _52501_ (_20082_, _20081_, _20080_);
  and _52502_ (_20083_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _52503_ (_20084_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _52504_ (_20085_, _20084_, _20083_);
  and _52505_ (_20086_, _20085_, _20082_);
  and _52506_ (_20087_, _20086_, _19741_);
  nor _52507_ (_20088_, _20087_, _20079_);
  nor _52508_ (_20089_, _20088_, _19896_);
  and _52509_ (_20090_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _52510_ (_20091_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _52511_ (_20092_, _20091_, _20090_);
  and _52512_ (_20093_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _52513_ (_20094_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _52514_ (_20095_, _20094_, _20093_);
  and _52515_ (_20096_, _20095_, _20092_);
  and _52516_ (_20097_, _20096_, _19742_);
  and _52517_ (_20098_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _52518_ (_20099_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _52519_ (_20100_, _20099_, _20098_);
  and _52520_ (_20101_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _52521_ (_20102_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _52522_ (_20103_, _20102_, _20101_);
  and _52523_ (_20104_, _20103_, _20100_);
  and _52524_ (_20105_, _20104_, _19741_);
  nor _52525_ (_20106_, _20105_, _20097_);
  nor _52526_ (_20107_, _20106_, _19745_);
  nor _52527_ (_20108_, _20107_, _20089_);
  and _52528_ (_20109_, _20108_, _19895_);
  and _52529_ (_20110_, _22752_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _52530_ (_20111_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _22747_);
  nor _52531_ (_20112_, _20111_, _20110_);
  not _52532_ (_20113_, _20112_);
  and _52533_ (_20114_, _20113_, _20109_);
  and _52534_ (_20115_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _52535_ (_20116_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _52536_ (_20117_, _20116_, _20115_);
  and _52537_ (_20118_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _52538_ (_20119_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _52539_ (_20120_, _20119_, _20118_);
  and _52540_ (_20121_, _20120_, _20117_);
  and _52541_ (_20122_, _20121_, _19742_);
  and _52542_ (_20123_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _52543_ (_20124_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _52544_ (_20125_, _20124_, _20123_);
  and _52545_ (_20126_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _52546_ (_20127_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _52547_ (_20128_, _20127_, _20126_);
  and _52548_ (_20129_, _20128_, _20125_);
  and _52549_ (_20130_, _20129_, _19741_);
  or _52550_ (_20131_, _20130_, _19745_);
  nor _52551_ (_20132_, _20131_, _20122_);
  and _52552_ (_20133_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _52553_ (_20134_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _52554_ (_20135_, _20134_, _20133_);
  and _52555_ (_20136_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _52556_ (_20137_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _52557_ (_20138_, _20137_, _20136_);
  and _52558_ (_20139_, _20138_, _20135_);
  nor _52559_ (_20140_, _20139_, _19741_);
  and _52560_ (_20141_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _52561_ (_20142_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _52562_ (_20143_, _20142_, _20141_);
  and _52563_ (_20144_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _52564_ (_20145_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _52565_ (_20146_, _20145_, _20144_);
  and _52566_ (_20147_, _20146_, _20143_);
  nor _52567_ (_20148_, _20147_, _19742_);
  or _52568_ (_20149_, _20148_, _20140_);
  and _52569_ (_20150_, _20149_, _19745_);
  nor _52570_ (_20151_, _20150_, _20132_);
  nor _52571_ (_20152_, _20151_, _19795_);
  and _52572_ (_20153_, _20152_, _22747_);
  and _52573_ (_20154_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _52574_ (_20155_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _52575_ (_20156_, _20155_, _20154_);
  and _52576_ (_20157_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _52577_ (_20158_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _52578_ (_20159_, _20158_, _20157_);
  and _52579_ (_20160_, _20159_, _20156_);
  and _52580_ (_20161_, _20160_, _19742_);
  and _52581_ (_20162_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _52582_ (_20163_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _52583_ (_20164_, _20163_, _20162_);
  and _52584_ (_20165_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _52585_ (_20166_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _52586_ (_20167_, _20166_, _20165_);
  and _52587_ (_20168_, _20167_, _20164_);
  and _52588_ (_20169_, _20168_, _19741_);
  or _52589_ (_20170_, _20169_, _19745_);
  nor _52590_ (_20171_, _20170_, _20161_);
  and _52591_ (_20172_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _52592_ (_20173_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor _52593_ (_20174_, _20173_, _20172_);
  and _52594_ (_20175_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _52595_ (_20176_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _52596_ (_20177_, _20176_, _20175_);
  and _52597_ (_20178_, _20177_, _20174_);
  nor _52598_ (_20179_, _20178_, _19741_);
  and _52599_ (_20180_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _52600_ (_20181_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _52601_ (_20182_, _20181_, _20180_);
  and _52602_ (_20183_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _52603_ (_20184_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _52604_ (_20185_, _20184_, _20183_);
  and _52605_ (_20186_, _20185_, _20182_);
  nor _52606_ (_20187_, _20186_, _19742_);
  or _52607_ (_20188_, _20187_, _20179_);
  and _52608_ (_20189_, _20188_, _19745_);
  nor _52609_ (_20190_, _20189_, _20171_);
  nor _52610_ (_20191_, _20190_, _19795_);
  and _52611_ (_20192_, _20191_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _52612_ (_20193_, _20152_, _22747_);
  nor _52613_ (_20194_, _20193_, _20153_);
  and _52614_ (_20195_, _20194_, _20192_);
  nor _52615_ (_20196_, _20195_, _20153_);
  nor _52616_ (_20197_, _20113_, _20109_);
  nor _52617_ (_20198_, _20197_, _20114_);
  not _52618_ (_20199_, _20198_);
  nor _52619_ (_20200_, _20199_, _20196_);
  nor _52620_ (_20201_, _20200_, _20114_);
  nor _52621_ (_20202_, _20201_, _20071_);
  nor _52622_ (_20203_, _20202_, _20068_);
  nor _52623_ (_20204_, _20024_, _20022_);
  nor _52624_ (_20205_, _20204_, _20025_);
  not _52625_ (_20206_, _20205_);
  nor _52626_ (_20207_, _20206_, _20203_);
  nor _52627_ (_20208_, _20207_, _20025_);
  nor _52628_ (_20209_, _20208_, _19984_);
  or _52629_ (_20210_, _20209_, _19983_);
  and _52630_ (_20211_, _20210_, _19941_);
  nor _52631_ (_20212_, _20211_, _19939_);
  nor _52632_ (_20213_, _20212_, _19894_);
  nor _52633_ (_20214_, _20213_, _19891_);
  nor _52634_ (_20215_, _19882_, _19833_);
  nor _52635_ (_20216_, _20215_, _19883_);
  not _52636_ (_20217_, _20216_);
  nor _52637_ (_20218_, _20217_, _20214_);
  and _52638_ (_20219_, _20218_, _19885_);
  or _52639_ (_20220_, _20219_, _19883_);
  nor _52640_ (_20221_, _20220_, _19880_);
  nor _52641_ (_20222_, _20221_, _19874_);
  and _52642_ (_20223_, _20222_, _19871_);
  or _52643_ (_20224_, _20223_, _19869_);
  nor _52644_ (_20225_, _20224_, _19865_);
  nor _52645_ (_20226_, _19859_, _19833_);
  nor _52646_ (_20227_, _20226_, _19860_);
  not _52647_ (_20228_, _20227_);
  nor _52648_ (_20229_, _20228_, _20225_);
  and _52649_ (_20230_, _20229_, _19862_);
  or _52650_ (_20231_, _20230_, _19860_);
  nor _52651_ (_20232_, _20231_, _19857_);
  nor _52652_ (_20233_, _19848_, _19833_);
  nor _52653_ (_20234_, _20233_, _19849_);
  not _52654_ (_20235_, _20234_);
  nor _52655_ (_20236_, _20235_, _20232_);
  nor _52656_ (_20237_, _20236_, _19849_);
  nor _52657_ (_20238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _52658_ (_20239_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _52659_ (_20240_, _20239_, _20238_);
  not _52660_ (_20241_, _20240_);
  nor _52661_ (_20242_, _20241_, _19847_);
  and _52662_ (_20243_, _20241_, _19847_);
  nor _52663_ (_20244_, _20243_, _20242_);
  not _52664_ (_20245_, _20244_);
  and _52665_ (_20246_, _20245_, _19833_);
  nor _52666_ (_20247_, _20245_, _19833_);
  nor _52667_ (_20248_, _20247_, _20246_);
  not _52668_ (_20249_, _20248_);
  nand _52669_ (_20250_, _20249_, _20237_);
  or _52670_ (_20251_, _20249_, _20237_);
  and _52671_ (_20252_, _20251_, _20250_);
  and _52672_ (_20253_, _20235_, _20232_);
  nor _52673_ (_20254_, _20253_, _20236_);
  nand _52674_ (_20255_, _20254_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or _52675_ (_20256_, _20254_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _52676_ (_20257_, _20256_, _20255_);
  nor _52677_ (_20258_, _20229_, _19860_);
  nor _52678_ (_20259_, _19855_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _52679_ (_20260_, _19855_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or _52680_ (_20261_, _20260_, _20259_);
  nand _52681_ (_20262_, _20261_, _19833_);
  or _52682_ (_20263_, _20261_, _19833_);
  and _52683_ (_20264_, _20263_, _20262_);
  not _52684_ (_20265_, _20264_);
  nand _52685_ (_20266_, _20265_, _20258_);
  or _52686_ (_20267_, _20265_, _20258_);
  and _52687_ (_20268_, _20267_, _20266_);
  and _52688_ (_20269_, _20228_, _20225_);
  nor _52689_ (_20270_, _20269_, _20229_);
  nor _52690_ (_20271_, _20270_, _22797_);
  and _52691_ (_20272_, _20270_, _22797_);
  nor _52692_ (_20273_, _20218_, _19883_);
  and _52693_ (_20274_, _20273_, _19885_);
  nor _52694_ (_20275_, _20273_, _19885_);
  nor _52695_ (_20276_, _20275_, _20274_);
  and _52696_ (_20277_, _20276_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _52697_ (_20278_, _20276_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _52698_ (_20279_, _20217_, _20214_);
  nor _52699_ (_20280_, _20279_, _20218_);
  nor _52700_ (_20281_, _20280_, _22780_);
  and _52701_ (_20282_, _20280_, _22780_);
  and _52702_ (_20283_, _20212_, _19894_);
  nor _52703_ (_20284_, _20283_, _20213_);
  and _52704_ (_20285_, _20284_, _26136_);
  nor _52705_ (_20286_, _20284_, _26136_);
  nor _52706_ (_20287_, _19983_, _19984_);
  nor _52707_ (_20288_, _20287_, _20208_);
  and _52708_ (_20289_, _20287_, _20208_);
  or _52709_ (_20290_, _20289_, _20288_);
  and _52710_ (_20291_, _20290_, _22767_);
  nor _52711_ (_20292_, _20290_, _22767_);
  and _52712_ (_20293_, _20206_, _20203_);
  nor _52713_ (_20294_, _20293_, _20207_);
  and _52714_ (_20295_, _20294_, _22762_);
  nor _52715_ (_20296_, _20294_, _22762_);
  and _52716_ (_20297_, _20201_, _20071_);
  nor _52717_ (_20298_, _20297_, _20202_);
  and _52718_ (_20299_, _20298_, _26149_);
  nor _52719_ (_20300_, _20298_, _26149_);
  and _52720_ (_20301_, _20199_, _20196_);
  nor _52721_ (_20302_, _20301_, _20200_);
  and _52722_ (_20303_, _20302_, _26153_);
  nor _52723_ (_20304_, _20302_, _26153_);
  and _52724_ (_20305_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _52725_ (_20306_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _52726_ (_20307_, _20306_, _20305_);
  not _52727_ (_20308_, _20307_);
  nand _52728_ (_20309_, _20308_, _20191_);
  or _52729_ (_20310_, _20308_, _20191_);
  and _52730_ (_20311_, _20310_, _20309_);
  nor _52731_ (_20312_, _20194_, _20192_);
  nor _52732_ (_20313_, _20312_, _20195_);
  and _52733_ (_20314_, _20313_, _09640_);
  or _52734_ (_20315_, _20314_, _20311_);
  nor _52735_ (_20316_, _20313_, _09640_);
  or _52736_ (_20317_, _20316_, _20315_);
  or _52737_ (_20318_, _20317_, _20304_);
  or _52738_ (_20319_, _20318_, _20303_);
  or _52739_ (_20320_, _20319_, _20300_);
  or _52740_ (_20321_, _20320_, _20299_);
  or _52741_ (_20322_, _20321_, _20296_);
  or _52742_ (_20323_, _20322_, _20295_);
  or _52743_ (_20324_, _20323_, _20292_);
  or _52744_ (_20325_, _20324_, _20291_);
  nor _52745_ (_20326_, _20210_, _19941_);
  nor _52746_ (_20327_, _20326_, _20211_);
  nor _52747_ (_20328_, _20327_, _22772_);
  and _52748_ (_20329_, _20327_, _22772_);
  or _52749_ (_20330_, _20329_, _20328_);
  or _52750_ (_20331_, _20330_, _20325_);
  or _52751_ (_20332_, _20331_, _20286_);
  or _52752_ (_20333_, _20332_, _20285_);
  or _52753_ (_20334_, _20333_, _20282_);
  or _52754_ (_20335_, _20334_, _20281_);
  or _52755_ (_20336_, _20335_, _20278_);
  or _52756_ (_20337_, _20336_, _20277_);
  and _52757_ (_20338_, _20221_, _19874_);
  nor _52758_ (_20339_, _20338_, _20222_);
  and _52759_ (_20340_, _20339_, _22789_);
  nor _52760_ (_20341_, _20339_, _22789_);
  or _52761_ (_20342_, _20341_, _20340_);
  nor _52762_ (_20343_, _20222_, _19869_);
  and _52763_ (_20344_, _19871_, _22793_);
  nor _52764_ (_20345_, _19871_, _22793_);
  nor _52765_ (_20346_, _20345_, _20344_);
  nand _52766_ (_20347_, _20346_, _20343_);
  or _52767_ (_20348_, _20346_, _20343_);
  and _52768_ (_20349_, _20348_, _20347_);
  or _52769_ (_20350_, _20349_, _20342_);
  or _52770_ (_20351_, _20350_, _20337_);
  or _52771_ (_20352_, _20351_, _20272_);
  or _52772_ (_20353_, _20352_, _20271_);
  or _52773_ (_20354_, _20353_, _20268_);
  or _52774_ (_20355_, _20354_, _20257_);
  or _52775_ (_20356_, _20355_, _20252_);
  and _52776_ (_20357_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _52777_ (_20358_, _20357_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _52778_ (_20359_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _52779_ (_20360_, _20359_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _52780_ (_20361_, _20360_, _20358_);
  not _52781_ (_20362_, _20361_);
  not _52782_ (_20363_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _52783_ (_20364_, _20358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _52784_ (_20365_, _20358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _52785_ (_20366_, _20365_, _20364_);
  nand _52786_ (_20367_, _20366_, _20363_);
  or _52787_ (_20368_, _20366_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _52788_ (_20369_, _20368_, _20367_);
  and _52789_ (_20370_, _20369_, _20362_);
  not _52790_ (_20371_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand _52791_ (_20372_, _20366_, _20371_);
  or _52792_ (_20373_, _20366_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _52793_ (_20374_, _20373_, _20361_);
  and _52794_ (_20375_, _20374_, _20372_);
  or _52795_ (_20376_, _20375_, _20370_);
  or _52796_ (_20377_, _20376_, _09640_);
  and _52797_ (_20378_, _26153_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _52798_ (_20379_, \oc8051_symbolic_cxrom1.regvalid [5], _26149_);
  and _52799_ (_20380_, \oc8051_symbolic_cxrom1.regvalid [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _52800_ (_20381_, _20380_, _20379_);
  and _52801_ (_20382_, _20381_, _20378_);
  or _52802_ (_20383_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _52803_ (_20384_, \oc8051_symbolic_cxrom1.regvalid [1], _26149_);
  and _52804_ (_20385_, _20384_, _20357_);
  and _52805_ (_20386_, _20385_, _20383_);
  or _52806_ (_20387_, _20386_, _20382_);
  nor _52807_ (_20388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _52808_ (_20389_, _20388_, _26153_);
  nor _52809_ (_20390_, _20389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _52810_ (_20391_, _20389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _52811_ (_20392_, _20391_, _20390_);
  and _52812_ (_20393_, _20392_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _52813_ (_20394_, _20388_, _26153_);
  nor _52814_ (_20395_, _20394_, _20389_);
  or _52815_ (_20396_, _05641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _52816_ (_20397_, _20396_, _20395_);
  or _52817_ (_20398_, _20397_, _20393_);
  and _52818_ (_20399_, _20398_, _09640_);
  nor _52819_ (_20400_, _20392_, _05634_);
  and _52820_ (_20401_, _20392_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _52821_ (_20402_, _20401_, _20400_);
  or _52822_ (_20403_, _20402_, _20395_);
  and _52823_ (_20404_, _20403_, _20399_);
  or _52824_ (_20405_, _20404_, _20387_);
  and _52825_ (_20406_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _52826_ (_20407_, \oc8051_symbolic_cxrom1.regvalid [6], _26149_);
  or _52827_ (_20408_, _20407_, _26153_);
  or _52828_ (_20409_, _20408_, _20406_);
  or _52829_ (_20410_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _52830_ (_20411_, \oc8051_symbolic_cxrom1.regvalid [10], _26149_);
  and _52831_ (_20412_, _20411_, _20410_);
  or _52832_ (_20413_, _20412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _52833_ (_20414_, _20413_, _20409_);
  and _52834_ (_20415_, _20414_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _52835_ (_20416_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _52836_ (_20417_, \oc8051_symbolic_cxrom1.regvalid [0], _26149_);
  or _52837_ (_20418_, _20417_, _20416_);
  and _52838_ (_20419_, _20418_, _26153_);
  and _52839_ (_20420_, \oc8051_symbolic_cxrom1.regvalid [4], _26149_);
  and _52840_ (_20421_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _52841_ (_20422_, _20421_, _20420_);
  and _52842_ (_20423_, _20422_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _52843_ (_20424_, _20423_, _20419_);
  and _52844_ (_20425_, _20424_, _09640_);
  or _52845_ (_20426_, _20425_, _20415_);
  and _52846_ (_20427_, _20426_, _09731_);
  and _52847_ (_20428_, _20378_, _20422_);
  or _52848_ (_20429_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _52849_ (_20430_, \oc8051_symbolic_cxrom1.regvalid [0], _26149_);
  and _52850_ (_20431_, _20430_, _20357_);
  and _52851_ (_20432_, _20431_, _20429_);
  or _52852_ (_20433_, _20432_, _20428_);
  and _52853_ (_20434_, _20414_, _09640_);
  or _52854_ (_20435_, _20434_, _20433_);
  and _52855_ (_20436_, _20435_, _20427_);
  not _52856_ (_20437_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand _52857_ (_20438_, _20366_, _20437_);
  or _52858_ (_20439_, _20366_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _52859_ (_20440_, _20439_, _20438_);
  and _52860_ (_20441_, _20440_, _20362_);
  not _52861_ (_20442_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nand _52862_ (_20443_, _20366_, _20442_);
  or _52863_ (_20444_, _20366_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _52864_ (_20445_, _20444_, _20361_);
  and _52865_ (_20446_, _20445_, _20443_);
  or _52866_ (_20447_, _20446_, _20441_);
  or _52867_ (_20448_, _20447_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _52868_ (_20449_, _20448_, _20436_);
  and _52869_ (_20450_, _20449_, _20405_);
  and _52870_ (_20451_, _20450_, _20377_);
  or _52871_ (_20452_, \oc8051_symbolic_cxrom1.regvalid [10], _09640_);
  or _52872_ (_20453_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _52873_ (_20454_, _20453_, _20452_);
  nand _52874_ (_20455_, _20454_, _20392_);
  or _52875_ (_20456_, \oc8051_symbolic_cxrom1.regvalid [2], _09640_);
  or _52876_ (_20457_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _52877_ (_20458_, _20457_, _20456_);
  or _52878_ (_20459_, _20458_, _20392_);
  and _52879_ (_20460_, _20459_, _20455_);
  or _52880_ (_20461_, _20460_, _20395_);
  nor _52881_ (_20462_, _20366_, _19774_);
  and _52882_ (_20463_, _20366_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _52883_ (_20464_, _20463_, _20462_);
  and _52884_ (_20465_, _20464_, _20362_);
  or _52885_ (_20466_, _20366_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _52886_ (_20467_, \oc8051_symbolic_cxrom1.regvalid [12], _26149_);
  and _52887_ (_20468_, _20467_, _20361_);
  and _52888_ (_20469_, _20468_, _20466_);
  or _52889_ (_20470_, _20469_, _09640_);
  or _52890_ (_20471_, _20470_, _20465_);
  nand _52891_ (_20472_, \oc8051_symbolic_cxrom1.regvalid [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _52892_ (_20473_, _20472_, _20396_);
  or _52893_ (_20474_, _20473_, _26153_);
  or _52894_ (_20475_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _52895_ (_20476_, \oc8051_symbolic_cxrom1.regvalid [11], _26149_);
  and _52896_ (_20477_, _20476_, _20475_);
  or _52897_ (_20478_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _52898_ (_20479_, _20478_, _20474_);
  and _52899_ (_20480_, _20479_, _20359_);
  and _52900_ (_20481_, _09640_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _52901_ (_20482_, _20381_, _26153_);
  or _52902_ (_20483_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _52903_ (_20484_, \oc8051_symbolic_cxrom1.regvalid [9], _26149_);
  and _52904_ (_20485_, _20484_, _20483_);
  or _52905_ (_20486_, _20485_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _52906_ (_20487_, _20486_, _20482_);
  and _52907_ (_20488_, _20487_, _20481_);
  or _52908_ (_20489_, _20488_, _20480_);
  and _52909_ (_20490_, _20479_, _09640_);
  or _52910_ (_20491_, _20490_, _20387_);
  and _52911_ (_20492_, _20491_, _20489_);
  and _52912_ (_20493_, _20492_, _20471_);
  and _52913_ (_20494_, _20493_, _20461_);
  or _52914_ (_20495_, _20366_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _52915_ (_20496_, \oc8051_symbolic_cxrom1.regvalid [14], _26149_);
  and _52916_ (_20497_, _20496_, _20495_);
  or _52917_ (_20498_, _20497_, _20362_);
  not _52918_ (_20499_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _52919_ (_20500_, _20366_, _20499_);
  or _52920_ (_20501_, _20366_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _52921_ (_20502_, _20501_, _20500_);
  or _52922_ (_20503_, _20502_, _20361_);
  and _52923_ (_20504_, _20503_, _20498_);
  or _52924_ (_20505_, _20504_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _52925_ (_20506_, _20392_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _52926_ (_20507_, _20407_, _09640_);
  or _52927_ (_20508_, _20507_, _20506_);
  and _52928_ (_20509_, _20392_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _52929_ (_20510_, _20420_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _52930_ (_20511_, _20510_, _20509_);
  nand _52931_ (_20512_, _20511_, _20508_);
  nand _52932_ (_20513_, _20512_, _20395_);
  and _52933_ (_20514_, _20513_, _20505_);
  and _52934_ (_20515_, _20514_, _20494_);
  or _52935_ (_20516_, _20515_, _20451_);
  nor _52936_ (_20517_, _19736_, _22752_);
  and _52937_ (_20518_, _20517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52938_ (_20519_, _20517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52939_ (_20520_, _20519_, _20518_);
  nand _52940_ (_20521_, _20520_, _20371_);
  and _52941_ (_20522_, _19736_, _22752_);
  nor _52942_ (_20523_, _20522_, _20517_);
  nor _52943_ (_20524_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _52944_ (_20525_, _20524_);
  and _52945_ (_20526_, _20525_, _20523_);
  and _52946_ (_20527_, _20526_, _20521_);
  nor _52947_ (_20528_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _52948_ (_20529_, _20363_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52949_ (_20530_, _20529_, _20528_);
  and _52950_ (_20531_, _20530_, _22752_);
  or _52951_ (_20532_, _20531_, _20527_);
  and _52952_ (_20533_, _20532_, _19736_);
  nand _52953_ (_20534_, _20520_, _05677_);
  nor _52954_ (_20535_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _52955_ (_20536_, _20535_);
  and _52956_ (_20537_, _20536_, _19738_);
  and _52957_ (_20538_, _20537_, _20534_);
  nand _52958_ (_20539_, _20520_, _20442_);
  nor _52959_ (_20540_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52960_ (_20541_, _20540_, _19757_);
  and _52961_ (_20542_, _20541_, _20539_);
  or _52962_ (_20543_, _20542_, _20538_);
  and _52963_ (_20544_, _20543_, _20523_);
  or _52964_ (_20545_, _20544_, _20533_);
  not _52965_ (_20546_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand _52966_ (_20547_, _20520_, _20546_);
  not _52967_ (_20548_, _20523_);
  nor _52968_ (_20549_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52969_ (_20550_, _20549_, _20548_);
  and _52970_ (_20551_, _20550_, _20547_);
  and _52971_ (_20552_, _20520_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _52972_ (_20553_, _20520_, _19774_);
  or _52973_ (_20554_, _20553_, _20552_);
  and _52974_ (_20555_, _20554_, _20548_);
  or _52975_ (_20556_, _20555_, _20551_);
  and _52976_ (_20557_, _20556_, _19781_);
  and _52977_ (_20558_, _20520_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _52978_ (_20559_, _20520_, _19787_);
  or _52979_ (_20560_, _20559_, _20558_);
  and _52980_ (_20561_, _20560_, _19738_);
  and _52981_ (_20562_, _20520_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _52982_ (_20563_, _20520_, _05653_);
  or _52983_ (_20564_, _20563_, _20562_);
  and _52984_ (_20565_, _20564_, _19756_);
  or _52985_ (_20566_, _20565_, _20561_);
  and _52986_ (_20567_, _20566_, _20548_);
  or _52987_ (_20568_, _20567_, _20557_);
  or _52988_ (_20569_, _20568_, _20545_);
  and _52989_ (_20570_, _05677_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52990_ (_20571_, _20570_, _22752_);
  and _52991_ (_20572_, _20571_, _20536_);
  and _52992_ (_20573_, _20499_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52993_ (_20574_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52994_ (_20575_, _20574_, _20573_);
  and _52995_ (_20576_, _20575_, _22752_);
  nor _52996_ (_20577_, _20576_, _20572_);
  nor _52997_ (_20578_, _20577_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _52998_ (_20579_, _20546_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _52999_ (_20580_, _20579_, _20549_);
  and _53000_ (_20581_, _20580_, _20110_);
  and _53001_ (_20582_, _19774_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53002_ (_20583_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53003_ (_20584_, _20583_, _22752_);
  nor _53004_ (_20585_, _20584_, _20582_);
  and _53005_ (_20586_, _20585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _53006_ (_20587_, _20586_, _20581_);
  not _53007_ (_20588_, _20587_);
  nor _53008_ (_20589_, _20588_, _20578_);
  nor _53009_ (_20590_, _20589_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _53010_ (_20591_, _20590_);
  and _53011_ (_20592_, _20371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53012_ (_20593_, _20592_, _22752_);
  and _53013_ (_20594_, _20593_, _20525_);
  nor _53014_ (_20595_, _20594_, _20531_);
  nor _53015_ (_20596_, _20595_, _19782_);
  not _53016_ (_20597_, _19739_);
  and _53017_ (_20598_, \oc8051_symbolic_cxrom1.regvalid [9], _22758_);
  and _53018_ (_20599_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53019_ (_20600_, _20599_, _20598_);
  nor _53020_ (_20601_, _20600_, _20597_);
  and _53021_ (_20602_, _19738_, _22752_);
  and _53022_ (_20603_, _20442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53023_ (_20604_, _20603_, _20540_);
  and _53024_ (_20605_, _20604_, _20602_);
  nor _53025_ (_20606_, _20605_, _20601_);
  not _53026_ (_20607_, _20606_);
  nor _53027_ (_20608_, _20607_, _20596_);
  and _53028_ (_20609_, _20608_, _20591_);
  and _53029_ (_20610_, _20604_, _20111_);
  nor _53030_ (_20611_, _20610_, _22742_);
  nor _53031_ (_20612_, _20595_, _22747_);
  nor _53032_ (_20613_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _53033_ (_20614_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _53034_ (_20615_, _20437_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53035_ (_20616_, _20615_, _20614_);
  and _53036_ (_20617_, _20616_, _20613_);
  nor _53037_ (_20618_, _20617_, _20612_);
  and _53038_ (_20619_, _20618_, _20611_);
  nor _53039_ (_20620_, _20577_, _22747_);
  nor _53040_ (_20621_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53041_ (_20622_, \oc8051_symbolic_cxrom1.regvalid [8], _22758_);
  nor _53042_ (_20623_, _20622_, _20621_);
  and _53043_ (_20624_, _20623_, _20613_);
  and _53044_ (_20625_, _20580_, _20111_);
  or _53045_ (_20626_, _20625_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _53046_ (_20627_, _20626_, _20624_);
  nor _53047_ (_20628_, _20627_, _20620_);
  nor _53048_ (_20629_, _20628_, _20619_);
  not _53049_ (_20630_, _22740_);
  nor _53050_ (_20631_, _20630_, first_instr);
  nand _53051_ (_20632_, _20631_, _20629_);
  or _53052_ (_20633_, _20632_, _20609_);
  nor _53053_ (_20634_, _20633_, _19795_);
  and _53054_ (_20635_, _20634_, _20569_);
  and _53055_ (_20636_, _20635_, _20516_);
  nor _53056_ (_20637_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53057_ (_20638_, _07573_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53058_ (_20639_, _20638_, _20637_);
  and _53059_ (_20640_, _20639_, _20613_);
  or _53060_ (_20641_, _20640_, _22758_);
  nor _53061_ (_20642_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53062_ (_20643_, _08484_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53063_ (_20644_, _20643_, _20642_);
  and _53064_ (_20645_, _20644_, _19834_);
  nor _53065_ (_20646_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53066_ (_20647_, _08117_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53067_ (_20648_, _20647_, _20646_);
  and _53068_ (_20649_, _20648_, _20111_);
  nor _53069_ (_20650_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53070_ (_20651_, _07816_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53071_ (_20652_, _20651_, _20650_);
  and _53072_ (_20653_, _20652_, _20110_);
  or _53073_ (_20654_, _20653_, _20649_);
  or _53074_ (_20655_, _20654_, _20645_);
  or _53075_ (_20656_, _20655_, _20641_);
  nor _53076_ (_20657_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53077_ (_20658_, _07046_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53078_ (_20659_, _20658_, _20657_);
  and _53079_ (_20660_, _20659_, _20111_);
  nor _53080_ (_20661_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53081_ (_20662_, _07310_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53082_ (_20663_, _20662_, _20661_);
  and _53083_ (_20664_, _20663_, _19834_);
  or _53084_ (_20665_, _20664_, _20660_);
  nor _53085_ (_20666_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53086_ (_20667_, _06545_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53087_ (_20668_, _20667_, _20666_);
  and _53088_ (_20669_, _20668_, _20613_);
  nor _53089_ (_20670_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53090_ (_20671_, _06790_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53091_ (_20672_, _20671_, _20670_);
  and _53092_ (_20673_, _20672_, _20110_);
  or _53093_ (_20674_, _20673_, _20669_);
  or _53094_ (_20675_, _20674_, _20665_);
  or _53095_ (_20676_, _20675_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _53096_ (_20677_, _20676_, _20656_);
  and _53097_ (_20678_, _20677_, _20629_);
  nor _53098_ (_20679_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53099_ (_20680_, _07294_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53100_ (_20681_, _20680_, _20679_);
  and _53101_ (_20682_, _20681_, _19834_);
  nor _53102_ (_20683_, _20682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53103_ (_20684_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53104_ (_20685_, _06518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53105_ (_20686_, _20685_, _20684_);
  and _53106_ (_20687_, _20686_, _20613_);
  not _53107_ (_20688_, _20687_);
  nor _53108_ (_20689_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53109_ (_20690_, _06775_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53110_ (_20691_, _20690_, _20689_);
  and _53111_ (_20692_, _20691_, _20110_);
  nor _53112_ (_20693_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53113_ (_20694_, _07023_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53114_ (_20695_, _20694_, _20693_);
  and _53115_ (_20696_, _20695_, _20111_);
  nor _53116_ (_20697_, _20696_, _20692_);
  and _53117_ (_20698_, _20697_, _20688_);
  and _53118_ (_20699_, _20698_, _20683_);
  nor _53119_ (_20700_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53120_ (_20701_, _08472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53121_ (_20702_, _20701_, _20700_);
  and _53122_ (_20703_, _20702_, _19834_);
  nor _53123_ (_20704_, _20703_, _22758_);
  nor _53124_ (_20705_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53125_ (_20706_, _07795_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53126_ (_20707_, _20706_, _20705_);
  and _53127_ (_20708_, _20707_, _20110_);
  not _53128_ (_20709_, _20708_);
  nor _53129_ (_20710_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53130_ (_20711_, _08104_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53131_ (_20712_, _20711_, _20710_);
  and _53132_ (_20713_, _20712_, _20111_);
  nor _53133_ (_20714_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53134_ (_20715_, _07556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53135_ (_20716_, _20715_, _20714_);
  and _53136_ (_20717_, _20716_, _20613_);
  nor _53137_ (_20718_, _20717_, _20713_);
  and _53138_ (_20719_, _20718_, _20709_);
  and _53139_ (_20720_, _20719_, _20704_);
  nor _53140_ (_20721_, _20720_, _20699_);
  and _53141_ (_20722_, _20721_, _20629_);
  nor _53142_ (_20723_, _20722_, _20678_);
  nor _53143_ (_20724_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53144_ (_20725_, _08179_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53145_ (_20726_, _20725_, _20724_);
  and _53146_ (_20727_, _20726_, _20111_);
  nor _53147_ (_20728_, _20727_, _22758_);
  nor _53148_ (_20729_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53149_ (_20730_, _07631_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53150_ (_20731_, _20730_, _20729_);
  and _53151_ (_20732_, _20731_, _20613_);
  nor _53152_ (_20733_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53153_ (_20734_, _07869_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53154_ (_20735_, _20734_, _20733_);
  and _53155_ (_20736_, _20735_, _20110_);
  nor _53156_ (_20737_, _20736_, _20732_);
  nor _53157_ (_20738_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53158_ (_20739_, _08547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53159_ (_20740_, _20739_, _20738_);
  and _53160_ (_20741_, _20740_, _19834_);
  not _53161_ (_20742_, _20741_);
  and _53162_ (_20743_, _20742_, _20737_);
  and _53163_ (_20744_, _20743_, _20728_);
  nor _53164_ (_20745_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53165_ (_20746_, _07112_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53166_ (_20747_, _20746_, _20745_);
  and _53167_ (_20748_, _20747_, _20111_);
  nor _53168_ (_20749_, _20748_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53169_ (_20750_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53170_ (_20751_, _06609_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53171_ (_20752_, _20751_, _20750_);
  and _53172_ (_20753_, _20752_, _20613_);
  nor _53173_ (_20754_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53174_ (_20755_, _06845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53175_ (_20756_, _20755_, _20754_);
  and _53176_ (_20757_, _20756_, _20110_);
  nor _53177_ (_20758_, _20757_, _20753_);
  nor _53178_ (_20759_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53179_ (_20760_, _07375_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53180_ (_20761_, _20760_, _20759_);
  and _53181_ (_20762_, _20761_, _19834_);
  not _53182_ (_20763_, _20762_);
  and _53183_ (_20764_, _20763_, _20758_);
  and _53184_ (_20765_, _20764_, _20749_);
  nor _53185_ (_20766_, _20765_, _20744_);
  and _53186_ (_20767_, _20766_, _20629_);
  nor _53187_ (_20768_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53188_ (_20769_, _08528_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53189_ (_20770_, _20769_, _20768_);
  and _53190_ (_20771_, _20770_, _19834_);
  nor _53191_ (_20772_, _20771_, _22758_);
  nor _53192_ (_20773_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53193_ (_20774_, _07616_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53194_ (_20775_, _20774_, _20773_);
  and _53195_ (_20776_, _20775_, _20613_);
  not _53196_ (_20777_, _20776_);
  nor _53197_ (_20778_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53198_ (_20779_, _07854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53199_ (_20780_, _20779_, _20778_);
  and _53200_ (_20781_, _20780_, _20110_);
  nor _53201_ (_20782_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53202_ (_20783_, _08162_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53203_ (_20784_, _20783_, _20782_);
  and _53204_ (_20785_, _20784_, _20111_);
  nor _53205_ (_20786_, _20785_, _20781_);
  and _53206_ (_20787_, _20786_, _20777_);
  and _53207_ (_20788_, _20787_, _20772_);
  nor _53208_ (_20789_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53209_ (_20790_, _07357_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53210_ (_20791_, _20790_, _20789_);
  and _53211_ (_20792_, _20791_, _19834_);
  nor _53212_ (_20793_, _20792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53213_ (_20794_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53214_ (_20795_, _06594_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53215_ (_20796_, _20795_, _20794_);
  and _53216_ (_20797_, _20796_, _20613_);
  not _53217_ (_20798_, _20797_);
  nor _53218_ (_20799_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53219_ (_20800_, _06832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53220_ (_20801_, _20800_, _20799_);
  and _53221_ (_20802_, _20801_, _20110_);
  nor _53222_ (_20803_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53223_ (_20804_, _07096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53224_ (_20805_, _20804_, _20803_);
  and _53225_ (_20806_, _20805_, _20111_);
  nor _53226_ (_20807_, _20806_, _20802_);
  and _53227_ (_20808_, _20807_, _20798_);
  and _53228_ (_20809_, _20808_, _20793_);
  nor _53229_ (_20810_, _20809_, _20788_);
  and _53230_ (_20811_, _20810_, _20629_);
  nor _53231_ (_20812_, _20811_, _20767_);
  and _53232_ (_20813_, _20812_, _20723_);
  nor _53233_ (_20814_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53234_ (_20815_, _06804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53235_ (_20816_, _20815_, _20814_);
  and _53236_ (_20817_, _20816_, _20110_);
  nor _53237_ (_20818_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53238_ (_20819_, _07063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53239_ (_20820_, _20819_, _20818_);
  and _53240_ (_20821_, _20820_, _20111_);
  nor _53241_ (_20822_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53242_ (_20823_, _06562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53243_ (_20824_, _20823_, _20822_);
  and _53244_ (_20825_, _20824_, _20613_);
  nor _53245_ (_20826_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53246_ (_20827_, _07329_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53247_ (_20828_, _20827_, _20826_);
  and _53248_ (_20829_, _20828_, _19834_);
  or _53249_ (_20830_, _20829_, _20825_);
  or _53250_ (_20831_, _20830_, _20821_);
  or _53251_ (_20832_, _20831_, _20817_);
  and _53252_ (_20833_, _20832_, _22758_);
  nor _53253_ (_20834_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53254_ (_20835_, _07828_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53255_ (_20836_, _20835_, _20834_);
  and _53256_ (_20837_, _20836_, _20110_);
  nor _53257_ (_20838_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53258_ (_20839_, _08134_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53259_ (_20840_, _20839_, _20838_);
  and _53260_ (_20841_, _20840_, _20111_);
  nor _53261_ (_20842_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53262_ (_20843_, _07590_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53263_ (_20844_, _20843_, _20842_);
  and _53264_ (_20845_, _20844_, _20613_);
  nor _53265_ (_20846_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53266_ (_20847_, _08498_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53267_ (_20848_, _20847_, _20846_);
  and _53268_ (_20849_, _20848_, _19834_);
  or _53269_ (_20850_, _20849_, _20845_);
  or _53270_ (_20851_, _20850_, _20841_);
  or _53271_ (_20852_, _20851_, _20837_);
  and _53272_ (_20853_, _20852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53273_ (_20854_, _20853_, _20833_);
  and _53274_ (_20855_, _20854_, _20629_);
  nor _53275_ (_20856_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53276_ (_20857_, _06818_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53277_ (_20858_, _20857_, _20856_);
  and _53278_ (_20859_, _20858_, _20110_);
  nor _53279_ (_20860_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53280_ (_20861_, _07078_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53281_ (_20862_, _20861_, _20860_);
  and _53282_ (_20863_, _20862_, _20111_);
  nor _53283_ (_20864_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53284_ (_20865_, _06578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53285_ (_20866_, _20865_, _20864_);
  and _53286_ (_20867_, _20866_, _20613_);
  nor _53287_ (_20868_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53288_ (_20869_, _07339_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53289_ (_20870_, _20869_, _20868_);
  and _53290_ (_20871_, _20870_, _19834_);
  or _53291_ (_20872_, _20871_, _20867_);
  or _53292_ (_20873_, _20872_, _20863_);
  or _53293_ (_20874_, _20873_, _20859_);
  and _53294_ (_20875_, _20874_, _22758_);
  nor _53295_ (_20876_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53296_ (_20877_, _07840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53297_ (_20878_, _20877_, _20876_);
  and _53298_ (_20879_, _20878_, _20110_);
  nor _53299_ (_20880_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53300_ (_20881_, _08148_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53301_ (_20882_, _20881_, _20880_);
  and _53302_ (_20883_, _20882_, _20111_);
  nor _53303_ (_20884_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53304_ (_20885_, _07602_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53305_ (_20886_, _20885_, _20884_);
  and _53306_ (_20887_, _20886_, _20613_);
  nor _53307_ (_20888_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53308_ (_20889_, _08512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53309_ (_20890_, _20889_, _20888_);
  and _53310_ (_20891_, _20890_, _19834_);
  or _53311_ (_20892_, _20891_, _20887_);
  or _53312_ (_20893_, _20892_, _20883_);
  or _53313_ (_20894_, _20893_, _20879_);
  and _53314_ (_20895_, _20894_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53315_ (_20896_, _20895_, _20875_);
  and _53316_ (_20897_, _20896_, _20629_);
  nor _53317_ (_20898_, _20897_, _20855_);
  nor _53318_ (_20899_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53319_ (_20900_, _06857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53320_ (_20901_, _20900_, _20899_);
  and _53321_ (_20902_, _20901_, _20110_);
  nor _53322_ (_20903_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53323_ (_20904_, _07127_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53324_ (_20905_, _20904_, _20903_);
  and _53325_ (_20906_, _20905_, _20111_);
  nor _53326_ (_20907_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53327_ (_20908_, _07384_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53328_ (_20909_, _20908_, _20907_);
  and _53329_ (_20910_, _20909_, _19834_);
  nor _53330_ (_20911_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53331_ (_20912_, _06625_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53332_ (_20913_, _20912_, _20911_);
  and _53333_ (_20914_, _20913_, _20613_);
  or _53334_ (_20915_, _20914_, _20910_);
  or _53335_ (_20916_, _20915_, _20906_);
  or _53336_ (_20917_, _20916_, _20902_);
  and _53337_ (_20918_, _20917_, _22758_);
  nor _53338_ (_20919_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53339_ (_20920_, _07887_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53340_ (_20921_, _20920_, _20919_);
  and _53341_ (_20922_, _20921_, _20110_);
  nor _53342_ (_20923_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53343_ (_20924_, _08192_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53344_ (_20925_, _20924_, _20923_);
  and _53345_ (_20926_, _20925_, _20111_);
  nor _53346_ (_20927_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53347_ (_20928_, _08564_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53348_ (_20929_, _20928_, _20927_);
  and _53349_ (_20930_, _20929_, _19834_);
  nor _53350_ (_20931_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53351_ (_20932_, _07647_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53352_ (_20933_, _20932_, _20931_);
  and _53353_ (_20934_, _20933_, _20613_);
  or _53354_ (_20935_, _20934_, _20930_);
  or _53355_ (_20936_, _20935_, _20926_);
  or _53356_ (_20937_, _20936_, _20922_);
  and _53357_ (_20938_, _20937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53358_ (_20939_, _20938_, _20918_);
  and _53359_ (_20940_, _20939_, _20629_);
  not _53360_ (_20941_, _20940_);
  nor _53361_ (_20942_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53362_ (_20943_, _05704_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53363_ (_20944_, _20943_, _20942_);
  and _53364_ (_20945_, _20944_, _20111_);
  nor _53365_ (_20946_, _20945_, _22758_);
  nor _53366_ (_20947_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53367_ (_20948_, _05709_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53368_ (_20949_, _20948_, _20947_);
  and _53369_ (_20950_, _20949_, _20613_);
  nor _53370_ (_20951_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53371_ (_20952_, _05697_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53372_ (_20953_, _20952_, _20951_);
  and _53373_ (_20954_, _20953_, _20110_);
  nor _53374_ (_20955_, _20954_, _20950_);
  nor _53375_ (_20956_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53376_ (_20957_, _05691_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53377_ (_20958_, _20957_, _20956_);
  and _53378_ (_20959_, _20958_, _19834_);
  not _53379_ (_20960_, _20959_);
  and _53380_ (_20961_, _20960_, _20955_);
  and _53381_ (_20962_, _20961_, _20946_);
  nor _53382_ (_20963_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53383_ (_20964_, _05732_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53384_ (_20965_, _20964_, _20963_);
  and _53385_ (_20966_, _20965_, _20111_);
  nor _53386_ (_20967_, _20966_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53387_ (_20968_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53388_ (_20969_, _05737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53389_ (_20970_, _20969_, _20968_);
  and _53390_ (_20971_, _20970_, _20613_);
  nor _53391_ (_20972_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53392_ (_20973_, _05719_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53393_ (_20974_, _20973_, _20972_);
  and _53394_ (_20975_, _20974_, _20110_);
  nor _53395_ (_20976_, _20975_, _20971_);
  nor _53396_ (_20977_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53397_ (_20978_, _05726_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53398_ (_20979_, _20978_, _20977_);
  and _53399_ (_20980_, _20979_, _19834_);
  not _53400_ (_20981_, _20980_);
  and _53401_ (_20982_, _20981_, _20976_);
  and _53402_ (_20983_, _20982_, _20967_);
  nor _53403_ (_20984_, _20983_, _20962_);
  and _53404_ (_20985_, _20984_, _20629_);
  and _53405_ (_20986_, _20985_, _20941_);
  and _53406_ (_20987_, _20986_, _20898_);
  and _53407_ (_20988_, _20987_, _20813_);
  and _53408_ (_20989_, _20988_, _20636_);
  and _53409_ (_20990_, _20989_, _20356_);
  and _53410_ (_20991_, _20695_, _20110_);
  or _53411_ (_20992_, _20991_, _20029_);
  and _53412_ (_20993_, _20686_, _19834_);
  and _53413_ (_20994_, _20691_, _20613_);
  and _53414_ (_20995_, _20681_, _20111_);
  or _53415_ (_20996_, _20995_, _20994_);
  or _53416_ (_20997_, _20996_, _20993_);
  or _53417_ (_20998_, _20997_, _20992_);
  and _53418_ (_20999_, _20712_, _20110_);
  or _53419_ (_21000_, _20999_, _20028_);
  and _53420_ (_21001_, _20707_, _20613_);
  and _53421_ (_21002_, _20702_, _20111_);
  and _53422_ (_21003_, _20716_, _19834_);
  or _53423_ (_21004_, _21003_, _21002_);
  or _53424_ (_21005_, _21004_, _21001_);
  or _53425_ (_21006_, _21005_, _21000_);
  nand _53426_ (_21007_, _21006_, _20998_);
  nor _53427_ (_21008_, _21007_, _20609_);
  nor _53428_ (_21009_, _21008_, _09731_);
  and _53429_ (_21010_, _21008_, _09731_);
  or _53430_ (_21011_, _21010_, _21009_);
  not _53431_ (_21012_, _20609_);
  and _53432_ (_21013_, _20659_, _20110_);
  and _53433_ (_21014_, _20663_, _20111_);
  nor _53434_ (_21015_, _21014_, _21013_);
  and _53435_ (_21016_, _20668_, _19834_);
  and _53436_ (_21017_, _20672_, _20613_);
  nor _53437_ (_21018_, _21017_, _21016_);
  and _53438_ (_21019_, _21018_, _21015_);
  and _53439_ (_21020_, _21019_, _20028_);
  and _53440_ (_21021_, _20644_, _20111_);
  and _53441_ (_21022_, _20639_, _19834_);
  and _53442_ (_21023_, _20648_, _20110_);
  or _53443_ (_21024_, _21023_, _21022_);
  nor _53444_ (_21025_, _21024_, _21021_);
  and _53445_ (_21026_, _20652_, _20613_);
  nor _53446_ (_21027_, _21026_, _20028_);
  and _53447_ (_21028_, _21027_, _21025_);
  nor _53448_ (_21029_, _21028_, _21020_);
  and _53449_ (_21030_, _21029_, _21012_);
  nor _53450_ (_21031_, _21030_, _09640_);
  and _53451_ (_21032_, _21030_, _09640_);
  or _53452_ (_21033_, _21032_, _21031_);
  or _53453_ (_21034_, _21033_, _21011_);
  and _53454_ (_21035_, _20878_, _20613_);
  and _53455_ (_21036_, _20890_, _20111_);
  and _53456_ (_21037_, _20882_, _20110_);
  and _53457_ (_21038_, _20886_, _19834_);
  or _53458_ (_21039_, _21038_, _21037_);
  or _53459_ (_21040_, _21039_, _21036_);
  or _53460_ (_21041_, _21040_, _21035_);
  and _53461_ (_21042_, _21041_, _20029_);
  and _53462_ (_21043_, _20858_, _20613_);
  and _53463_ (_21044_, _20870_, _20111_);
  and _53464_ (_21045_, _20866_, _19834_);
  and _53465_ (_21046_, _20862_, _20110_);
  or _53466_ (_21047_, _21046_, _21045_);
  or _53467_ (_21048_, _21047_, _21044_);
  or _53468_ (_21049_, _21048_, _21043_);
  and _53469_ (_21050_, _21049_, _20028_);
  or _53470_ (_21051_, _21050_, _21042_);
  and _53471_ (_21052_, _21051_, _21012_);
  nand _53472_ (_21053_, _21052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53473_ (_21054_, _21052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53474_ (_21055_, _21054_, _21053_);
  and _53475_ (_21056_, _20836_, _20613_);
  and _53476_ (_21057_, _20848_, _20111_);
  and _53477_ (_21058_, _20844_, _19834_);
  and _53478_ (_21059_, _20840_, _20110_);
  or _53479_ (_21060_, _21059_, _21058_);
  or _53480_ (_21061_, _21060_, _21057_);
  or _53481_ (_21062_, _21061_, _21056_);
  and _53482_ (_21063_, _21062_, _20029_);
  and _53483_ (_21064_, _20816_, _20613_);
  and _53484_ (_21065_, _20828_, _20111_);
  and _53485_ (_21066_, _20824_, _19834_);
  and _53486_ (_21067_, _20820_, _20110_);
  or _53487_ (_21068_, _21067_, _21066_);
  or _53488_ (_21069_, _21068_, _21065_);
  or _53489_ (_21070_, _21069_, _21064_);
  and _53490_ (_21071_, _21070_, _20028_);
  or _53491_ (_21072_, _21071_, _21063_);
  and _53492_ (_21073_, _21072_, _21012_);
  nor _53493_ (_21074_, _21073_, _26153_);
  and _53494_ (_21075_, _21073_, _26153_);
  or _53495_ (_21076_, _21075_, _21074_);
  or _53496_ (_21077_, _21076_, _21055_);
  or _53497_ (_21078_, _21077_, _21034_);
  and _53498_ (_21079_, _20958_, _20111_);
  and _53499_ (_21080_, _20944_, _20110_);
  nor _53500_ (_21081_, _21080_, _21079_);
  and _53501_ (_21082_, _20949_, _19834_);
  and _53502_ (_21083_, _20953_, _20613_);
  nor _53503_ (_21084_, _21083_, _21082_);
  and _53504_ (_21085_, _21084_, _21081_);
  and _53505_ (_21086_, _21085_, _20029_);
  and _53506_ (_21087_, _20979_, _20111_);
  and _53507_ (_21088_, _20970_, _19834_);
  and _53508_ (_21089_, _20965_, _20110_);
  or _53509_ (_21090_, _21089_, _21088_);
  nor _53510_ (_21091_, _21090_, _21087_);
  and _53511_ (_21092_, _20974_, _20613_);
  nor _53512_ (_21093_, _21092_, _20029_);
  and _53513_ (_21094_, _21093_, _21091_);
  nor _53514_ (_21095_, _21094_, _21086_);
  and _53515_ (_21096_, _21095_, _21012_);
  nand _53516_ (_21097_, _21096_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or _53517_ (_21098_, _21096_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _53518_ (_21099_, _21098_, _21097_);
  and _53519_ (_21100_, _20905_, _20110_);
  and _53520_ (_21101_, _20909_, _20111_);
  and _53521_ (_21102_, _20913_, _19834_);
  or _53522_ (_21103_, _21102_, _21101_);
  or _53523_ (_21104_, _21103_, _21100_);
  and _53524_ (_21105_, _20901_, _20613_);
  or _53525_ (_21106_, _21105_, _20029_);
  or _53526_ (_21107_, _21106_, _21104_);
  and _53527_ (_21108_, _20925_, _20110_);
  or _53528_ (_21109_, _21108_, _20028_);
  and _53529_ (_21110_, _20933_, _19834_);
  and _53530_ (_21111_, _20921_, _20613_);
  and _53531_ (_21112_, _20929_, _20111_);
  or _53532_ (_21113_, _21112_, _21111_);
  or _53533_ (_21114_, _21113_, _21110_);
  or _53534_ (_21115_, _21114_, _21109_);
  nand _53535_ (_21116_, _21115_, _21107_);
  nor _53536_ (_21117_, _21116_, _20609_);
  nand _53537_ (_21118_, _21117_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or _53538_ (_21119_, _21117_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _53539_ (_21120_, _21119_, _21118_);
  or _53540_ (_21121_, _21120_, _21099_);
  and _53541_ (_21122_, _20747_, _20110_);
  or _53542_ (_21123_, _21122_, _20029_);
  and _53543_ (_21124_, _20752_, _19834_);
  and _53544_ (_21125_, _20756_, _20613_);
  and _53545_ (_21126_, _20761_, _20111_);
  or _53546_ (_21127_, _21126_, _21125_);
  or _53547_ (_21128_, _21127_, _21124_);
  or _53548_ (_21129_, _21128_, _21123_);
  and _53549_ (_21130_, _20740_, _20111_);
  or _53550_ (_21131_, _21130_, _20028_);
  and _53551_ (_21132_, _20735_, _20613_);
  and _53552_ (_21133_, _20731_, _19834_);
  or _53553_ (_21134_, _21133_, _21132_);
  and _53554_ (_21135_, _20726_, _20110_);
  or _53555_ (_21136_, _21135_, _21134_);
  or _53556_ (_21137_, _21136_, _21131_);
  nand _53557_ (_21138_, _21137_, _21129_);
  nor _53558_ (_21139_, _21138_, _20609_);
  nand _53559_ (_21140_, _21139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or _53560_ (_21141_, _21139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _53561_ (_21142_, _21141_, _21140_);
  and _53562_ (_21143_, _20805_, _20110_);
  or _53563_ (_21144_, _21143_, _20029_);
  and _53564_ (_21145_, _20796_, _19834_);
  and _53565_ (_21146_, _20801_, _20613_);
  and _53566_ (_21147_, _20791_, _20111_);
  or _53567_ (_21148_, _21147_, _21146_);
  or _53568_ (_21149_, _21148_, _21145_);
  or _53569_ (_21150_, _21149_, _21144_);
  and _53570_ (_21151_, _20784_, _20110_);
  or _53571_ (_21152_, _21151_, _20028_);
  and _53572_ (_21153_, _20775_, _19834_);
  and _53573_ (_21154_, _20780_, _20613_);
  and _53574_ (_21155_, _20770_, _20111_);
  or _53575_ (_21156_, _21155_, _21154_);
  or _53576_ (_21157_, _21156_, _21153_);
  or _53577_ (_21158_, _21157_, _21152_);
  nand _53578_ (_21159_, _21158_, _21150_);
  nor _53579_ (_21160_, _21159_, _20609_);
  nor _53580_ (_21161_, _21160_, _22762_);
  and _53581_ (_21162_, _21160_, _22762_);
  or _53582_ (_21163_, _21162_, _21161_);
  or _53583_ (_21164_, _21163_, _21142_);
  or _53584_ (_21165_, _21164_, _21121_);
  or _53585_ (_21166_, _21165_, _21078_);
  nor _53586_ (_21167_, _20152_, _26128_);
  and _53587_ (_21168_, _20152_, _26128_);
  or _53588_ (_21169_, _21168_, _21167_);
  and _53589_ (_21170_, _20191_, _22780_);
  nor _53590_ (_21171_, _20191_, _22780_);
  or _53591_ (_21172_, _21171_, _21170_);
  or _53592_ (_21173_, _21172_, _21169_);
  or _53593_ (_21174_, _20067_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _53594_ (_21175_, _20067_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _53595_ (_21176_, _21175_, _21174_);
  nor _53596_ (_21177_, _20109_, _22789_);
  and _53597_ (_21178_, _20109_, _22789_);
  or _53598_ (_21179_, _21178_, _21177_);
  or _53599_ (_21180_, _21179_, _21176_);
  or _53600_ (_21181_, _21180_, _21173_);
  or _53601_ (_21182_, _19979_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _53602_ (_21183_, _19979_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _53603_ (_21184_, _21183_, _21182_);
  and _53604_ (_21185_, _20022_, _22797_);
  nor _53605_ (_21186_, _20022_, _22797_);
  or _53606_ (_21187_, _21186_, _21185_);
  or _53607_ (_21188_, _21187_, _21184_);
  nor _53608_ (_21189_, _19833_, _04912_);
  and _53609_ (_21190_, _19833_, _04912_);
  or _53610_ (_21191_, _21190_, _21189_);
  nor _53611_ (_21192_, _19935_, _22806_);
  and _53612_ (_21193_, _19935_, _22806_);
  or _53613_ (_21194_, _21193_, _21192_);
  or _53614_ (_21195_, _21194_, _21191_);
  or _53615_ (_21196_, _21195_, _21188_);
  or _53616_ (_21197_, _21196_, _21181_);
  or _53617_ (_21198_, _21197_, _21166_);
  nor _53618_ (_21199_, _20985_, _20940_);
  not _53619_ (_21200_, _20767_);
  not _53620_ (_21201_, _20722_);
  and _53621_ (_21202_, _20898_, _21201_);
  and _53622_ (_21203_, _21202_, _20678_);
  and _53623_ (_21204_, _21203_, _21200_);
  and _53624_ (_21205_, _21204_, _21199_);
  and _53625_ (_21206_, _21205_, _20636_);
  and _53626_ (_21207_, _21206_, _21198_);
  nor _53627_ (_21208_, _20152_, _09640_);
  and _53628_ (_21209_, _20152_, _09640_);
  or _53629_ (_21210_, _21209_, _21208_);
  nor _53630_ (_21211_, _19935_, _22772_);
  nor _53631_ (_21212_, _20767_, _22780_);
  and _53632_ (_21213_, _20767_, _22780_);
  or _53633_ (_21214_, _21213_, _21212_);
  nor _53634_ (_21215_, _20940_, _26128_);
  and _53635_ (_21216_, _20940_, _26128_);
  or _53636_ (_21217_, _21216_, _21215_);
  or _53637_ (_21218_, _21217_, _21214_);
  or _53638_ (_21219_, _19864_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _53639_ (_21220_, _19864_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _53640_ (_21221_, _21220_, _21219_);
  and _53641_ (_21222_, _20985_, _22789_);
  nor _53642_ (_21223_, _20985_, _22789_);
  or _53643_ (_21224_, _21223_, _21222_);
  or _53644_ (_21225_, _21224_, _21221_);
  or _53645_ (_21226_, _21225_, _21218_);
  or _53646_ (_21227_, _21226_, _21211_);
  or _53647_ (_21228_, _21227_, _21210_);
  and _53648_ (_21229_, _20022_, _22762_);
  nor _53649_ (_21230_, _20022_, _22762_);
  or _53650_ (_21231_, _21230_, _21229_);
  nor _53651_ (_21232_, _19859_, _22797_);
  and _53652_ (_21233_, _19859_, _22797_);
  or _53653_ (_21234_, _21233_, _21232_);
  or _53654_ (_21235_, _21234_, _20261_);
  and _53655_ (_21236_, _19848_, _22806_);
  nor _53656_ (_21237_, _19848_, _22806_);
  or _53657_ (_21238_, _21237_, _21236_);
  or _53658_ (_21239_, _21238_, _20245_);
  or _53659_ (_21240_, _21239_, _21235_);
  or _53660_ (_21241_, _21240_, _21231_);
  or _53661_ (_21242_, _21241_, _21228_);
  and _53662_ (_21243_, _19935_, _22772_);
  and _53663_ (_21244_, _19833_, _26136_);
  nor _53664_ (_21245_, _19833_, _26136_);
  or _53665_ (_21246_, _21245_, _21244_);
  or _53666_ (_21247_, _21246_, _21243_);
  nor _53667_ (_21248_, _20067_, _26149_);
  and _53668_ (_21249_, _20109_, _26153_);
  or _53669_ (_21250_, _21249_, _21248_);
  and _53670_ (_21251_, _20067_, _26149_);
  nor _53671_ (_21252_, _19979_, _22767_);
  or _53672_ (_21253_, _21252_, _21251_);
  or _53673_ (_21254_, _21253_, _21250_);
  and _53674_ (_21255_, _20191_, _09731_);
  nor _53675_ (_21256_, _20109_, _26153_);
  or _53676_ (_21257_, _21256_, _21255_);
  nor _53677_ (_21258_, _20191_, _09731_);
  and _53678_ (_21259_, _19979_, _22767_);
  or _53679_ (_21260_, _21259_, _21258_);
  or _53680_ (_21261_, _21260_, _21257_);
  or _53681_ (_21262_, _21261_, _21254_);
  or _53682_ (_21263_, _21262_, _21247_);
  or _53683_ (_21264_, _21263_, _21242_);
  not _53684_ (_21265_, _20678_);
  and _53685_ (_21266_, _20722_, _21265_);
  and _53686_ (_21267_, _21266_, _20898_);
  and _53687_ (_21268_, _21267_, _21264_);
  not _53688_ (_21269_, _20985_);
  and _53689_ (_21270_, _20855_, _20678_);
  and _53690_ (_21271_, _21270_, _20811_);
  and _53691_ (_21272_, _21271_, _20767_);
  not _53692_ (_21273_, _20896_);
  and _53693_ (_21274_, _21273_, _20855_);
  and _53694_ (_21275_, _21274_, _20723_);
  and _53695_ (_21276_, _20811_, _20766_);
  and _53696_ (_21277_, _21276_, _20896_);
  or _53697_ (_21278_, _21277_, _21275_);
  or _53698_ (_21279_, _21278_, _21203_);
  or _53699_ (_21280_, _21279_, _21272_);
  and _53700_ (_21281_, _21280_, _20940_);
  and _53701_ (_21282_, _21274_, _21265_);
  and _53702_ (_21283_, _20941_, _20767_);
  and _53703_ (_21284_, _21283_, _21282_);
  and _53704_ (_21285_, _21282_, _20722_);
  and _53705_ (_21286_, _21285_, _21200_);
  or _53706_ (_21287_, _21286_, _21284_);
  or _53707_ (_21288_, _21287_, _21281_);
  and _53708_ (_21289_, _21288_, _21269_);
  and _53709_ (_21290_, _20940_, _21200_);
  and _53710_ (_21291_, _21290_, _21202_);
  or _53711_ (_21292_, _21291_, _21204_);
  not _53712_ (_21293_, _20766_);
  and _53713_ (_21294_, _20811_, _21293_);
  and _53714_ (_21295_, _21282_, _21294_);
  and _53715_ (_21296_, _21202_, _20766_);
  not _53716_ (_21297_, _20810_);
  and _53717_ (_21298_, _20897_, _21297_);
  not _53718_ (_21299_, _20811_);
  and _53719_ (_21300_, _21270_, _21299_);
  or _53720_ (_21301_, _21300_, _21298_);
  or _53721_ (_21302_, _21301_, _21296_);
  or _53722_ (_21303_, _21302_, _21295_);
  and _53723_ (_21304_, _21303_, _20941_);
  or _53724_ (_21305_, _21304_, _21292_);
  and _53725_ (_21306_, _21305_, _20985_);
  and _53726_ (_21307_, _21285_, _20940_);
  nand _53727_ (_21308_, _20985_, _20767_);
  nand _53728_ (_21309_, _21308_, _20810_);
  and _53729_ (_21310_, _21309_, _21307_);
  or _53730_ (_21311_, _21310_, _21306_);
  or _53731_ (_21312_, _21311_, _21289_);
  nor _53732_ (_21313_, _19868_, _22789_);
  nor _53733_ (_21314_, _19982_, _22767_);
  and _53734_ (_21315_, _19982_, _22767_);
  or _53735_ (_21316_, _21315_, _21314_);
  nor _53736_ (_21317_, _19889_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _53737_ (_21318_, _19889_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or _53738_ (_21319_, _21318_, _21317_);
  or _53739_ (_21320_, _21319_, _21316_);
  or _53740_ (_21321_, _21320_, _21313_);
  or _53741_ (_21322_, _19882_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _53742_ (_21323_, _19882_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _53743_ (_21324_, _21323_, _21322_);
  and _53744_ (_21325_, _19868_, _22789_);
  or _53745_ (_21326_, _21325_, _21324_);
  or _53746_ (_21327_, _21326_, _21321_);
  or _53747_ (_21328_, _19878_, _26128_);
  nand _53748_ (_21329_, _19878_, _26128_);
  and _53749_ (_21330_, _21329_, _21328_);
  nor _53750_ (_21331_, _19938_, _22772_);
  and _53751_ (_21332_, _20028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _53752_ (_21333_, _20028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53753_ (_21334_, _21333_, _21332_);
  nor _53754_ (_21335_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _53755_ (_21336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _53756_ (_21337_, _21336_, _21335_);
  nand _53757_ (_21338_, _21337_, _20307_);
  nor _53758_ (_21339_, _20112_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53759_ (_21340_, _20112_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _53760_ (_21341_, _21340_, _21339_);
  or _53761_ (_21342_, _21341_, _21338_);
  or _53762_ (_21343_, _21342_, _21334_);
  nor _53763_ (_21344_, _20024_, _22762_);
  and _53764_ (_21345_, _20024_, _22762_);
  or _53765_ (_21346_, _21345_, _21344_);
  or _53766_ (_21347_, _21346_, _21343_);
  and _53767_ (_21348_, _19938_, _22772_);
  or _53768_ (_21349_, _21348_, _21347_);
  or _53769_ (_21350_, _21349_, _21331_);
  or _53770_ (_21351_, _21350_, _21221_);
  or _53771_ (_21352_, _21351_, _21330_);
  or _53772_ (_21353_, _21352_, _21327_);
  or _53773_ (_21354_, _21353_, _21240_);
  and _53774_ (_21355_, _21354_, _21312_);
  and _53775_ (_21356_, _20898_, _20723_);
  and _53776_ (_21357_, _21356_, _21294_);
  and _53777_ (_21358_, _21286_, _21297_);
  or _53778_ (_21359_, _21358_, _21357_);
  and _53779_ (_21360_, _21359_, _20986_);
  not _53780_ (_21361_, _21276_);
  or _53781_ (_21362_, _21307_, _21361_);
  and _53782_ (_21363_, _20722_, _20678_);
  and _53783_ (_21364_, _21363_, _20898_);
  and _53784_ (_21365_, _21364_, _20940_);
  or _53785_ (_21366_, _21365_, _21276_);
  and _53786_ (_21367_, _21366_, _21269_);
  and _53787_ (_21368_, _21367_, _21362_);
  or _53788_ (_21369_, _21368_, _21360_);
  and _53789_ (_21370_, _20518_, _19838_);
  and _53790_ (_21371_, _21370_, _19842_);
  and _53791_ (_21372_, _21371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _53792_ (_21373_, _21372_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _53793_ (_21374_, _21373_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _53794_ (_21375_, _21373_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _53795_ (_21376_, _21375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _53796_ (_21377_, _21376_, _20240_);
  nor _53797_ (_21378_, _21377_, _21374_);
  and _53798_ (_21379_, _21374_, _20241_);
  and _53799_ (_21380_, _20518_, _19837_);
  nor _53800_ (_21381_, _21380_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _53801_ (_21382_, _21381_, _21370_);
  and _53802_ (_21383_, _21382_, _26136_);
  nor _53803_ (_21384_, _21382_, _26136_);
  or _53804_ (_21385_, _21384_, _21383_);
  and _53805_ (_21386_, _20518_, _19836_);
  nor _53806_ (_21387_, _21386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _53807_ (_21389_, _21387_, _21380_);
  nor _53808_ (_21390_, _21389_, _22772_);
  and _53809_ (_21391_, _21370_, _19840_);
  and _53810_ (_21392_, _21370_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _53811_ (_21393_, _21392_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _53812_ (_21394_, _21393_, _21391_);
  nor _53813_ (_21395_, _21394_, _26128_);
  and _53814_ (_21396_, _21389_, _22772_);
  or _53815_ (_21397_, _21396_, _21395_);
  or _53816_ (_21398_, _21397_, _21390_);
  and _53817_ (_21399_, _20518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _53818_ (_21400_, _20518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _53819_ (_21401_, _21400_, _21399_);
  nand _53820_ (_21402_, _21401_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _53821_ (_21403_, _21401_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _53822_ (_21404_, _21403_, _21402_);
  nor _53823_ (_21405_, _21370_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _53824_ (_21406_, _21405_, _21392_);
  and _53825_ (_21407_, _21406_, _22780_);
  or _53826_ (_21408_, _21407_, _21404_);
  nor _53827_ (_21409_, _21399_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _53828_ (_21410_, _21409_, _21386_);
  and _53829_ (_21411_, _21410_, _22767_);
  nor _53830_ (_21412_, _21410_, _22767_);
  or _53831_ (_21413_, _21412_, _21411_);
  or _53832_ (_21414_, _21413_, _21408_);
  and _53833_ (_21415_, _21394_, _26128_);
  nor _53834_ (_21416_, _21406_, _22780_);
  or _53835_ (_21417_, _20520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _53836_ (_21418_, _20520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53837_ (_21419_, _21418_, _21417_);
  nor _53838_ (_21420_, _19756_, _19781_);
  nor _53839_ (_21421_, _21420_, _09640_);
  and _53840_ (_21422_, _21420_, _09640_);
  nor _53841_ (_21423_, _21422_, _21421_);
  nand _53842_ (_21424_, _21423_, _20308_);
  nor _53843_ (_21425_, _20523_, _26153_);
  and _53844_ (_21426_, _20523_, _26153_);
  or _53845_ (_21427_, _21426_, _21425_);
  or _53846_ (_21428_, _21427_, _21424_);
  or _53847_ (_21429_, _21428_, _21419_);
  or _53848_ (_21430_, _21429_, _21416_);
  or _53849_ (_21431_, _21430_, _21415_);
  or _53850_ (_21432_, _21431_, _21414_);
  or _53851_ (_21433_, _21432_, _21398_);
  or _53852_ (_21434_, _21433_, _21385_);
  or _53853_ (_21435_, _21434_, _21379_);
  nor _53854_ (_21436_, _21372_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _53855_ (_21437_, _21436_, _21373_);
  nor _53856_ (_21438_, _21437_, _26114_);
  and _53857_ (_21439_, _21437_, _26114_);
  or _53858_ (_21440_, _21439_, _21438_);
  or _53859_ (_21441_, _21440_, _21435_);
  or _53860_ (_21442_, _21375_, _21374_);
  and _53861_ (_21443_, _21442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _53862_ (_21444_, _21371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _53863_ (_21445_, _21444_, _21372_);
  nor _53864_ (_21446_, _21445_, _22797_);
  and _53865_ (_21447_, _21445_, _22797_);
  and _53866_ (_21448_, _21370_, _19841_);
  or _53867_ (_21449_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nand _53868_ (_21450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _53869_ (_21451_, _21450_, _21449_);
  or _53870_ (_21452_, _21451_, _21448_);
  nand _53871_ (_21453_, _21451_, _21448_);
  and _53872_ (_21454_, _21453_, _21452_);
  nor _53873_ (_21455_, _21391_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _53874_ (_21456_, _21455_, _21448_);
  nor _53875_ (_21457_, _21456_, _22789_);
  and _53876_ (_21458_, _21456_, _22789_);
  or _53877_ (_21459_, _21458_, _21457_);
  or _53878_ (_21460_, _21459_, _21454_);
  or _53879_ (_21461_, _21460_, _21447_);
  or _53880_ (_21462_, _21461_, _21446_);
  or _53881_ (_21463_, _21462_, _21443_);
  or _53882_ (_21464_, _21463_, _21441_);
  or _53883_ (_21465_, _21464_, _21378_);
  and _53884_ (_21466_, _21465_, _21369_);
  nor _53885_ (_21467_, _20897_, _20767_);
  and _53886_ (_21468_, _21467_, _21271_);
  not _53887_ (_21469_, _20984_);
  or _53888_ (_21470_, _21294_, _21469_);
  and _53889_ (_21471_, _20941_, _20897_);
  and _53890_ (_21472_, _21471_, _21470_);
  or _53891_ (_21473_, _21472_, _21468_);
  and _53892_ (_21474_, _21469_, _20897_);
  not _53893_ (_21475_, _20721_);
  and _53894_ (_21476_, _20855_, _21475_);
  and _53895_ (_21477_, _21476_, _21199_);
  or _53896_ (_21478_, _21477_, _21474_);
  and _53897_ (_21479_, _21478_, _21293_);
  and _53898_ (_21480_, _21298_, _20940_);
  or _53899_ (_21481_, _20896_, _21475_);
  nand _53900_ (_21482_, _20984_, _20678_);
  nor _53901_ (_21483_, _21482_, _21481_);
  or _53902_ (_21484_, _21483_, _21300_);
  and _53903_ (_21485_, _21484_, _20940_);
  or _53904_ (_21486_, _21485_, _21480_);
  or _53905_ (_21487_, _21486_, _21479_);
  or _53906_ (_21488_, _21487_, _21473_);
  and _53907_ (_21489_, _21284_, _21299_);
  or _53908_ (_21490_, _21274_, _20767_);
  and _53909_ (_21491_, _21481_, _20940_);
  and _53910_ (_21492_, _21491_, _21490_);
  or _53911_ (_21493_, _21492_, _21489_);
  and _53912_ (_21494_, _21493_, _20985_);
  and _53913_ (_21495_, _21275_, _20812_);
  or _53914_ (_21496_, _21495_, _21364_);
  or _53915_ (_21497_, _21270_, _20813_);
  and _53916_ (_21498_, _21497_, _21269_);
  or _53917_ (_21499_, _21498_, _21496_);
  and _53918_ (_21500_, _21499_, _20941_);
  or _53919_ (_21501_, _21500_, _21494_);
  or _53920_ (_21502_, _21501_, _21488_);
  and _53921_ (_21503_, _19852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53922_ (_21504_, _21503_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _53923_ (_21505_, _21504_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _53924_ (_21506_, _21505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _53925_ (_21507_, _21505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _53926_ (_21508_, _21507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _53927_ (_21509_, _21508_, _20240_);
  nor _53928_ (_21510_, _21509_, _21506_);
  nand _53929_ (_21511_, _20240_, _22806_);
  and _53930_ (_21512_, _21511_, _21506_);
  and _53931_ (_21513_, _19838_, _19743_);
  and _53932_ (_21514_, _21513_, _19842_);
  and _53933_ (_21515_, _21514_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _53934_ (_21516_, _21515_, _22802_);
  and _53935_ (_21517_, _21515_, _22802_);
  nor _53936_ (_21518_, _21517_, _21516_);
  and _53937_ (_21520_, _21518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _53938_ (_21521_, _21507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or _53939_ (_21522_, _21521_, _21520_);
  or _53940_ (_21523_, _21522_, _21512_);
  nor _53941_ (_21524_, _21503_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _53942_ (_21525_, _21524_, _21504_);
  and _53943_ (_21526_, _21525_, _22797_);
  nor _53944_ (_21527_, _21525_, _22797_);
  and _53945_ (_21528_, _21513_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _53946_ (_21529_, _21513_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _53947_ (_21530_, _21529_, _21528_);
  nand _53948_ (_21531_, _21530_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or _53949_ (_21532_, _21530_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _53950_ (_21533_, _21532_, _21531_);
  and _53951_ (_21534_, _19886_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53952_ (_21535_, _19836_, _19743_);
  nor _53953_ (_21536_, _21535_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _53954_ (_21537_, _21536_, _21534_);
  nor _53955_ (_21538_, _21537_, _22772_);
  and _53956_ (_21539_, _21537_, _22772_);
  or _53957_ (_21540_, _21539_, _21538_);
  and _53958_ (_21541_, _19743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _53959_ (_21542_, _19743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _53960_ (_21543_, _21542_, _21541_);
  nand _53961_ (_21544_, _21543_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _53962_ (_21545_, _21543_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _53963_ (_21546_, _21545_, _21544_);
  or _53964_ (_21547_, _19745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _53965_ (_21548_, _19745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53966_ (_21549_, _21548_, _21547_);
  or _53967_ (_21550_, _21549_, _21546_);
  or _53968_ (_21551_, _21550_, _21540_);
  or _53969_ (_21552_, _21551_, _21533_);
  and _53970_ (_21553_, _21513_, _19841_);
  and _53971_ (_21554_, _21513_, _19840_);
  nor _53972_ (_21555_, _21554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _53973_ (_21556_, _21555_, _21553_);
  nor _53974_ (_21557_, _21556_, _22789_);
  and _53975_ (_21558_, _21556_, _22789_);
  or _53976_ (_21559_, _21558_, _21557_);
  or _53977_ (_21560_, _21559_, _21552_);
  or _53978_ (_21561_, _21560_, _21527_);
  or _53979_ (_21562_, _21561_, _21526_);
  nor _53980_ (_21563_, _21518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _53981_ (_21564_, _21528_, _22784_);
  and _53982_ (_21565_, _21528_, _22784_);
  nor _53983_ (_21566_, _21565_, _21564_);
  nor _53984_ (_21567_, _21566_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _53985_ (_21568_, _21566_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _53986_ (_21569_, _21534_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _53987_ (_21570_, _21569_, _21513_);
  nor _53988_ (_21571_, _21570_, _26136_);
  or _53989_ (_21572_, _19741_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _53990_ (_21573_, _19741_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53991_ (_21574_, _21573_, _21572_);
  nor _53992_ (_21575_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _53993_ (_21576_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or _53994_ (_21577_, _21576_, _21575_);
  and _53995_ (_21578_, _21577_, _21541_);
  nor _53996_ (_21579_, _21577_, _21541_);
  or _53997_ (_21580_, _21579_, _21578_);
  or _53998_ (_21581_, _21423_, _20307_);
  or _53999_ (_21582_, _21581_, _21580_);
  or _54000_ (_21583_, _21582_, _21574_);
  or _54001_ (_21584_, _21583_, _21571_);
  and _54002_ (_21585_, _21570_, _26136_);
  or _54003_ (_21586_, _21553_, _21451_);
  nand _54004_ (_21587_, _21553_, _21451_);
  and _54005_ (_21588_, _21587_, _21586_);
  or _54006_ (_21589_, _21588_, _21585_);
  or _54007_ (_21590_, _21589_, _21584_);
  or _54008_ (_21591_, _21590_, _21568_);
  or _54009_ (_21592_, _21591_, _21567_);
  or _54010_ (_21593_, _21592_, _21563_);
  or _54011_ (_21594_, _21593_, _21562_);
  or _54012_ (_21595_, _21594_, _21523_);
  or _54013_ (_21596_, _21595_, _21510_);
  and _54014_ (_21597_, _21596_, _21502_);
  or _54015_ (_21598_, _21597_, _21466_);
  or _54016_ (_21599_, _21598_, _21355_);
  or _54017_ (_21600_, _21599_, _21268_);
  and _54018_ (_21601_, _21600_, _20636_);
  or _54019_ (_21602_, _21601_, _21207_);
  or _54020_ (property_invalid, _21602_, _20990_);
  and _54021_ (_21603_, _24017_, _23548_);
  and _54022_ (_21604_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or _54023_ (_12202_, _21604_, _21603_);
  and _54024_ (_21605_, _20630_, first_instr);
  or _54025_ (_00000_, _21605_, rst);
  and _54026_ (_21606_, _16026_, _24051_);
  and _54027_ (_21607_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or _54028_ (_12224_, _21607_, _21606_);
  and _54029_ (_21608_, _03033_, _23996_);
  and _54030_ (_21609_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or _54031_ (_12251_, _21609_, _21608_);
  and _54032_ (_21610_, _16008_, _23996_);
  and _54033_ (_21611_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or _54034_ (_12261_, _21611_, _21610_);
  and _54035_ (_21612_, _03033_, _24134_);
  and _54036_ (_21613_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or _54037_ (_12268_, _21613_, _21612_);
  and _54038_ (_21614_, _05442_, _23583_);
  and _54039_ (_21615_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _54040_ (_12274_, _21615_, _21614_);
  and _54041_ (_21616_, _05438_, _23996_);
  and _54042_ (_21617_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _54043_ (_12280_, _21617_, _21616_);
  and _54044_ (_21618_, _05438_, _23583_);
  and _54045_ (_21619_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _54046_ (_12293_, _21619_, _21618_);
  and _54047_ (_21621_, _02964_, _24051_);
  and _54048_ (_21622_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _54049_ (_27186_, _21622_, _21621_);
  and _54050_ (_21623_, _03355_, _23996_);
  and _54051_ (_21624_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _54052_ (_12301_, _21624_, _21623_);
  or _54053_ (_21625_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _54054_ (_21626_, _21625_, _22731_);
  nand _54055_ (_21627_, _24189_, _23542_);
  and _54056_ (_12316_, _21627_, _21626_);
  nand _54057_ (_21628_, _24210_, _24184_);
  or _54058_ (_21629_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _54059_ (_21630_, _21629_, _22731_);
  and _54060_ (_12325_, _21630_, _21628_);
  and _54061_ (_21631_, _05442_, _24134_);
  and _54062_ (_21632_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _54063_ (_12332_, _21632_, _21631_);
  and _54064_ (_21633_, _03287_, _24219_);
  and _54065_ (_21634_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or _54066_ (_12334_, _21634_, _21633_);
  and _54067_ (_21635_, _03287_, _23548_);
  and _54068_ (_21636_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or _54069_ (_12340_, _21636_, _21635_);
  and _54070_ (_21637_, _05485_, _23583_);
  and _54071_ (_21638_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _54072_ (_12342_, _21638_, _21637_);
  and _54073_ (_21639_, _16026_, _23548_);
  and _54074_ (_21640_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or _54075_ (_12344_, _21640_, _21639_);
  and _54076_ (_21641_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _54077_ (_21643_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _54078_ (_21644_, _21643_, _21641_);
  and _54079_ (_21645_, _21644_, _09792_);
  and _54080_ (_21646_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and _54081_ (_21647_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _54082_ (_21648_, _21647_, _21646_);
  and _54083_ (_21649_, _21648_, _05549_);
  or _54084_ (_21650_, _21649_, _21645_);
  or _54085_ (_21651_, _21650_, _09791_);
  and _54086_ (_21652_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and _54087_ (_21653_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _54088_ (_21654_, _21653_, _21652_);
  and _54089_ (_21655_, _21654_, _09792_);
  and _54090_ (_21656_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and _54091_ (_21657_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _54092_ (_21658_, _21657_, _21656_);
  and _54093_ (_21659_, _21658_, _05549_);
  or _54094_ (_21660_, _21659_, _21655_);
  or _54095_ (_21661_, _21660_, _05535_);
  and _54096_ (_21662_, _21661_, _09805_);
  and _54097_ (_21663_, _21662_, _21651_);
  or _54098_ (_21664_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _54099_ (_21665_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and _54100_ (_21666_, _21665_, _21664_);
  and _54101_ (_21667_, _21666_, _09792_);
  or _54102_ (_21668_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _54103_ (_21669_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and _54104_ (_21670_, _21669_, _21668_);
  and _54105_ (_21671_, _21670_, _05549_);
  or _54106_ (_21672_, _21671_, _21667_);
  or _54107_ (_21673_, _21672_, _09791_);
  or _54108_ (_21674_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _54109_ (_21675_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and _54110_ (_21676_, _21675_, _21674_);
  and _54111_ (_21677_, _21676_, _09792_);
  or _54112_ (_21678_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _54113_ (_21679_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and _54114_ (_21680_, _21679_, _21678_);
  and _54115_ (_21681_, _21680_, _05549_);
  or _54116_ (_21682_, _21681_, _21677_);
  or _54117_ (_21683_, _21682_, _05535_);
  and _54118_ (_21684_, _21683_, _05542_);
  and _54119_ (_21685_, _21684_, _21673_);
  or _54120_ (_21686_, _21685_, _21663_);
  and _54121_ (_21687_, _21686_, _05518_);
  and _54122_ (_21688_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and _54123_ (_21689_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _54124_ (_21690_, _21689_, _21688_);
  and _54125_ (_21691_, _21690_, _09792_);
  and _54126_ (_21692_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and _54127_ (_21693_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _54128_ (_21694_, _21693_, _21692_);
  and _54129_ (_21695_, _21694_, _05549_);
  or _54130_ (_21696_, _21695_, _21691_);
  or _54131_ (_21697_, _21696_, _09791_);
  and _54132_ (_21698_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and _54133_ (_21699_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _54134_ (_21700_, _21699_, _21698_);
  and _54135_ (_21701_, _21700_, _09792_);
  and _54136_ (_21702_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and _54137_ (_21703_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _54138_ (_21704_, _21703_, _21702_);
  and _54139_ (_21705_, _21704_, _05549_);
  or _54140_ (_21706_, _21705_, _21701_);
  or _54141_ (_21707_, _21706_, _05535_);
  and _54142_ (_21708_, _21707_, _09805_);
  and _54143_ (_21709_, _21708_, _21697_);
  or _54144_ (_21710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _54145_ (_21711_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and _54146_ (_21712_, _21711_, _05549_);
  and _54147_ (_21713_, _21712_, _21710_);
  or _54148_ (_21714_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _54149_ (_21715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and _54150_ (_21716_, _21715_, _09792_);
  and _54151_ (_21717_, _21716_, _21714_);
  or _54152_ (_21718_, _21717_, _21713_);
  or _54153_ (_21719_, _21718_, _09791_);
  or _54154_ (_21720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _54155_ (_21721_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and _54156_ (_21722_, _21721_, _05549_);
  and _54157_ (_21723_, _21722_, _21720_);
  or _54158_ (_21724_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _54159_ (_21725_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and _54160_ (_21726_, _21725_, _09792_);
  and _54161_ (_21727_, _21726_, _21724_);
  or _54162_ (_21728_, _21727_, _21723_);
  or _54163_ (_21729_, _21728_, _05535_);
  and _54164_ (_21730_, _21729_, _05542_);
  and _54165_ (_21731_, _21730_, _21719_);
  or _54166_ (_21732_, _21731_, _21709_);
  and _54167_ (_21733_, _21732_, _09850_);
  or _54168_ (_21734_, _21733_, _21687_);
  and _54169_ (_21735_, _21734_, _09790_);
  and _54170_ (_21736_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and _54171_ (_21737_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _54172_ (_21738_, _21737_, _21736_);
  and _54173_ (_21739_, _21738_, _09792_);
  and _54174_ (_21740_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and _54175_ (_21741_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _54176_ (_21742_, _21741_, _21740_);
  and _54177_ (_21743_, _21742_, _05549_);
  or _54178_ (_21744_, _21743_, _21739_);
  and _54179_ (_21745_, _21744_, _05535_);
  and _54180_ (_21746_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _54181_ (_21747_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _54182_ (_21748_, _21747_, _21746_);
  and _54183_ (_21749_, _21748_, _09792_);
  and _54184_ (_21750_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and _54185_ (_21751_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _54186_ (_21752_, _21751_, _21750_);
  and _54187_ (_21753_, _21752_, _05549_);
  or _54188_ (_21754_, _21753_, _21749_);
  and _54189_ (_21755_, _21754_, _09791_);
  or _54190_ (_21756_, _21755_, _21745_);
  and _54191_ (_21757_, _21756_, _09805_);
  or _54192_ (_21758_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _54193_ (_21759_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _54194_ (_21760_, _21759_, _05549_);
  and _54195_ (_21761_, _21760_, _21758_);
  or _54196_ (_21762_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _54197_ (_21763_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _54198_ (_21764_, _21763_, _09792_);
  and _54199_ (_21765_, _21764_, _21762_);
  or _54200_ (_21766_, _21765_, _21761_);
  and _54201_ (_21767_, _21766_, _05535_);
  or _54202_ (_21768_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _54203_ (_21769_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _54204_ (_21770_, _21769_, _05549_);
  and _54205_ (_21771_, _21770_, _21768_);
  or _54206_ (_21772_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _54207_ (_21773_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _54208_ (_21774_, _21773_, _09792_);
  and _54209_ (_21775_, _21774_, _21772_);
  or _54210_ (_21776_, _21775_, _21771_);
  and _54211_ (_21777_, _21776_, _09791_);
  or _54212_ (_21778_, _21777_, _21767_);
  and _54213_ (_21779_, _21778_, _05542_);
  or _54214_ (_21780_, _21779_, _21757_);
  and _54215_ (_21781_, _21780_, _09850_);
  and _54216_ (_21782_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and _54217_ (_21783_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _54218_ (_21784_, _21783_, _21782_);
  and _54219_ (_21785_, _21784_, _09792_);
  and _54220_ (_21786_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and _54221_ (_21787_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _54222_ (_21788_, _21787_, _21786_);
  and _54223_ (_21789_, _21788_, _05549_);
  or _54224_ (_21790_, _21789_, _21785_);
  and _54225_ (_21791_, _21790_, _05535_);
  and _54226_ (_21792_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and _54227_ (_21793_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _54228_ (_21794_, _21793_, _21792_);
  and _54229_ (_21795_, _21794_, _09792_);
  and _54230_ (_21796_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and _54231_ (_21797_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _54232_ (_21798_, _21797_, _21796_);
  and _54233_ (_21799_, _21798_, _05549_);
  or _54234_ (_21800_, _21799_, _21795_);
  and _54235_ (_21801_, _21800_, _09791_);
  or _54236_ (_21802_, _21801_, _21791_);
  and _54237_ (_21803_, _21802_, _09805_);
  or _54238_ (_21804_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _54239_ (_21805_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and _54240_ (_21806_, _21805_, _21804_);
  and _54241_ (_21807_, _21806_, _09792_);
  or _54242_ (_21808_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _54243_ (_21809_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and _54244_ (_21810_, _21809_, _21808_);
  and _54245_ (_21811_, _21810_, _05549_);
  or _54246_ (_21812_, _21811_, _21807_);
  and _54247_ (_21813_, _21812_, _05535_);
  or _54248_ (_21814_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _54249_ (_21815_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and _54250_ (_21816_, _21815_, _21814_);
  and _54251_ (_21817_, _21816_, _09792_);
  or _54252_ (_21818_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _54253_ (_21819_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and _54254_ (_21820_, _21819_, _21818_);
  and _54255_ (_21821_, _21820_, _05549_);
  or _54256_ (_21822_, _21821_, _21817_);
  and _54257_ (_21823_, _21822_, _09791_);
  or _54258_ (_21824_, _21823_, _21813_);
  and _54259_ (_21825_, _21824_, _05542_);
  or _54260_ (_21826_, _21825_, _21803_);
  and _54261_ (_21827_, _21826_, _05518_);
  or _54262_ (_21828_, _21827_, _21781_);
  and _54263_ (_21829_, _21828_, _05520_);
  or _54264_ (_21830_, _21829_, _21735_);
  or _54265_ (_21831_, _21830_, _05526_);
  and _54266_ (_21832_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and _54267_ (_21833_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _54268_ (_21834_, _21833_, _21832_);
  and _54269_ (_21835_, _21834_, _09792_);
  and _54270_ (_21836_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and _54271_ (_21837_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _54272_ (_21838_, _21837_, _21836_);
  and _54273_ (_21839_, _21838_, _05549_);
  or _54274_ (_21840_, _21839_, _21835_);
  or _54275_ (_21841_, _21840_, _09791_);
  and _54276_ (_21842_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and _54277_ (_21843_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _54278_ (_21844_, _21843_, _21842_);
  and _54279_ (_21845_, _21844_, _09792_);
  and _54280_ (_21846_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and _54281_ (_21847_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _54282_ (_21848_, _21847_, _21846_);
  and _54283_ (_21849_, _21848_, _05549_);
  or _54284_ (_21850_, _21849_, _21845_);
  or _54285_ (_21851_, _21850_, _05535_);
  and _54286_ (_21852_, _21851_, _09805_);
  and _54287_ (_21853_, _21852_, _21841_);
  or _54288_ (_21854_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _54289_ (_21855_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and _54290_ (_21856_, _21855_, _05549_);
  and _54291_ (_21857_, _21856_, _21854_);
  or _54292_ (_21858_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _54293_ (_21859_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and _54294_ (_21860_, _21859_, _09792_);
  and _54295_ (_21861_, _21860_, _21858_);
  or _54296_ (_21862_, _21861_, _21857_);
  or _54297_ (_21863_, _21862_, _09791_);
  or _54298_ (_21864_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _54299_ (_21865_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and _54300_ (_21866_, _21865_, _05549_);
  and _54301_ (_21867_, _21866_, _21864_);
  or _54302_ (_21868_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _54303_ (_21869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and _54304_ (_21870_, _21869_, _09792_);
  and _54305_ (_21871_, _21870_, _21868_);
  or _54306_ (_21872_, _21871_, _21867_);
  or _54307_ (_21873_, _21872_, _05535_);
  and _54308_ (_21874_, _21873_, _05542_);
  and _54309_ (_21875_, _21874_, _21863_);
  or _54310_ (_21876_, _21875_, _21853_);
  and _54311_ (_21877_, _21876_, _09850_);
  and _54312_ (_21878_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and _54313_ (_21879_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _54314_ (_21880_, _21879_, _21878_);
  and _54315_ (_21881_, _21880_, _09792_);
  and _54316_ (_21882_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and _54317_ (_21883_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _54318_ (_21884_, _21883_, _21882_);
  and _54319_ (_21885_, _21884_, _05549_);
  or _54320_ (_21886_, _21885_, _21881_);
  or _54321_ (_21887_, _21886_, _09791_);
  and _54322_ (_21888_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and _54323_ (_21889_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _54324_ (_21890_, _21889_, _21888_);
  and _54325_ (_21891_, _21890_, _09792_);
  and _54326_ (_21892_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and _54327_ (_21893_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _54328_ (_21894_, _21893_, _21892_);
  and _54329_ (_21895_, _21894_, _05549_);
  or _54330_ (_21896_, _21895_, _21891_);
  or _54331_ (_21897_, _21896_, _05535_);
  and _54332_ (_21898_, _21897_, _09805_);
  and _54333_ (_21899_, _21898_, _21887_);
  or _54334_ (_21900_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _54335_ (_21901_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and _54336_ (_21902_, _21901_, _21900_);
  and _54337_ (_21903_, _21902_, _09792_);
  or _54338_ (_21904_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _54339_ (_21905_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _54340_ (_21906_, _21905_, _21904_);
  and _54341_ (_21907_, _21906_, _05549_);
  or _54342_ (_21908_, _21907_, _21903_);
  or _54343_ (_21909_, _21908_, _09791_);
  or _54344_ (_21910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _54345_ (_21911_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and _54346_ (_21912_, _21911_, _21910_);
  and _54347_ (_21913_, _21912_, _09792_);
  or _54348_ (_21914_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _54349_ (_21915_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and _54350_ (_21916_, _21915_, _21914_);
  and _54351_ (_21917_, _21916_, _05549_);
  or _54352_ (_21918_, _21917_, _21913_);
  or _54353_ (_21919_, _21918_, _05535_);
  and _54354_ (_21920_, _21919_, _05542_);
  and _54355_ (_21921_, _21920_, _21909_);
  or _54356_ (_21922_, _21921_, _21899_);
  and _54357_ (_21923_, _21922_, _05518_);
  or _54358_ (_21924_, _21923_, _21877_);
  and _54359_ (_21925_, _21924_, _09790_);
  or _54360_ (_21926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _54361_ (_21927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and _54362_ (_21928_, _21927_, _21926_);
  and _54363_ (_21929_, _21928_, _09792_);
  or _54364_ (_21930_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _54365_ (_21931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and _54366_ (_21932_, _21931_, _21930_);
  and _54367_ (_21933_, _21932_, _05549_);
  or _54368_ (_21934_, _21933_, _21929_);
  and _54369_ (_21935_, _21934_, _09791_);
  or _54370_ (_21936_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _54371_ (_21937_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and _54372_ (_21938_, _21937_, _21936_);
  and _54373_ (_21939_, _21938_, _09792_);
  or _54374_ (_21940_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _54375_ (_21941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and _54376_ (_21942_, _21941_, _21940_);
  and _54377_ (_21943_, _21942_, _05549_);
  or _54378_ (_21944_, _21943_, _21939_);
  and _54379_ (_21945_, _21944_, _05535_);
  or _54380_ (_21946_, _21945_, _21935_);
  and _54381_ (_21947_, _21946_, _05542_);
  and _54382_ (_21948_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and _54383_ (_21949_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _54384_ (_21950_, _21949_, _21948_);
  and _54385_ (_21951_, _21950_, _09792_);
  and _54386_ (_21952_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and _54387_ (_21953_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _54388_ (_21954_, _21953_, _21952_);
  and _54389_ (_21955_, _21954_, _05549_);
  or _54390_ (_21956_, _21955_, _21951_);
  and _54391_ (_21957_, _21956_, _09791_);
  and _54392_ (_21958_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and _54393_ (_21959_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _54394_ (_21960_, _21959_, _21958_);
  and _54395_ (_21961_, _21960_, _09792_);
  and _54396_ (_21962_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and _54397_ (_21963_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _54398_ (_21964_, _21963_, _21962_);
  and _54399_ (_21965_, _21964_, _05549_);
  or _54400_ (_21966_, _21965_, _21961_);
  and _54401_ (_21967_, _21966_, _05535_);
  or _54402_ (_21968_, _21967_, _21957_);
  and _54403_ (_21969_, _21968_, _09805_);
  or _54404_ (_21970_, _21969_, _21947_);
  and _54405_ (_21971_, _21970_, _05518_);
  or _54406_ (_21972_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _54407_ (_21973_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and _54408_ (_21974_, _21973_, _05549_);
  and _54409_ (_21975_, _21974_, _21972_);
  or _54410_ (_21976_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or _54411_ (_21977_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and _54412_ (_21978_, _21977_, _09792_);
  and _54413_ (_21979_, _21978_, _21976_);
  or _54414_ (_21980_, _21979_, _21975_);
  and _54415_ (_21981_, _21980_, _09791_);
  or _54416_ (_21982_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _54417_ (_21983_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and _54418_ (_21984_, _21983_, _05549_);
  and _54419_ (_21985_, _21984_, _21982_);
  or _54420_ (_21986_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or _54421_ (_21987_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and _54422_ (_21988_, _21987_, _09792_);
  and _54423_ (_21989_, _21988_, _21986_);
  or _54424_ (_21990_, _21989_, _21985_);
  and _54425_ (_21991_, _21990_, _05535_);
  or _54426_ (_21992_, _21991_, _21981_);
  and _54427_ (_21993_, _21992_, _05542_);
  and _54428_ (_21994_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and _54429_ (_21995_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _54430_ (_21996_, _21995_, _21994_);
  and _54431_ (_21997_, _21996_, _09792_);
  and _54432_ (_21998_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and _54433_ (_21999_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _54434_ (_22000_, _21999_, _21998_);
  and _54435_ (_22001_, _22000_, _05549_);
  or _54436_ (_22002_, _22001_, _21997_);
  and _54437_ (_22003_, _22002_, _09791_);
  and _54438_ (_22004_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and _54439_ (_22005_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or _54440_ (_22006_, _22005_, _22004_);
  and _54441_ (_22007_, _22006_, _09792_);
  and _54442_ (_22008_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and _54443_ (_22009_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _54444_ (_22010_, _22009_, _22008_);
  and _54445_ (_22011_, _22010_, _05549_);
  or _54446_ (_22012_, _22011_, _22007_);
  and _54447_ (_22013_, _22012_, _05535_);
  or _54448_ (_22014_, _22013_, _22003_);
  and _54449_ (_22015_, _22014_, _09805_);
  or _54450_ (_22016_, _22015_, _21993_);
  and _54451_ (_22017_, _22016_, _09850_);
  or _54452_ (_22018_, _22017_, _21971_);
  and _54453_ (_22019_, _22018_, _05520_);
  or _54454_ (_22020_, _22019_, _21925_);
  or _54455_ (_22021_, _22020_, _10033_);
  and _54456_ (_22022_, _22021_, _21831_);
  or _54457_ (_22023_, _22022_, _00143_);
  and _54458_ (_22024_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and _54459_ (_22025_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _54460_ (_22026_, _22025_, _22024_);
  and _54461_ (_22027_, _22026_, _09792_);
  and _54462_ (_22028_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and _54463_ (_22029_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _54464_ (_22030_, _22029_, _22028_);
  and _54465_ (_22031_, _22030_, _05549_);
  or _54466_ (_22032_, _22031_, _22027_);
  or _54467_ (_22033_, _22032_, _09791_);
  and _54468_ (_22034_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and _54469_ (_22035_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _54470_ (_22036_, _22035_, _22034_);
  and _54471_ (_22037_, _22036_, _09792_);
  and _54472_ (_22038_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and _54473_ (_22039_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _54474_ (_22040_, _22039_, _22038_);
  and _54475_ (_22041_, _22040_, _05549_);
  or _54476_ (_22042_, _22041_, _22037_);
  or _54477_ (_22043_, _22042_, _05535_);
  and _54478_ (_22044_, _22043_, _09805_);
  and _54479_ (_22045_, _22044_, _22033_);
  or _54480_ (_22046_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _54481_ (_22047_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and _54482_ (_22048_, _22047_, _22046_);
  and _54483_ (_22049_, _22048_, _09792_);
  or _54484_ (_22050_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _54485_ (_22051_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and _54486_ (_22052_, _22051_, _22050_);
  and _54487_ (_22053_, _22052_, _05549_);
  or _54488_ (_22054_, _22053_, _22049_);
  or _54489_ (_22055_, _22054_, _09791_);
  or _54490_ (_22056_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _54491_ (_22057_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and _54492_ (_22058_, _22057_, _22056_);
  and _54493_ (_22059_, _22058_, _09792_);
  or _54494_ (_22060_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _54495_ (_22061_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and _54496_ (_22062_, _22061_, _22060_);
  and _54497_ (_22063_, _22062_, _05549_);
  or _54498_ (_22064_, _22063_, _22059_);
  or _54499_ (_22065_, _22064_, _05535_);
  and _54500_ (_22066_, _22065_, _05542_);
  and _54501_ (_22067_, _22066_, _22055_);
  or _54502_ (_22068_, _22067_, _22045_);
  and _54503_ (_22069_, _22068_, _05518_);
  and _54504_ (_22070_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _54505_ (_22071_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _54506_ (_22072_, _22071_, _22070_);
  and _54507_ (_22073_, _22072_, _09792_);
  and _54508_ (_22074_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _54509_ (_22075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _54510_ (_22076_, _22075_, _22074_);
  and _54511_ (_22077_, _22076_, _05549_);
  or _54512_ (_22078_, _22077_, _22073_);
  or _54513_ (_22079_, _22078_, _09791_);
  and _54514_ (_22080_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _54515_ (_22081_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _54516_ (_22082_, _22081_, _22080_);
  and _54517_ (_22083_, _22082_, _09792_);
  and _54518_ (_22084_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _54519_ (_22085_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _54520_ (_22086_, _22085_, _22084_);
  and _54521_ (_22087_, _22086_, _05549_);
  or _54522_ (_22088_, _22087_, _22083_);
  or _54523_ (_22089_, _22088_, _05535_);
  and _54524_ (_22090_, _22089_, _09805_);
  and _54525_ (_22091_, _22090_, _22079_);
  or _54526_ (_22092_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _54527_ (_22093_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _54528_ (_22094_, _22093_, _05549_);
  and _54529_ (_22095_, _22094_, _22092_);
  or _54530_ (_22096_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or _54531_ (_22097_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _54532_ (_22098_, _22097_, _09792_);
  and _54533_ (_22099_, _22098_, _22096_);
  or _54534_ (_22100_, _22099_, _22095_);
  or _54535_ (_22101_, _22100_, _09791_);
  or _54536_ (_22102_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or _54537_ (_22103_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _54538_ (_22104_, _22103_, _05549_);
  and _54539_ (_22105_, _22104_, _22102_);
  or _54540_ (_22106_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _54541_ (_22107_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and _54542_ (_22108_, _22107_, _09792_);
  and _54543_ (_22109_, _22108_, _22106_);
  or _54544_ (_22110_, _22109_, _22105_);
  or _54545_ (_22111_, _22110_, _05535_);
  and _54546_ (_22112_, _22111_, _05542_);
  and _54547_ (_22113_, _22112_, _22101_);
  or _54548_ (_22114_, _22113_, _22091_);
  and _54549_ (_22115_, _22114_, _09850_);
  or _54550_ (_22116_, _22115_, _22069_);
  and _54551_ (_22117_, _22116_, _09790_);
  and _54552_ (_22118_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and _54553_ (_22119_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _54554_ (_22120_, _22119_, _22118_);
  and _54555_ (_22121_, _22120_, _09792_);
  and _54556_ (_22122_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and _54557_ (_22123_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _54558_ (_22124_, _22123_, _22122_);
  and _54559_ (_22125_, _22124_, _05549_);
  or _54560_ (_22126_, _22125_, _22121_);
  and _54561_ (_22127_, _22126_, _05535_);
  and _54562_ (_22128_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and _54563_ (_22129_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or _54564_ (_22130_, _22129_, _22128_);
  and _54565_ (_22131_, _22130_, _09792_);
  and _54566_ (_22132_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and _54567_ (_22133_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or _54568_ (_22134_, _22133_, _22132_);
  and _54569_ (_22135_, _22134_, _05549_);
  or _54570_ (_22136_, _22135_, _22131_);
  and _54571_ (_22137_, _22136_, _09791_);
  or _54572_ (_22138_, _22137_, _22127_);
  and _54573_ (_22139_, _22138_, _09805_);
  or _54574_ (_22140_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or _54575_ (_22141_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _54576_ (_22142_, _22141_, _05549_);
  and _54577_ (_22143_, _22142_, _22140_);
  or _54578_ (_22144_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or _54579_ (_22145_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and _54580_ (_22146_, _22145_, _09792_);
  and _54581_ (_22147_, _22146_, _22144_);
  or _54582_ (_22148_, _22147_, _22143_);
  and _54583_ (_22149_, _22148_, _05535_);
  or _54584_ (_22150_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or _54585_ (_22151_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and _54586_ (_22152_, _22151_, _05549_);
  and _54587_ (_22153_, _22152_, _22150_);
  or _54588_ (_22154_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or _54589_ (_22155_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and _54590_ (_22156_, _22155_, _09792_);
  and _54591_ (_22157_, _22156_, _22154_);
  or _54592_ (_22158_, _22157_, _22153_);
  and _54593_ (_22159_, _22158_, _09791_);
  or _54594_ (_22160_, _22159_, _22149_);
  and _54595_ (_22161_, _22160_, _05542_);
  or _54596_ (_22162_, _22161_, _22139_);
  and _54597_ (_22163_, _22162_, _09850_);
  and _54598_ (_22164_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and _54599_ (_22165_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _54600_ (_22166_, _22165_, _22164_);
  and _54601_ (_22167_, _22166_, _09792_);
  and _54602_ (_22168_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _54603_ (_22169_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _54604_ (_22170_, _22169_, _22168_);
  and _54605_ (_22171_, _22170_, _05549_);
  or _54606_ (_22172_, _22171_, _22167_);
  and _54607_ (_22173_, _22172_, _05535_);
  and _54608_ (_22174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and _54609_ (_22175_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _54610_ (_22176_, _22175_, _22174_);
  and _54611_ (_22177_, _22176_, _09792_);
  and _54612_ (_22178_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and _54613_ (_22179_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _54614_ (_22180_, _22179_, _22178_);
  and _54615_ (_22181_, _22180_, _05549_);
  or _54616_ (_22182_, _22181_, _22177_);
  and _54617_ (_22183_, _22182_, _09791_);
  or _54618_ (_22184_, _22183_, _22173_);
  and _54619_ (_22185_, _22184_, _09805_);
  or _54620_ (_22186_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _54621_ (_22187_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and _54622_ (_22188_, _22187_, _22186_);
  and _54623_ (_22189_, _22188_, _09792_);
  or _54624_ (_22190_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _54625_ (_22191_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _54626_ (_22192_, _22191_, _22190_);
  and _54627_ (_22193_, _22192_, _05549_);
  or _54628_ (_22194_, _22193_, _22189_);
  and _54629_ (_22195_, _22194_, _05535_);
  or _54630_ (_22196_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _54631_ (_22197_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _54632_ (_22198_, _22197_, _22196_);
  and _54633_ (_22199_, _22198_, _09792_);
  or _54634_ (_22200_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _54635_ (_22201_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and _54636_ (_22202_, _22201_, _22200_);
  and _54637_ (_22203_, _22202_, _05549_);
  or _54638_ (_22204_, _22203_, _22199_);
  and _54639_ (_22205_, _22204_, _09791_);
  or _54640_ (_22206_, _22205_, _22195_);
  and _54641_ (_22207_, _22206_, _05542_);
  or _54642_ (_22208_, _22207_, _22185_);
  and _54643_ (_22209_, _22208_, _05518_);
  or _54644_ (_22210_, _22209_, _22163_);
  and _54645_ (_22211_, _22210_, _05520_);
  or _54646_ (_22212_, _22211_, _22117_);
  or _54647_ (_22213_, _22212_, _05526_);
  and _54648_ (_22214_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and _54649_ (_22215_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _54650_ (_22216_, _22215_, _22214_);
  and _54651_ (_22217_, _22216_, _09792_);
  and _54652_ (_22218_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and _54653_ (_22219_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _54654_ (_22220_, _22219_, _22218_);
  and _54655_ (_22221_, _22220_, _05549_);
  or _54656_ (_22222_, _22221_, _22217_);
  or _54657_ (_22223_, _22222_, _09791_);
  and _54658_ (_22224_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and _54659_ (_22225_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _54660_ (_22226_, _22225_, _22224_);
  and _54661_ (_22227_, _22226_, _09792_);
  and _54662_ (_22228_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and _54663_ (_22229_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _54664_ (_22230_, _22229_, _22228_);
  and _54665_ (_22231_, _22230_, _05549_);
  or _54666_ (_22232_, _22231_, _22227_);
  or _54667_ (_22233_, _22232_, _05535_);
  and _54668_ (_22234_, _22233_, _09805_);
  and _54669_ (_22235_, _22234_, _22223_);
  or _54670_ (_22236_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _54671_ (_22237_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and _54672_ (_22238_, _22237_, _05549_);
  and _54673_ (_22239_, _22238_, _22236_);
  or _54674_ (_22240_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _54675_ (_22241_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and _54676_ (_22242_, _22241_, _09792_);
  and _54677_ (_22243_, _22242_, _22240_);
  or _54678_ (_22244_, _22243_, _22239_);
  or _54679_ (_22245_, _22244_, _09791_);
  or _54680_ (_22246_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _54681_ (_22247_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and _54682_ (_22248_, _22247_, _05549_);
  and _54683_ (_22249_, _22248_, _22246_);
  or _54684_ (_22250_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _54685_ (_22251_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and _54686_ (_22252_, _22251_, _09792_);
  and _54687_ (_22253_, _22252_, _22250_);
  or _54688_ (_22254_, _22253_, _22249_);
  or _54689_ (_22255_, _22254_, _05535_);
  and _54690_ (_22256_, _22255_, _05542_);
  and _54691_ (_22257_, _22256_, _22245_);
  or _54692_ (_22258_, _22257_, _22235_);
  and _54693_ (_22259_, _22258_, _09850_);
  and _54694_ (_22260_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and _54695_ (_22261_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _54696_ (_22262_, _22261_, _22260_);
  and _54697_ (_22263_, _22262_, _09792_);
  and _54698_ (_22264_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _54699_ (_22265_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or _54700_ (_22266_, _22265_, _22264_);
  and _54701_ (_22267_, _22266_, _05549_);
  or _54702_ (_22268_, _22267_, _22263_);
  or _54703_ (_22269_, _22268_, _09791_);
  and _54704_ (_22270_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and _54705_ (_22271_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or _54706_ (_22272_, _22271_, _22270_);
  and _54707_ (_22273_, _22272_, _09792_);
  and _54708_ (_22274_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and _54709_ (_22275_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _54710_ (_22276_, _22275_, _22274_);
  and _54711_ (_22277_, _22276_, _05549_);
  or _54712_ (_22278_, _22277_, _22273_);
  or _54713_ (_22279_, _22278_, _05535_);
  and _54714_ (_22280_, _22279_, _09805_);
  and _54715_ (_22281_, _22280_, _22269_);
  or _54716_ (_22282_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _54717_ (_22283_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _54718_ (_22284_, _22283_, _22282_);
  and _54719_ (_22285_, _22284_, _09792_);
  or _54720_ (_22286_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _54721_ (_22287_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and _54722_ (_22288_, _22287_, _22286_);
  and _54723_ (_22289_, _22288_, _05549_);
  or _54724_ (_22290_, _22289_, _22285_);
  or _54725_ (_22291_, _22290_, _09791_);
  or _54726_ (_22292_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _54727_ (_22293_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _54728_ (_22294_, _22293_, _22292_);
  and _54729_ (_22295_, _22294_, _09792_);
  or _54730_ (_22296_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _54731_ (_22297_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _54732_ (_22298_, _22297_, _22296_);
  and _54733_ (_22299_, _22298_, _05549_);
  or _54734_ (_22300_, _22299_, _22295_);
  or _54735_ (_22301_, _22300_, _05535_);
  and _54736_ (_22302_, _22301_, _05542_);
  and _54737_ (_22303_, _22302_, _22291_);
  or _54738_ (_22304_, _22303_, _22281_);
  and _54739_ (_22305_, _22304_, _05518_);
  or _54740_ (_22306_, _22305_, _22259_);
  and _54741_ (_22307_, _22306_, _09790_);
  or _54742_ (_22308_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _54743_ (_22309_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _54744_ (_22310_, _22309_, _22308_);
  and _54745_ (_22311_, _22310_, _09792_);
  or _54746_ (_22312_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _54747_ (_22313_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and _54748_ (_22314_, _22313_, _22312_);
  and _54749_ (_22315_, _22314_, _05549_);
  or _54750_ (_22316_, _22315_, _22311_);
  and _54751_ (_22317_, _22316_, _09791_);
  or _54752_ (_22318_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _54753_ (_22319_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _54754_ (_22320_, _22319_, _22318_);
  and _54755_ (_22321_, _22320_, _09792_);
  or _54756_ (_22322_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or _54757_ (_22323_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _54758_ (_22324_, _22323_, _22322_);
  and _54759_ (_22325_, _22324_, _05549_);
  or _54760_ (_22326_, _22325_, _22321_);
  and _54761_ (_22327_, _22326_, _05535_);
  or _54762_ (_22328_, _22327_, _22317_);
  and _54763_ (_22329_, _22328_, _05542_);
  and _54764_ (_22330_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and _54765_ (_22331_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _54766_ (_22332_, _22331_, _22330_);
  and _54767_ (_22333_, _22332_, _09792_);
  and _54768_ (_22334_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _54769_ (_22335_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _54770_ (_22336_, _22335_, _22334_);
  and _54771_ (_22337_, _22336_, _05549_);
  or _54772_ (_22338_, _22337_, _22333_);
  and _54773_ (_22339_, _22338_, _09791_);
  and _54774_ (_22340_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _54775_ (_22341_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _54776_ (_22342_, _22341_, _22340_);
  and _54777_ (_22343_, _22342_, _09792_);
  and _54778_ (_22344_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _54779_ (_22345_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _54780_ (_22346_, _22345_, _22344_);
  and _54781_ (_22347_, _22346_, _05549_);
  or _54782_ (_22348_, _22347_, _22343_);
  and _54783_ (_22349_, _22348_, _05535_);
  or _54784_ (_22350_, _22349_, _22339_);
  and _54785_ (_22351_, _22350_, _09805_);
  or _54786_ (_22352_, _22351_, _22329_);
  and _54787_ (_22353_, _22352_, _05518_);
  or _54788_ (_22354_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or _54789_ (_22355_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and _54790_ (_22356_, _22355_, _05549_);
  and _54791_ (_22357_, _22356_, _22354_);
  or _54792_ (_22358_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _54793_ (_22359_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and _54794_ (_22360_, _22359_, _09792_);
  and _54795_ (_22361_, _22360_, _22358_);
  or _54796_ (_22362_, _22361_, _22357_);
  and _54797_ (_22363_, _22362_, _09791_);
  or _54798_ (_22364_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or _54799_ (_22365_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and _54800_ (_22366_, _22365_, _05549_);
  and _54801_ (_22367_, _22366_, _22364_);
  or _54802_ (_22368_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _54803_ (_22369_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and _54804_ (_22370_, _22369_, _09792_);
  and _54805_ (_22371_, _22370_, _22368_);
  or _54806_ (_22372_, _22371_, _22367_);
  and _54807_ (_22373_, _22372_, _05535_);
  or _54808_ (_22374_, _22373_, _22363_);
  and _54809_ (_22375_, _22374_, _05542_);
  and _54810_ (_22376_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and _54811_ (_22377_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _54812_ (_22378_, _22377_, _22376_);
  and _54813_ (_22379_, _22378_, _09792_);
  and _54814_ (_22380_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and _54815_ (_22381_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or _54816_ (_22382_, _22381_, _22380_);
  and _54817_ (_22383_, _22382_, _05549_);
  or _54818_ (_22384_, _22383_, _22379_);
  and _54819_ (_22385_, _22384_, _09791_);
  and _54820_ (_22386_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and _54821_ (_22387_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or _54822_ (_22388_, _22387_, _22386_);
  and _54823_ (_22389_, _22388_, _09792_);
  and _54824_ (_22390_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and _54825_ (_22391_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _54826_ (_22392_, _22391_, _22390_);
  and _54827_ (_22393_, _22392_, _05549_);
  or _54828_ (_22394_, _22393_, _22389_);
  and _54829_ (_22395_, _22394_, _05535_);
  or _54830_ (_22396_, _22395_, _22385_);
  and _54831_ (_22397_, _22396_, _09805_);
  or _54832_ (_22398_, _22397_, _22375_);
  and _54833_ (_22399_, _22398_, _09850_);
  or _54834_ (_22400_, _22399_, _22353_);
  and _54835_ (_22401_, _22400_, _05520_);
  or _54836_ (_22402_, _22401_, _22307_);
  or _54837_ (_22403_, _22402_, _10033_);
  and _54838_ (_22404_, _22403_, _22213_);
  or _54839_ (_22405_, _22404_, _04413_);
  and _54840_ (_22406_, _22405_, _22023_);
  or _54841_ (_22407_, _22406_, _05563_);
  or _54842_ (_22408_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and _54843_ (_22409_, _22408_, _22731_);
  and _54844_ (_12348_, _22409_, _22407_);
  and _54845_ (_22410_, _02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _54846_ (_22411_, _22410_, _02306_);
  and _54847_ (_22412_, _22411_, _02195_);
  nor _54848_ (_22413_, _22412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _54849_ (_22414_, _22412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _54850_ (_22415_, _22414_, _22413_);
  and _54851_ (_22416_, _22415_, _02198_);
  and _54852_ (_22417_, _01818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _54853_ (_22418_, _22417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _54854_ (_22419_, _11221_);
  and _54855_ (_22420_, _01829_, _22419_);
  and _54856_ (_22421_, _22420_, _22418_);
  or _54857_ (_22422_, _11203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _54858_ (_22423_, _11211_, _02320_);
  and _54859_ (_22424_, _22423_, _22422_);
  or _54860_ (_22425_, _22424_, _22421_);
  or _54861_ (_22426_, _22425_, _22416_);
  or _54862_ (_22427_, _22426_, _01814_);
  nand _54863_ (_22428_, _01814_, _23542_);
  and _54864_ (_22429_, _22428_, _22427_);
  or _54865_ (_22430_, _22429_, _01816_);
  or _54866_ (_22431_, _02300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _54867_ (_22432_, _22431_, _22731_);
  and _54868_ (_12351_, _22432_, _22430_);
  and _54869_ (_22433_, _02488_, _24134_);
  and _54870_ (_22434_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or _54871_ (_12353_, _22434_, _22433_);
  nand _54872_ (_22435_, _01814_, _24210_);
  and _54873_ (_22436_, _08225_, _02195_);
  or _54874_ (_22437_, _22436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _54875_ (_22438_, _11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _54876_ (_22439_, _22438_, _02198_);
  and _54877_ (_22440_, _22439_, _22437_);
  or _54878_ (_22441_, _01818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _54879_ (_22442_, _22441_, _01829_);
  nor _54880_ (_22443_, _22442_, _22417_);
  or _54881_ (_22444_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _54882_ (_22445_, _11203_, _02320_);
  and _54883_ (_22446_, _22445_, _22444_);
  or _54884_ (_22447_, _22446_, _22443_);
  or _54885_ (_22448_, _22447_, _22440_);
  or _54886_ (_22449_, _22448_, _01814_);
  and _54887_ (_22450_, _22449_, _22435_);
  or _54888_ (_22451_, _22450_, _01816_);
  or _54889_ (_22452_, _02300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _54890_ (_22453_, _22452_, _22731_);
  and _54891_ (_12355_, _22453_, _22451_);
  and _54892_ (_22454_, _12438_, _23996_);
  and _54893_ (_22455_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or _54894_ (_12357_, _22455_, _22454_);
  and _54895_ (_22456_, _12438_, _24219_);
  and _54896_ (_22457_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or _54897_ (_27190_, _22457_, _22456_);
  and _54898_ (_22458_, _16026_, _24219_);
  and _54899_ (_22459_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or _54900_ (_12369_, _22459_, _22458_);
  and _54901_ (_22460_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _54902_ (_22461_, _01814_, _24126_);
  and _54903_ (_22462_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _54904_ (_22463_, _22462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _54905_ (_22464_, _22462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _54906_ (_22465_, _22464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _54907_ (_22466_, _22465_, _22463_);
  and _54908_ (_22467_, _02210_, _02302_);
  or _54909_ (_22468_, _22467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _54910_ (_22469_, _02318_, _02320_);
  and _54911_ (_22470_, _22469_, _22468_);
  and _54912_ (_22471_, _08225_, _02302_);
  or _54913_ (_22472_, _22471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _54914_ (_22473_, _02308_, _02197_);
  and _54915_ (_22474_, _22473_, _22472_);
  or _54916_ (_22475_, _22474_, _22470_);
  or _54917_ (_22476_, _22475_, _22466_);
  or _54918_ (_22477_, _22476_, _01814_);
  and _54919_ (_22478_, _22477_, _02300_);
  and _54920_ (_22479_, _22478_, _22461_);
  or _54921_ (_22480_, _22479_, _22460_);
  and _54922_ (_12384_, _22480_, _22731_);
  and _54923_ (_22481_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _54924_ (_22482_, _01814_, _24043_);
  nand _54925_ (_22483_, _08225_, _01823_);
  nor _54926_ (_22484_, _22483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _54927_ (_22485_, _22484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not _54928_ (_22486_, _22471_);
  or _54929_ (_22487_, _22486_, _02196_);
  and _54930_ (_22488_, _22487_, _02198_);
  and _54931_ (_22489_, _22488_, _22485_);
  or _54932_ (_22490_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not _54933_ (_22491_, _01825_);
  and _54934_ (_22492_, _01829_, _22491_);
  and _54935_ (_22493_, _22492_, _22490_);
  and _54936_ (_22494_, _02210_, _01823_);
  or _54937_ (_22495_, _22494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _54938_ (_22496_, _22467_, _02320_);
  and _54939_ (_22497_, _22496_, _22495_);
  or _54940_ (_22498_, _22497_, _22493_);
  or _54941_ (_22499_, _22498_, _22489_);
  or _54942_ (_22500_, _22499_, _01814_);
  and _54943_ (_22501_, _22500_, _02300_);
  and _54944_ (_22502_, _22501_, _22482_);
  or _54945_ (_22503_, _22502_, _22481_);
  and _54946_ (_12387_, _22503_, _22731_);
  and _54947_ (_22504_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _54948_ (_22505_, _01814_, _24082_);
  and _54949_ (_22506_, _08225_, _01822_);
  or _54950_ (_22507_, _22506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _54951_ (_22508_, _22483_, _02197_);
  and _54952_ (_22509_, _22508_, _22507_);
  and _54953_ (_22510_, _02210_, _01822_);
  or _54954_ (_22511_, _22510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _54955_ (_22512_, _22494_, _02320_);
  and _54956_ (_22513_, _22512_, _22511_);
  and _54957_ (_22514_, _01822_, _01818_);
  and _54958_ (_22515_, _22514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _54959_ (_22516_, _22515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _54960_ (_22517_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _54961_ (_22518_, _22517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _54962_ (_22519_, _22518_, _22516_);
  or _54963_ (_22520_, _22519_, _22513_);
  or _54964_ (_22521_, _22520_, _22509_);
  or _54965_ (_22522_, _22521_, _01814_);
  and _54966_ (_22523_, _22522_, _02300_);
  and _54967_ (_22524_, _22523_, _22505_);
  or _54968_ (_22525_, _22524_, _22504_);
  and _54969_ (_12390_, _22525_, _22731_);
  not _54970_ (_22526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _54971_ (_22527_, _22414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _54972_ (_22528_, _22527_, _22526_);
  and _54973_ (_22529_, _22527_, _22526_);
  or _54974_ (_22530_, _22529_, _22528_);
  and _54975_ (_22531_, _22530_, _02198_);
  or _54976_ (_22532_, _11218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _54977_ (_22533_, _22514_);
  and _54978_ (_22534_, _01829_, _22533_);
  and _54979_ (_22535_, _22534_, _22532_);
  or _54980_ (_22536_, _11214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _54981_ (_22537_, _22510_, _02320_);
  and _54982_ (_22538_, _22537_, _22536_);
  or _54983_ (_22539_, _22538_, _22535_);
  or _54984_ (_22540_, _22539_, _01814_);
  or _54985_ (_22541_, _22540_, _22531_);
  or _54986_ (_22542_, _02193_, _23577_);
  and _54987_ (_22543_, _22542_, _22541_);
  or _54988_ (_22544_, _22543_, _01816_);
  nand _54989_ (_22545_, _01816_, _22526_);
  and _54990_ (_22546_, _22545_, _22731_);
  and _54991_ (_12391_, _22546_, _22544_);
  and _54992_ (_22547_, _25637_, _23583_);
  and _54993_ (_22548_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _54994_ (_12393_, _22548_, _22547_);
  and _54995_ (_22549_, _12438_, _23583_);
  and _54996_ (_22550_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or _54997_ (_12397_, _22550_, _22549_);
  and _54998_ (_22551_, _05442_, _24219_);
  and _54999_ (_22552_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _55000_ (_12399_, _22552_, _22551_);
  and _55001_ (_22553_, _03355_, _23583_);
  and _55002_ (_22554_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _55003_ (_12404_, _22554_, _22553_);
  and _55004_ (_22555_, _03033_, _23887_);
  and _55005_ (_22556_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or _55006_ (_27161_, _22556_, _22555_);
  or _55007_ (_22557_, _02300_, _23880_);
  nor _55008_ (_22558_, _11184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _55009_ (_22559_, _22558_, _11185_);
  and _55010_ (_22560_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _55011_ (_22561_, _22560_, _22559_);
  nor _55012_ (_22562_, _22561_, _01814_);
  and _55013_ (_22563_, _01814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _55014_ (_22564_, _22563_, _22562_);
  or _55015_ (_22565_, _22564_, _01816_);
  and _55016_ (_22566_, _22565_, _22731_);
  and _55017_ (_12412_, _22566_, _22557_);
  nand _55018_ (_22567_, _01816_, _23542_);
  and _55019_ (_22568_, _02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _55020_ (_22569_, _22568_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _55021_ (_22570_, _22569_, _11184_);
  and _55022_ (_22571_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _55023_ (_22572_, _22571_, _22570_);
  nor _55024_ (_22573_, _22572_, _01814_);
  and _55025_ (_22574_, _01814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _55026_ (_22575_, _22574_, _22573_);
  or _55027_ (_22576_, _22575_, _01816_);
  and _55028_ (_22577_, _22576_, _22731_);
  and _55029_ (_12413_, _22577_, _22567_);
  and _55030_ (_22578_, _02488_, _24051_);
  and _55031_ (_22579_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or _55032_ (_12416_, _22579_, _22578_);
  nor _55033_ (_22580_, _02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _55034_ (_22581_, _22580_, _22568_);
  and _55035_ (_22582_, _11205_, _02196_);
  nor _55036_ (_22583_, _22582_, _22581_);
  nor _55037_ (_22584_, _22583_, _01814_);
  and _55038_ (_22585_, _01814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or _55039_ (_22586_, _22585_, _22584_);
  or _55040_ (_22587_, _22586_, _01816_);
  nand _55041_ (_22588_, _01816_, _24210_);
  and _55042_ (_22589_, _22588_, _22731_);
  and _55043_ (_12417_, _22589_, _22587_);
  and _55044_ (_22590_, _02045_, _24219_);
  and _55045_ (_22591_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _55046_ (_12420_, _22591_, _22590_);
  and _55047_ (_22592_, _24510_, _24219_);
  and _55048_ (_22593_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _55049_ (_12422_, _22593_, _22592_);
  and _55050_ (_22594_, _24510_, _23583_);
  and _55051_ (_22595_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _55052_ (_12424_, _22595_, _22594_);
  and _55053_ (_22596_, _12429_, _24219_);
  and _55054_ (_22597_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or _55055_ (_27182_, _22597_, _22596_);
  nand _55056_ (_22598_, _01816_, _24082_);
  nand _55057_ (_22599_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _55058_ (_22600_, _02210_);
  nand _55059_ (_22601_, _11191_, _22600_);
  and _55060_ (_22602_, _22601_, _22599_);
  nor _55061_ (_22603_, _22602_, _01814_);
  or _55062_ (_22604_, _22600_, _01814_);
  and _55063_ (_22605_, _22604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _55064_ (_22606_, _22605_, _22603_);
  or _55065_ (_22607_, _22606_, _01816_);
  and _55066_ (_22608_, _22607_, _22731_);
  and _55067_ (_12432_, _22608_, _22598_);
  and _55068_ (_22609_, _03043_, _23996_);
  and _55069_ (_22610_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or _55070_ (_27252_, _22610_, _22609_);
  dff _55071_ (first_instr, _00000_, clk);
  dff _55072_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _26823_[0], clk);
  dff _55073_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _26823_[1], clk);
  dff _55074_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _26823_[2], clk);
  dff _55075_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _26823_[3], clk);
  dff _55076_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _26823_[4], clk);
  dff _55077_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _26823_[5], clk);
  dff _55078_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _26823_[6], clk);
  dff _55079_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _26823_[7], clk);
  dff _55080_ (\oc8051_symbolic_cxrom1.regvalid [0], _26839_, clk);
  dff _55081_ (\oc8051_symbolic_cxrom1.regvalid [1], _26822_[1], clk);
  dff _55082_ (\oc8051_symbolic_cxrom1.regvalid [2], _26822_[2], clk);
  dff _55083_ (\oc8051_symbolic_cxrom1.regvalid [3], _26822_[3], clk);
  dff _55084_ (\oc8051_symbolic_cxrom1.regvalid [4], _26822_[4], clk);
  dff _55085_ (\oc8051_symbolic_cxrom1.regvalid [5], _26822_[5], clk);
  dff _55086_ (\oc8051_symbolic_cxrom1.regvalid [6], _26822_[6], clk);
  dff _55087_ (\oc8051_symbolic_cxrom1.regvalid [7], _26822_[7], clk);
  dff _55088_ (\oc8051_symbolic_cxrom1.regvalid [8], _26822_[8], clk);
  dff _55089_ (\oc8051_symbolic_cxrom1.regvalid [9], _26822_[9], clk);
  dff _55090_ (\oc8051_symbolic_cxrom1.regvalid [10], _26822_[10], clk);
  dff _55091_ (\oc8051_symbolic_cxrom1.regvalid [11], _26822_[11], clk);
  dff _55092_ (\oc8051_symbolic_cxrom1.regvalid [12], _26822_[12], clk);
  dff _55093_ (\oc8051_symbolic_cxrom1.regvalid [13], _26822_[13], clk);
  dff _55094_ (\oc8051_symbolic_cxrom1.regvalid [14], _26822_[14], clk);
  dff _55095_ (\oc8051_symbolic_cxrom1.regvalid [15], _26822_[15], clk);
  dff _55096_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _26830_[0], clk);
  dff _55097_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _26830_[1], clk);
  dff _55098_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _26830_[2], clk);
  dff _55099_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _26830_[3], clk);
  dff _55100_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _26830_[4], clk);
  dff _55101_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _26830_[5], clk);
  dff _55102_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _26830_[6], clk);
  dff _55103_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _26830_[7], clk);
  dff _55104_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _26831_[0], clk);
  dff _55105_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _26831_[1], clk);
  dff _55106_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _26831_[2], clk);
  dff _55107_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _26831_[3], clk);
  dff _55108_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _26831_[4], clk);
  dff _55109_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _26831_[5], clk);
  dff _55110_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _26831_[6], clk);
  dff _55111_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _26831_[7], clk);
  dff _55112_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _26832_[0], clk);
  dff _55113_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _26832_[1], clk);
  dff _55114_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _26832_[2], clk);
  dff _55115_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _26832_[3], clk);
  dff _55116_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _26832_[4], clk);
  dff _55117_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _26832_[5], clk);
  dff _55118_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _26832_[6], clk);
  dff _55119_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _26832_[7], clk);
  dff _55120_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _26833_[0], clk);
  dff _55121_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _26833_[1], clk);
  dff _55122_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _26833_[2], clk);
  dff _55123_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _26833_[3], clk);
  dff _55124_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _26833_[4], clk);
  dff _55125_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _26833_[5], clk);
  dff _55126_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _26833_[6], clk);
  dff _55127_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _26833_[7], clk);
  dff _55128_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _26834_[0], clk);
  dff _55129_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _26834_[1], clk);
  dff _55130_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _26834_[2], clk);
  dff _55131_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _26834_[3], clk);
  dff _55132_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _26834_[4], clk);
  dff _55133_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _26834_[5], clk);
  dff _55134_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _26834_[6], clk);
  dff _55135_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _26834_[7], clk);
  dff _55136_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _26835_[0], clk);
  dff _55137_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _26835_[1], clk);
  dff _55138_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _26835_[2], clk);
  dff _55139_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _26835_[3], clk);
  dff _55140_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _26835_[4], clk);
  dff _55141_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _26835_[5], clk);
  dff _55142_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _26835_[6], clk);
  dff _55143_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _26835_[7], clk);
  dff _55144_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _26836_[0], clk);
  dff _55145_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _26836_[1], clk);
  dff _55146_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _26836_[2], clk);
  dff _55147_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _26836_[3], clk);
  dff _55148_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _26836_[4], clk);
  dff _55149_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _26836_[5], clk);
  dff _55150_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _26836_[6], clk);
  dff _55151_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _26836_[7], clk);
  dff _55152_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _26837_[0], clk);
  dff _55153_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _26837_[1], clk);
  dff _55154_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _26837_[2], clk);
  dff _55155_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _26837_[3], clk);
  dff _55156_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _26837_[4], clk);
  dff _55157_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _26837_[5], clk);
  dff _55158_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _26837_[6], clk);
  dff _55159_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _26837_[7], clk);
  dff _55160_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _26838_[0], clk);
  dff _55161_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _26838_[1], clk);
  dff _55162_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _26838_[2], clk);
  dff _55163_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _26838_[3], clk);
  dff _55164_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _26838_[4], clk);
  dff _55165_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _26838_[5], clk);
  dff _55166_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _26838_[6], clk);
  dff _55167_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _26838_[7], clk);
  dff _55168_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _26824_[0], clk);
  dff _55169_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _26824_[1], clk);
  dff _55170_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _26824_[2], clk);
  dff _55171_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _26824_[3], clk);
  dff _55172_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _26824_[4], clk);
  dff _55173_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _26824_[5], clk);
  dff _55174_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _26824_[6], clk);
  dff _55175_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _26824_[7], clk);
  dff _55176_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _26825_[0], clk);
  dff _55177_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _26825_[1], clk);
  dff _55178_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _26825_[2], clk);
  dff _55179_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _26825_[3], clk);
  dff _55180_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _26825_[4], clk);
  dff _55181_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _26825_[5], clk);
  dff _55182_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _26825_[6], clk);
  dff _55183_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _26825_[7], clk);
  dff _55184_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _26826_[0], clk);
  dff _55185_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _26826_[1], clk);
  dff _55186_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _26826_[2], clk);
  dff _55187_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _26826_[3], clk);
  dff _55188_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _26826_[4], clk);
  dff _55189_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _26826_[5], clk);
  dff _55190_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _26826_[6], clk);
  dff _55191_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _26826_[7], clk);
  dff _55192_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _26827_[0], clk);
  dff _55193_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _26827_[1], clk);
  dff _55194_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _26827_[2], clk);
  dff _55195_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _26827_[3], clk);
  dff _55196_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _26827_[4], clk);
  dff _55197_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _26827_[5], clk);
  dff _55198_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _26827_[6], clk);
  dff _55199_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _26827_[7], clk);
  dff _55200_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _26828_[0], clk);
  dff _55201_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _26828_[1], clk);
  dff _55202_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _26828_[2], clk);
  dff _55203_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _26828_[3], clk);
  dff _55204_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _26828_[4], clk);
  dff _55205_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _26828_[5], clk);
  dff _55206_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _26828_[6], clk);
  dff _55207_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _26828_[7], clk);
  dff _55208_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _26829_[0], clk);
  dff _55209_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _26829_[1], clk);
  dff _55210_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _26829_[2], clk);
  dff _55211_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _26829_[3], clk);
  dff _55212_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _26829_[4], clk);
  dff _55213_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _26829_[5], clk);
  dff _55214_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _26829_[6], clk);
  dff _55215_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _26829_[7], clk);
  dff _55216_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _11336_, clk);
  dff _55217_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _11315_, clk);
  dff _55218_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _09141_, clk);
  dff _55219_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _11283_, clk);
  dff _55220_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _11332_, clk);
  dff _55221_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _09148_, clk);
  dff _55222_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _09152_, clk);
  dff _55223_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _09133_, clk);
  dff _55224_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _11514_, clk);
  dff _55225_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11408_, clk);
  dff _55226_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _11487_, clk);
  dff _55227_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11475_, clk);
  dff _55228_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _11517_, clk);
  dff _55229_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _11510_, clk);
  dff _55230_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _11407_, clk);
  dff _55231_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _09145_, clk);
  dff _55232_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11708_, clk);
  dff _55233_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22676_, clk);
  dff _55234_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11721_, clk);
  dff _55235_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11934_, clk);
  dff _55236_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11726_, clk);
  dff _55237_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11738_, clk);
  dff _55238_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11716_, clk);
  dff _55239_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11728_, clk);
  dff _55240_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11734_, clk);
  dff _55241_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _11740_, clk);
  dff _55242_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11736_, clk);
  dff _55243_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11730_, clk);
  dff _55244_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11723_, clk);
  dff _55245_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11746_, clk);
  dff _55246_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11742_, clk);
  dff _55247_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11776_, clk);
  dff _55248_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _26840_[0], clk);
  dff _55249_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _26840_[1], clk);
  dff _55250_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _26840_[2], clk);
  dff _55251_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _26840_[3], clk);
  dff _55252_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _26840_[4], clk);
  dff _55253_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _26840_[5], clk);
  dff _55254_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _26840_[6], clk);
  dff _55255_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _26840_[7], clk);
  dff _55256_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _26867_[0], clk);
  dff _55257_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _26867_[1], clk);
  dff _55258_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _26867_[2], clk);
  dff _55259_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _26867_[3], clk);
  dff _55260_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _26867_[4], clk);
  dff _55261_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _26867_[5], clk);
  dff _55262_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _26867_[6], clk);
  dff _55263_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _26867_[7], clk);
  dff _55264_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _26877_[0], clk);
  dff _55265_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _26877_[1], clk);
  dff _55266_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _26877_[2], clk);
  dff _55267_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _26877_[3], clk);
  dff _55268_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _26877_[4], clk);
  dff _55269_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _26877_[5], clk);
  dff _55270_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _26877_[6], clk);
  dff _55271_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _26877_[7], clk);
  dff _55272_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _26847_[0], clk);
  dff _55273_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _26847_[1], clk);
  dff _55274_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _26848_[0], clk);
  dff _55275_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _26848_[1], clk);
  dff _55276_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _26848_[2], clk);
  dff _55277_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _26849_[0], clk);
  dff _55278_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _26849_[1], clk);
  dff _55279_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _26849_[2], clk);
  dff _55280_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _26850_[0], clk);
  dff _55281_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _26850_[1], clk);
  dff _55282_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _26851_[0], clk);
  dff _55283_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _26851_[1], clk);
  dff _55284_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _26851_[2], clk);
  dff _55285_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _26851_[3], clk);
  dff _55286_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _26852_[0], clk);
  dff _55287_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _26852_[1], clk);
  dff _55288_ (\oc8051_top_1.oc8051_decoder1.wr , _26853_, clk);
  dff _55289_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _26841_[0], clk);
  dff _55290_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _26841_[1], clk);
  dff _55291_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _26841_[2], clk);
  dff _55292_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _26842_[0], clk);
  dff _55293_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _26842_[1], clk);
  dff _55294_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _26842_[2], clk);
  dff _55295_ (\oc8051_top_1.oc8051_decoder1.state [0], _26843_[0], clk);
  dff _55296_ (\oc8051_top_1.oc8051_decoder1.state [1], _26843_[1], clk);
  dff _55297_ (\oc8051_top_1.oc8051_decoder1.op [0], _26844_[0], clk);
  dff _55298_ (\oc8051_top_1.oc8051_decoder1.op [1], _26844_[1], clk);
  dff _55299_ (\oc8051_top_1.oc8051_decoder1.op [2], _26844_[2], clk);
  dff _55300_ (\oc8051_top_1.oc8051_decoder1.op [3], _26844_[3], clk);
  dff _55301_ (\oc8051_top_1.oc8051_decoder1.op [4], _26844_[4], clk);
  dff _55302_ (\oc8051_top_1.oc8051_decoder1.op [5], _26844_[5], clk);
  dff _55303_ (\oc8051_top_1.oc8051_decoder1.op [6], _26844_[6], clk);
  dff _55304_ (\oc8051_top_1.oc8051_decoder1.op [7], _26844_[7], clk);
  dff _55305_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _26845_, clk);
  dff _55306_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _26846_[0], clk);
  dff _55307_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _26846_[1], clk);
  dff _55308_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _26892_, clk);
  dff _55309_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _26854_[0], clk);
  dff _55310_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _26854_[1], clk);
  dff _55311_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _26854_[2], clk);
  dff _55312_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _26854_[3], clk);
  dff _55313_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _26854_[4], clk);
  dff _55314_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _26854_[5], clk);
  dff _55315_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _26854_[6], clk);
  dff _55316_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _26854_[7], clk);
  dff _55317_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _26855_[0], clk);
  dff _55318_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _26855_[1], clk);
  dff _55319_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _26855_[2], clk);
  dff _55320_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _26855_[3], clk);
  dff _55321_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _26855_[4], clk);
  dff _55322_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _26855_[5], clk);
  dff _55323_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _26855_[6], clk);
  dff _55324_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _26855_[7], clk);
  dff _55325_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _26856_[0], clk);
  dff _55326_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _26856_[1], clk);
  dff _55327_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _26856_[2], clk);
  dff _55328_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _26856_[3], clk);
  dff _55329_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _26856_[4], clk);
  dff _55330_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _26856_[5], clk);
  dff _55331_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _26856_[6], clk);
  dff _55332_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _26856_[7], clk);
  dff _55333_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _26857_[0], clk);
  dff _55334_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _26857_[1], clk);
  dff _55335_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _26857_[2], clk);
  dff _55336_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _26857_[3], clk);
  dff _55337_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _26857_[4], clk);
  dff _55338_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _26857_[5], clk);
  dff _55339_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _26857_[6], clk);
  dff _55340_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _26857_[7], clk);
  dff _55341_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _26858_[0], clk);
  dff _55342_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _26858_[1], clk);
  dff _55343_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _26858_[2], clk);
  dff _55344_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _26858_[3], clk);
  dff _55345_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _26858_[4], clk);
  dff _55346_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _26858_[5], clk);
  dff _55347_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _26858_[6], clk);
  dff _55348_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _26858_[7], clk);
  dff _55349_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _26859_[0], clk);
  dff _55350_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _26859_[1], clk);
  dff _55351_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _26859_[2], clk);
  dff _55352_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _26859_[3], clk);
  dff _55353_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _26859_[4], clk);
  dff _55354_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _26859_[5], clk);
  dff _55355_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _26859_[6], clk);
  dff _55356_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _26859_[7], clk);
  dff _55357_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _26860_[0], clk);
  dff _55358_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _26860_[1], clk);
  dff _55359_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _26860_[2], clk);
  dff _55360_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _26860_[3], clk);
  dff _55361_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _26860_[4], clk);
  dff _55362_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _26860_[5], clk);
  dff _55363_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _26860_[6], clk);
  dff _55364_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _26860_[7], clk);
  dff _55365_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _26861_[0], clk);
  dff _55366_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _26861_[1], clk);
  dff _55367_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _26861_[2], clk);
  dff _55368_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _26861_[3], clk);
  dff _55369_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _26861_[4], clk);
  dff _55370_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _26861_[5], clk);
  dff _55371_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _26861_[6], clk);
  dff _55372_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _26861_[7], clk);
  dff _55373_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _26865_[0], clk);
  dff _55374_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _26865_[1], clk);
  dff _55375_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _26865_[2], clk);
  dff _55376_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _26865_[3], clk);
  dff _55377_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _26865_[4], clk);
  dff _55378_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _26862_[0], clk);
  dff _55379_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _26862_[1], clk);
  dff _55380_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _26862_[2], clk);
  dff _55381_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _26862_[3], clk);
  dff _55382_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _26862_[4], clk);
  dff _55383_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _26862_[5], clk);
  dff _55384_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _26862_[6], clk);
  dff _55385_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _26862_[7], clk);
  dff _55386_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _26862_[8], clk);
  dff _55387_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _26862_[9], clk);
  dff _55388_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _26862_[10], clk);
  dff _55389_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _26862_[11], clk);
  dff _55390_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _26862_[12], clk);
  dff _55391_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _26862_[13], clk);
  dff _55392_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _26862_[14], clk);
  dff _55393_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _26862_[15], clk);
  dff _55394_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _26863_[0], clk);
  dff _55395_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26863_[1], clk);
  dff _55396_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26863_[2], clk);
  dff _55397_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _26863_[3], clk);
  dff _55398_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _26863_[4], clk);
  dff _55399_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _26863_[5], clk);
  dff _55400_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _26863_[6], clk);
  dff _55401_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _26863_[7], clk);
  dff _55402_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _26863_[8], clk);
  dff _55403_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _26863_[9], clk);
  dff _55404_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _26863_[10], clk);
  dff _55405_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26863_[11], clk);
  dff _55406_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _26863_[12], clk);
  dff _55407_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _26863_[13], clk);
  dff _55408_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _26863_[14], clk);
  dff _55409_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _26863_[15], clk);
  dff _55410_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _26883_[0], clk);
  dff _55411_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _26883_[1], clk);
  dff _55412_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _26883_[2], clk);
  dff _55413_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _26883_[3], clk);
  dff _55414_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _26883_[4], clk);
  dff _55415_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _26883_[5], clk);
  dff _55416_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _26883_[6], clk);
  dff _55417_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _26883_[7], clk);
  dff _55418_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _26883_[8], clk);
  dff _55419_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _26883_[9], clk);
  dff _55420_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _26883_[10], clk);
  dff _55421_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _26883_[11], clk);
  dff _55422_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _26883_[12], clk);
  dff _55423_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _26883_[13], clk);
  dff _55424_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _26883_[14], clk);
  dff _55425_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _26883_[15], clk);
  dff _55426_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _26883_[16], clk);
  dff _55427_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _26883_[17], clk);
  dff _55428_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _26883_[18], clk);
  dff _55429_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _26883_[19], clk);
  dff _55430_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _26883_[20], clk);
  dff _55431_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _26883_[21], clk);
  dff _55432_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _26883_[22], clk);
  dff _55433_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _26883_[23], clk);
  dff _55434_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _26883_[24], clk);
  dff _55435_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _26883_[25], clk);
  dff _55436_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _26883_[26], clk);
  dff _55437_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _26883_[27], clk);
  dff _55438_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _26883_[28], clk);
  dff _55439_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _26883_[29], clk);
  dff _55440_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _26883_[30], clk);
  dff _55441_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _26883_[31], clk);
  dff _55442_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _26864_, clk);
  dff _55443_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _26866_[0], clk);
  dff _55444_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _26866_[1], clk);
  dff _55445_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _26866_[2], clk);
  dff _55446_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _26866_[3], clk);
  dff _55447_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _26866_[4], clk);
  dff _55448_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _26866_[5], clk);
  dff _55449_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _26866_[6], clk);
  dff _55450_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _26866_[7], clk);
  dff _55451_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _26868_, clk);
  dff _55452_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _26869_, clk);
  dff _55453_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _26870_[0], clk);
  dff _55454_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _26870_[1], clk);
  dff _55455_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _26870_[2], clk);
  dff _55456_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _26870_[3], clk);
  dff _55457_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _26870_[4], clk);
  dff _55458_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _26870_[5], clk);
  dff _55459_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _26870_[6], clk);
  dff _55460_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _26870_[7], clk);
  dff _55461_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _26870_[8], clk);
  dff _55462_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _26870_[9], clk);
  dff _55463_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _26870_[10], clk);
  dff _55464_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _26870_[11], clk);
  dff _55465_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _26870_[12], clk);
  dff _55466_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _26870_[13], clk);
  dff _55467_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _26870_[14], clk);
  dff _55468_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _26870_[15], clk);
  dff _55469_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _26871_[0], clk);
  dff _55470_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _26871_[1], clk);
  dff _55471_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _26871_[2], clk);
  dff _55472_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _26871_[3], clk);
  dff _55473_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _26871_[4], clk);
  dff _55474_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _26871_[5], clk);
  dff _55475_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _26871_[6], clk);
  dff _55476_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _26871_[7], clk);
  dff _55477_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _26871_[8], clk);
  dff _55478_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _26871_[9], clk);
  dff _55479_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _26871_[10], clk);
  dff _55480_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _26871_[11], clk);
  dff _55481_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _26871_[12], clk);
  dff _55482_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _26871_[13], clk);
  dff _55483_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _26871_[14], clk);
  dff _55484_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _26871_[15], clk);
  dff _55485_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _26872_, clk);
  dff _55486_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _26874_, clk);
  dff _55487_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _26873_, clk);
  dff _55488_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _26875_[0], clk);
  dff _55489_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _26875_[1], clk);
  dff _55490_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _26875_[2], clk);
  dff _55491_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _26875_[3], clk);
  dff _55492_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _26875_[4], clk);
  dff _55493_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _26875_[5], clk);
  dff _55494_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _26875_[6], clk);
  dff _55495_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _26875_[7], clk);
  dff _55496_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _26876_[0], clk);
  dff _55497_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26876_[1], clk);
  dff _55498_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _26876_[2], clk);
  dff _55499_ (\oc8051_top_1.oc8051_memory_interface1.reti , _26878_, clk);
  dff _55500_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _26879_[0], clk);
  dff _55501_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _26879_[1], clk);
  dff _55502_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _26879_[2], clk);
  dff _55503_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _26879_[3], clk);
  dff _55504_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _26879_[4], clk);
  dff _55505_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _26879_[5], clk);
  dff _55506_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _26879_[6], clk);
  dff _55507_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _26879_[7], clk);
  dff _55508_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _26880_, clk);
  dff _55509_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _26881_, clk);
  dff _55510_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _26882_[0], clk);
  dff _55511_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _26882_[1], clk);
  dff _55512_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _26882_[2], clk);
  dff _55513_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _26882_[3], clk);
  dff _55514_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _26884_[0], clk);
  dff _55515_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _26884_[1], clk);
  dff _55516_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _26884_[2], clk);
  dff _55517_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _26884_[3], clk);
  dff _55518_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _26884_[4], clk);
  dff _55519_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _26884_[5], clk);
  dff _55520_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _26884_[6], clk);
  dff _55521_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _26884_[7], clk);
  dff _55522_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _26884_[8], clk);
  dff _55523_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _26884_[9], clk);
  dff _55524_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _26884_[10], clk);
  dff _55525_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _26884_[11], clk);
  dff _55526_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _26884_[12], clk);
  dff _55527_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _26884_[13], clk);
  dff _55528_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _26884_[14], clk);
  dff _55529_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _26884_[15], clk);
  dff _55530_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _26884_[16], clk);
  dff _55531_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _26884_[17], clk);
  dff _55532_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _26884_[18], clk);
  dff _55533_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _26884_[19], clk);
  dff _55534_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _26884_[20], clk);
  dff _55535_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _26884_[21], clk);
  dff _55536_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _26884_[22], clk);
  dff _55537_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _26884_[23], clk);
  dff _55538_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _26884_[24], clk);
  dff _55539_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _26884_[25], clk);
  dff _55540_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _26884_[26], clk);
  dff _55541_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _26884_[27], clk);
  dff _55542_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _26884_[28], clk);
  dff _55543_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _26884_[29], clk);
  dff _55544_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _26884_[30], clk);
  dff _55545_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _26884_[31], clk);
  dff _55546_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _26885_, clk);
  dff _55547_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _26886_, clk);
  dff _55548_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _26887_, clk);
  dff _55549_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _26888_[0], clk);
  dff _55550_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _26888_[1], clk);
  dff _55551_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _26888_[2], clk);
  dff _55552_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _26888_[3], clk);
  dff _55553_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _26889_, clk);
  dff _55554_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _26890_, clk);
  dff _55555_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26891_[0], clk);
  dff _55556_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26891_[1], clk);
  dff _55557_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26891_[2], clk);
  dff _55558_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26891_[3], clk);
  dff _55559_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26891_[4], clk);
  dff _55560_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26891_[5], clk);
  dff _55561_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26891_[6], clk);
  dff _55562_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _26891_[7], clk);
  dff _55563_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _26893_[0], clk);
  dff _55564_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _26893_[1], clk);
  dff _55565_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _26893_[2], clk);
  dff _55566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _23339_, clk);
  dff _55567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _26970_, clk);
  dff _55568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _23165_, clk);
  dff _55569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _23153_, clk);
  dff _55570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _11688_, clk);
  dff _55571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _26971_, clk);
  dff _55572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _26972_, clk);
  dff _55573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _23014_, clk);
  dff _55574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _23431_, clk);
  dff _55575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _26951_, clk);
  dff _55576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _23435_, clk);
  dff _55577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _11292_, clk);
  dff _55578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _11440_, clk);
  dff _55579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _11455_, clk);
  dff _55580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _23303_, clk);
  dff _55581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _26952_, clk);
  dff _55582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _23725_, clk);
  dff _55583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _26932_, clk);
  dff _55584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _23866_, clk);
  dff _55585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _23849_, clk);
  dff _55586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _11661_, clk);
  dff _55587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _23394_, clk);
  dff _55588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _23389_, clk);
  dff _55589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _26933_, clk);
  dff _55590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _23956_, clk);
  dff _55591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _23942_, clk);
  dff _55592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _26917_, clk);
  dff _55593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _24010_, clk);
  dff _55594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _24046_, clk);
  dff _55595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _24012_, clk);
  dff _55596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _11294_, clk);
  dff _55597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _23678_, clk);
  dff _55598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _22955_, clk);
  dff _55599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _23046_, clk);
  dff _55600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _23077_, clk);
  dff _55601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _11289_, clk);
  dff _55602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _22770_, clk);
  dff _55603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _26986_, clk);
  dff _55604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _22729_, clk);
  dff _55605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _22873_, clk);
  dff _55606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _11296_, clk);
  dff _55607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _27311_, clk);
  dff _55608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _24090_, clk);
  dff _55609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _11656_, clk);
  dff _55610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _27312_, clk);
  dff _55611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _24168_, clk);
  dff _55612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _24138_, clk);
  dff _55613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _11638_, clk);
  dff _55614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _04945_, clk);
  dff _55615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _27171_, clk);
  dff _55616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _10382_, clk);
  dff _55617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _10250_, clk);
  dff _55618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _11792_, clk);
  dff _55619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _05029_, clk);
  dff _55620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _05024_, clk);
  dff _55621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _05093_, clk);
  dff _55622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _27154_, clk);
  dff _55623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _10796_, clk);
  dff _55624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _10780_, clk);
  dff _55625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _10764_, clk);
  dff _55626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _11778_, clk);
  dff _55627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _11161_, clk);
  dff _55628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _27155_, clk);
  dff _55629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _27156_, clk);
  dff _55630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _12637_, clk);
  dff _55631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _15619_, clk);
  dff _55632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _15213_, clk);
  dff _55633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _11761_, clk);
  dff _55634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _27122_, clk);
  dff _55635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _11589_, clk);
  dff _55636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _12266_, clk);
  dff _55637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _12243_, clk);
  dff _55638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _09970_, clk);
  dff _55639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _07588_, clk);
  dff _55640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _08947_, clk);
  dff _55641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _27209_, clk);
  dff _55642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _10001_, clk);
  dff _55643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _04842_, clk);
  dff _55644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _27210_, clk);
  dff _55645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _11526_, clk);
  dff _55646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _08369_, clk);
  dff _55647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _08381_, clk);
  dff _55648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _27207_, clk);
  dff _55649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _27208_, clk);
  dff _55650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _22681_, clk);
  dff _55651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _08629_, clk);
  dff _55652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _08634_, clk);
  dff _55653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _09980_, clk);
  dff _55654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _27205_, clk);
  dff _55655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _26065_, clk);
  dff _55656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _11383_, clk);
  dff _55657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _07499_, clk);
  dff _55658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _06869_, clk);
  dff _55659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _21620_, clk);
  dff _55660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _09230_, clk);
  dff _55661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _27206_, clk);
  dff _55662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _09896_, clk);
  dff _55663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _27203_, clk);
  dff _55664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _09891_, clk);
  dff _55665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _03584_, clk);
  dff _55666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _27204_, clk);
  dff _55667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _06614_, clk);
  dff _55668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _07503_, clk);
  dff _55669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _03063_, clk);
  dff _55670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _09600_, clk);
  dff _55671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _09745_, clk);
  dff _55672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _11081_, clk);
  dff _55673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _09809_, clk);
  dff _55674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _11077_, clk);
  dff _55675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _09986_, clk);
  dff _55676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _11215_, clk);
  dff _55677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _27202_, clk);
  dff _55678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _11237_, clk);
  dff _55679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _27201_, clk);
  dff _55680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _09448_, clk);
  dff _55681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _11088_, clk);
  dff _55682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _09479_, clk);
  dff _55683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _11085_, clk);
  dff _55684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _09499_, clk);
  dff _55685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _11176_, clk);
  dff _55686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _11180_, clk);
  dff _55687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _09008_, clk);
  dff _55688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _11103_, clk);
  dff _55689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _09032_, clk);
  dff _55690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _11178_, clk);
  dff _55691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _09093_, clk);
  dff _55692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _27200_, clk);
  dff _55693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _11091_, clk);
  dff _55694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _27197_, clk);
  dff _55695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _11240_, clk);
  dff _55696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _08606_, clk);
  dff _55697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _11106_, clk);
  dff _55698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _27198_, clk);
  dff _55699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _27199_, clk);
  dff _55700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _08724_, clk);
  dff _55701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _08971_, clk);
  dff _55702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _08294_, clk);
  dff _55703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _11190_, clk);
  dff _55704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _08378_, clk);
  dff _55705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _11109_, clk);
  dff _55706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _08397_, clk);
  dff _55707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _11188_, clk);
  dff _55708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _08490_, clk);
  dff _55709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _27196_, clk);
  dff _55710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _08087_, clk);
  dff _55711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _11115_, clk);
  dff _55712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _11222_, clk);
  dff _55713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _08123_, clk);
  dff _55714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _11113_, clk);
  dff _55715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _08142_, clk);
  dff _55716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _11192_, clk);
  dff _55717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _08169_, clk);
  dff _55718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _07645_, clk);
  dff _55719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _07762_, clk);
  dff _55720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _11121_, clk);
  dff _55721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _11224_, clk);
  dff _55722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _07812_, clk);
  dff _55723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _07923_, clk);
  dff _55724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _11117_, clk);
  dff _55725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _07944_, clk);
  dff _55726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _27305_, clk);
  dff _55727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _07972_, clk);
  dff _55728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _27306_, clk);
  dff _55729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _08275_, clk);
  dff _55730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _27307_, clk);
  dff _55731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _27308_, clk);
  dff _55732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _10812_, clk);
  dff _55733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _07968_, clk);
  dff _55734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _27300_, clk);
  dff _55735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _27301_, clk);
  dff _55736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _10720_, clk);
  dff _55737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _27302_, clk);
  dff _55738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _07975_, clk);
  dff _55739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _08814_, clk);
  dff _55740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _27303_, clk);
  dff _55741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _27304_, clk);
  dff _55742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _10607_, clk);
  dff _55743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _27299_, clk);
  dff _55744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _07983_, clk);
  dff _55745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _10656_, clk);
  dff _55746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _07981_, clk);
  dff _55747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _10671_, clk);
  dff _55748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _08290_, clk);
  dff _55749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _10688_, clk);
  dff _55750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _10534_, clk);
  dff _55751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _10562_, clk);
  dff _55752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _07990_, clk);
  dff _55753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _10583_, clk);
  dff _55754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _07988_, clk);
  dff _55755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _27298_, clk);
  dff _55756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _08694_, clk);
  dff _55757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _08855_, clk);
  dff _55758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _07997_, clk);
  dff _55759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _10379_, clk);
  dff _55760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _10446_, clk);
  dff _55761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _07995_, clk);
  dff _55762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _27296_, clk);
  dff _55763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _07993_, clk);
  dff _55764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _10508_, clk);
  dff _55765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _27297_, clk);
  dff _55766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _10173_, clk);
  dff _55767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _27295_, clk);
  dff _55768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _08005_, clk);
  dff _55769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _10186_, clk);
  dff _55770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _10196_, clk);
  dff _55771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _10242_, clk);
  dff _55772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _08002_, clk);
  dff _55773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _10260_, clk);
  dff _55774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _08851_, clk);
  dff _55775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _09770_, clk);
  dff _55776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _27292_, clk);
  dff _55777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _09844_, clk);
  dff _55778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _08247_, clk);
  dff _55779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _27293_, clk);
  dff _55780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _08809_, clk);
  dff _55781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _27294_, clk);
  dff _55782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _10115_, clk);
  dff _55783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _08799_, clk);
  dff _55784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _10126_, clk);
  dff _55785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _10140_, clk);
  dff _55786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _09226_, clk);
  dff _55787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _27291_, clk);
  dff _55788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _09748_, clk);
  dff _55789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _09211_, clk);
  dff _55790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _03196_, clk);
  dff _55791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _06574_, clk);
  dff _55792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _27246_, clk);
  dff _55793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _27247_, clk);
  dff _55794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _22743_, clk);
  dff _55795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _22787_, clk);
  dff _55796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _22677_, clk);
  dff _55797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _22679_, clk);
  dff _55798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _08847_, clk);
  dff _55799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _10040_, clk);
  dff _55800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _10061_, clk);
  dff _55801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _08802_, clk);
  dff _55802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _10070_, clk);
  dff _55803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _27287_, clk);
  dff _55804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _08012_, clk);
  dff _55805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _27288_, clk);
  dff _55806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _10428_, clk);
  dff _55807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _26904_, clk);
  dff _55808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _10461_, clk);
  dff _55809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _10523_, clk);
  dff _55810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _08932_, clk);
  dff _55811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _09180_, clk);
  dff _55812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _10528_, clk);
  dff _55813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _26905_, clk);
  dff _55814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _08986_, clk);
  dff _55815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _10201_, clk);
  dff _55816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _09112_, clk);
  dff _55817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _26902_, clk);
  dff _55818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _10337_, clk);
  dff _55819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _26903_, clk);
  dff _55820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _09198_, clk);
  dff _55821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _10375_, clk);
  dff _55822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _10166_, clk);
  dff _55823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _08992_, clk);
  dff _55824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _10170_, clk);
  dff _55825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _09113_, clk);
  dff _55826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _10179_, clk);
  dff _55827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _26901_, clk);
  dff _55828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _08989_, clk);
  dff _55829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _09183_, clk);
  dff _55830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _09191_, clk);
  dff _55831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _09768_, clk);
  dff _55832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _09810_, clk);
  dff _55833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _09048_, clk);
  dff _55834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _26899_, clk);
  dff _55835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _26900_, clk);
  dff _55836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _09854_, clk);
  dff _55837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _09130_, clk);
  dff _55838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _10964_, clk);
  dff _55839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _22616_, clk);
  dff _55840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _22688_, clk);
  dff _55841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _11056_, clk);
  dff _55842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _23972_, clk);
  dff _55843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _26923_, clk);
  dff _55844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _11011_, clk);
  dff _55845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _23949_, clk);
  dff _55846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _10978_, clk);
  dff _55847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _22611_, clk);
  dff _55848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _08728_, clk);
  dff _55849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _05116_, clk);
  dff _55850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _10933_, clk);
  dff _55851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _08393_, clk);
  dff _55852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _22620_, clk);
  dff _55853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _10967_, clk);
  dff _55854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _26921_, clk);
  dff _55855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _11030_, clk);
  dff _55856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _23787_, clk);
  dff _55857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _26922_, clk);
  dff _55858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _10951_, clk);
  dff _55859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _10944_, clk);
  dff _55860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _10980_, clk);
  dff _55861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _10993_, clk);
  dff _55862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _24326_, clk);
  dff _55863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _27176_, clk);
  dff _55864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _26004_, clk);
  dff _55865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _27177_, clk);
  dff _55866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _06994_, clk);
  dff _55867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _26026_, clk);
  dff _55868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _26009_, clk);
  dff _55869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _24429_, clk);
  dff _55870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _25883_, clk);
  dff _55871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _24483_, clk);
  dff _55872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _25972_, clk);
  dff _55873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _04929_, clk);
  dff _55874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _25966_, clk);
  dff _55875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _22724_, clk);
  dff _55876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _23502_, clk);
  dff _55877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _22668_, clk);
  dff _55878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _25927_, clk);
  dff _55879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _10560_, clk);
  dff _55880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _10899_, clk);
  dff _55881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _25953_, clk);
  dff _55882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _24432_, clk);
  dff _55883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _25993_, clk);
  dff _55884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _24423_, clk);
  dff _55885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _02554_, clk);
  dff _55886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _07425_, clk);
  dff _55887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _27174_, clk);
  dff _55888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _07399_, clk);
  dff _55889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _01662_, clk);
  dff _55890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _24390_, clk);
  dff _55891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _24498_, clk);
  dff _55892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _11442_, clk);
  dff _55893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _27175_, clk);
  dff _55894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _07511_, clk);
  dff _55895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _07501_, clk);
  dff _55896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _07550_, clk);
  dff _55897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _27172_, clk);
  dff _55898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _07554_, clk);
  dff _55899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _24191_, clk);
  dff _55900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _27173_, clk);
  dff _55901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _07306_, clk);
  dff _55902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _27169_, clk);
  dff _55903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _24199_, clk);
  dff _55904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _07868_, clk);
  dff _55905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _07646_, clk);
  dff _55906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _27170_, clk);
  dff _55907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _08240_, clk);
  dff _55908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _07904_, clk);
  dff _55909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _24195_, clk);
  dff _55910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _09224_, clk);
  dff _55911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _09220_, clk);
  dff _55912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _09159_, clk);
  dff _55913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _24205_, clk);
  dff _55914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _08272_, clk);
  dff _55915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _08261_, clk);
  dff _55916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _08256_, clk);
  dff _55917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _08903_, clk);
  dff _55918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _24222_, clk);
  dff _55919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _27166_, clk);
  dff _55920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _27167_, clk);
  dff _55921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _27168_, clk);
  dff _55922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _00541_, clk);
  dff _55923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _09061_, clk);
  dff _55924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _09059_, clk);
  dff _55925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _09004_, clk);
  dff _55926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _10705_, clk);
  dff _55927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _10703_, clk);
  dff _55928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _00302_, clk);
  dff _55929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _10810_, clk);
  dff _55930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _24227_, clk);
  dff _55931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _10175_, clk);
  dff _55932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _00527_, clk);
  dff _55933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _27165_, clk);
  dff _55934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _24241_, clk);
  dff _55935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _11111_, clk);
  dff _55936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _27164_, clk);
  dff _55937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _11199_, clk);
  dff _55938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _10915_, clk);
  dff _55939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _10893_, clk);
  dff _55940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _10982_, clk);
  dff _55941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _00215_, clk);
  dff _55942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _11539_, clk);
  dff _55943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _11605_, clk);
  dff _55944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _11711_, clk);
  dff _55945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _11685_, clk);
  dff _55946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _26105_, clk);
  dff _55947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _11331_, clk);
  dff _55948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _27163_, clk);
  dff _55949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _11436_, clk);
  dff _55950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _12334_, clk);
  dff _55951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _12340_, clk);
  dff _55952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _24280_, clk);
  dff _55953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _11906_, clk);
  dff _55954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _12092_, clk);
  dff _55955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _11937_, clk);
  dff _55956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _24252_, clk);
  dff _55957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _24466_, clk);
  dff _55958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _02342_, clk);
  dff _55959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _05861_, clk);
  dff _55960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _27244_, clk);
  dff _55961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _22944_, clk);
  dff _55962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _10686_, clk);
  dff _55963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _22667_, clk);
  dff _55964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _27245_, clk);
  dff _55965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _10713_, clk);
  dff _55966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _26075_, clk);
  dff _55967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _26030_, clk);
  dff _55968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _27161_, clk);
  dff _55969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _26046_, clk);
  dff _55970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _23326_, clk);
  dff _55971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _27162_, clk);
  dff _55972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _12268_, clk);
  dff _55973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _12251_, clk);
  dff _55974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _02457_, clk);
  dff _55975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _12065_, clk);
  dff _55976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _02454_, clk);
  dff _55977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _27159_, clk);
  dff _55978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _27160_, clk);
  dff _55979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _02721_, clk);
  dff _55980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _10936_, clk);
  dff _55981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _10910_, clk);
  dff _55982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _06923_, clk);
  dff _55983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _02466_, clk);
  dff _55984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _07214_, clk);
  dff _55985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _02464_, clk);
  dff _55986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _05330_, clk);
  dff _55987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _27157_, clk);
  dff _55988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _11920_, clk);
  dff _55989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _27158_, clk);
  dff _55990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _22664_, clk);
  dff _55991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _22662_, clk);
  dff _55992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _02477_, clk);
  dff _55993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _22661_, clk);
  dff _55994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _27151_, clk);
  dff _55995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _27152_, clk);
  dff _55996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _27153_, clk);
  dff _55997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _02725_, clk);
  dff _55998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _27147_, clk);
  dff _55999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _22669_, clk);
  dff _56000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _27148_, clk);
  dff _56001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _02487_, clk);
  dff _56002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _27149_, clk);
  dff _56003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _02482_, clk);
  dff _56004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _22666_, clk);
  dff _56005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _27150_, clk);
  dff _56006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _27144_, clk);
  dff _56007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _27145_, clk);
  dff _56008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _22678_, clk);
  dff _56009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _02496_, clk);
  dff _56010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _22672_, clk);
  dff _56011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _02493_, clk);
  dff _56012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _22671_, clk);
  dff _56013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _27146_, clk);
  dff _56014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _27142_, clk);
  dff _56015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _02736_, clk);
  dff _56016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _22723_, clk);
  dff _56017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _22686_, clk);
  dff _56018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _02510_, clk);
  dff _56019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _22685_, clk);
  dff _56020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _02506_, clk);
  dff _56021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _27143_, clk);
  dff _56022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _25079_, clk);
  dff _56023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _27140_, clk);
  dff _56024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _22929_, clk);
  dff _56025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _02529_, clk);
  dff _56026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _22915_, clk);
  dff _56027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _27141_, clk);
  dff _56028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _22860_, clk);
  dff _56029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _22739_, clk);
  dff _56030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _09328_, clk);
  dff _56031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _27137_, clk);
  dff _56032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _02747_, clk);
  dff _56033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _27138_, clk);
  dff _56034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _02538_, clk);
  dff _56035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _25774_, clk);
  dff _56036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _27139_, clk);
  dff _56037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _25762_, clk);
  dff _56038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _27133_, clk);
  dff _56039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _10690_, clk);
  dff _56040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _27134_, clk);
  dff _56041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _12342_, clk);
  dff _56042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _27135_, clk);
  dff _56043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _00019_, clk);
  dff _56044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _27136_, clk);
  dff _56045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _07444_, clk);
  dff _56046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _00994_, clk);
  dff _56047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _10681_, clk);
  dff _56048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _01254_, clk);
  dff _56049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _01235_, clk);
  dff _56050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _10675_, clk);
  dff _56051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _07540_, clk);
  dff _56052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _19907_, clk);
  dff _56053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _06071_, clk);
  dff _56054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _02547_, clk);
  dff _56055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _26621_, clk);
  dff _56056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _27129_, clk);
  dff _56057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _26604_, clk);
  dff _56058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _27130_, clk);
  dff _56059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _02741_, clk);
  dff _56060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _27131_, clk);
  dff _56061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _27132_, clk);
  dff _56062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _00007_, clk);
  dff _56063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _02559_, clk);
  dff _56064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _26785_, clk);
  dff _56065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _27125_, clk);
  dff _56066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _27126_, clk);
  dff _56067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _27127_, clk);
  dff _56068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _26746_, clk);
  dff _56069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _27128_, clk);
  dff _56070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _05450_, clk);
  dff _56071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _05383_, clk);
  dff _56072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _10609_, clk);
  dff _56073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _03511_, clk);
  dff _56074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _03297_, clk);
  dff _56075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _03262_, clk);
  dff _56076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _04262_, clk);
  dff _56077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _27242_, clk);
  dff _56078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _07370_, clk);
  dff _56079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _01407_, clk);
  dff _56080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _01392_, clk);
  dff _56081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _10658_, clk);
  dff _56082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _02099_, clk);
  dff _56083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _01495_, clk);
  dff _56084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _10650_, clk);
  dff _56085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _00985_, clk);
  dff _56086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _02575_, clk);
  dff _56087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _00515_, clk);
  dff _56088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _27123_, clk);
  dff _56089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _11519_, clk);
  dff _56090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _00087_, clk);
  dff _56091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _02567_, clk);
  dff _56092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _27124_, clk);
  dff _56093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _00032_, clk);
  dff _56094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _27118_, clk);
  dff _56095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _27119_, clk);
  dff _56096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _05764_, clk);
  dff _56097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _27120_, clk);
  dff _56098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _04562_, clk);
  dff _56099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _08410_, clk);
  dff _56100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _02579_, clk);
  dff _56101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _27121_, clk);
  dff _56102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _27117_, clk);
  dff _56103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _04931_, clk);
  dff _56104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _24445_, clk);
  dff _56105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _04934_, clk);
  dff _56106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _05168_, clk);
  dff _56107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _24477_, clk);
  dff _56108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _24488_, clk);
  dff _56109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _05052_, clk);
  dff _56110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _07544_, clk);
  dff _56111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _09691_, clk);
  dff _56112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _09688_, clk);
  dff _56113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _10589_, clk);
  dff _56114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _09721_, clk);
  dff _56115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _07391_, clk);
  dff _56116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _05783_, clk);
  dff _56117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _05703_, clk);
  dff _56118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _06787_, clk);
  dff _56119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _07103_, clk);
  dff _56120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _27241_, clk);
  dff _56121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _07870_, clk);
  dff _56122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _07961_, clk);
  dff _56123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _04889_, clk);
  dff _56124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _04839_, clk);
  dff _56125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _04811_, clk);
  dff _56126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _27234_, clk);
  dff _56127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _12140_, clk);
  dff _56128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _12154_, clk);
  dff _56129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _12142_, clk);
  dff _56130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _07403_, clk);
  dff _56131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _27235_, clk);
  dff _56132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _10958_, clk);
  dff _56133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _10941_, clk);
  dff _56134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _11228_, clk);
  dff _56135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _27236_, clk);
  dff _56136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _10513_, clk);
  dff _56137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _07546_, clk);
  dff _56138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _10833_, clk);
  dff _56139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _27237_, clk);
  dff _56140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _27238_, clk);
  dff _56141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _27239_, clk);
  dff _56142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _25887_, clk);
  dff _56143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _25904_, clk);
  dff _56144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _25889_, clk);
  dff _56145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _27080_, clk);
  dff _56146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _25949_, clk);
  dff _56147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _11553_, clk);
  dff _56148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _25731_, clk);
  dff _56149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _25742_, clk);
  dff _56150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _12420_, clk);
  dff _56151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _00074_, clk);
  dff _56152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _22663_, clk);
  dff _56153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _27232_, clk);
  dff _56154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _22628_, clk);
  dff _56155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _22635_, clk);
  dff _56156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _07414_, clk);
  dff _56157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _27233_, clk);
  dff _56158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _11463_, clk);
  dff _56159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _04174_, clk);
  dff _56160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _11462_, clk);
  dff _56161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _04075_, clk);
  dff _56162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _04101_, clk);
  dff _56163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _11466_, clk);
  dff _56164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _03992_, clk);
  dff _56165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _26894_, clk);
  dff _56166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _25399_, clk);
  dff _56167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _25389_, clk);
  dff _56168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _25439_, clk);
  dff _56169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _27213_, clk);
  dff _56170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _25427_, clk);
  dff _56171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _11300_, clk);
  dff _56172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _25317_, clk);
  dff _56173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _25304_, clk);
  dff _56174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _25537_, clk);
  dff _56175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _25530_, clk);
  dff _56176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _25570_, clk);
  dff _56177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _25559_, clk);
  dff _56178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _11446_, clk);
  dff _56179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _25468_, clk);
  dff _56180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _25464_, clk);
  dff _56181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _25498_, clk);
  dff _56182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _25857_, clk);
  dff _56183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _11563_, clk);
  dff _56184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _11390_, clk);
  dff _56185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _25667_, clk);
  dff _56186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _25653_, clk);
  dff _56187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _11592_, clk);
  dff _56188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _25702_, clk);
  dff _56189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _27189_, clk);
  dff _56190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _27258_, clk);
  dff _56191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _11630_, clk);
  dff _56192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _24435_, clk);
  dff _56193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _27259_, clk);
  dff _56194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _27260_, clk);
  dff _56195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _24338_, clk);
  dff _56196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _24335_, clk);
  dff _56197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _24356_, clk);
  dff _56198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _24463_, clk);
  dff _56199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _24456_, clk);
  dff _56200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _27243_, clk);
  dff _56201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _24524_, clk);
  dff _56202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _24506_, clk);
  dff _56203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _24501_, clk);
  dff _56204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _11298_, clk);
  dff _56205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _24366_, clk);
  dff _56206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _25348_, clk);
  dff _56207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _11603_, clk);
  dff _56208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _25239_, clk);
  dff _56209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _25237_, clk);
  dff _56210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _25031_, clk);
  dff _56211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _11611_, clk);
  dff _56212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _27228_, clk);
  dff _56213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _25265_, clk);
  dff _56214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _11632_, clk);
  dff _56215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _27289_, clk);
  dff _56216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _27290_, clk);
  dff _56217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _24211_, clk);
  dff _56218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _24202_, clk);
  dff _56219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _24288_, clk);
  dff _56220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _24285_, clk);
  dff _56221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _24256_, clk);
  dff _56222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _04958_, clk);
  dff _56223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _04962_, clk);
  dff _56224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _05005_, clk);
  dff _56225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _04954_, clk);
  dff _56226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _24213_, clk);
  dff _56227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _04863_, clk);
  dff _56228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _24215_, clk);
  dff _56229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _24183_, clk);
  dff _56230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _03336_, clk);
  dff _56231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _04487_, clk);
  dff _56232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _03509_, clk);
  dff _56233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _05113_, clk);
  dff _56234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _27116_, clk);
  dff _56235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _05089_, clk);
  dff _56236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _04873_, clk);
  dff _56237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _04914_, clk);
  dff _56238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _03352_, clk);
  dff _56239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _04381_, clk);
  dff _56240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _27114_, clk);
  dff _56241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _04424_, clk);
  dff _56242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _03345_, clk);
  dff _56243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _27115_, clk);
  dff _56244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _04455_, clk);
  dff _56245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _03339_, clk);
  dff _56246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _04310_, clk);
  dff _56247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _27111_, clk);
  dff _56248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _04316_, clk);
  dff _56249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _03519_, clk);
  dff _56250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _04324_, clk);
  dff _56251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _27112_, clk);
  dff _56252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _27113_, clk);
  dff _56253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _03598_, clk);
  dff _56254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _03389_, clk);
  dff _56255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _27109_, clk);
  dff _56256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _03533_, clk);
  dff _56257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _04254_, clk);
  dff _56258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _04271_, clk);
  dff _56259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _03529_, clk);
  dff _56260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _04282_, clk);
  dff _56261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _27110_, clk);
  dff _56262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _27108_, clk);
  dff _56263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _04171_, clk);
  dff _56264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _04189_, clk);
  dff _56265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _03401_, clk);
  dff _56266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _03605_, clk);
  dff _56267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _04194_, clk);
  dff _56268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _04208_, clk);
  dff _56269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _03399_, clk);
  dff _56270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _27106_, clk);
  dff _56271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _04087_, clk);
  dff _56272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _04112_, clk);
  dff _56273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _03427_, clk);
  dff _56274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _04116_, clk);
  dff _56275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _03539_, clk);
  dff _56276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _27107_, clk);
  dff _56277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _04162_, clk);
  dff _56278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _03749_, clk);
  dff _56279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _27101_, clk);
  dff _56280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _27102_, clk);
  dff _56281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _27103_, clk);
  dff _56282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _27104_, clk);
  dff _56283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _04040_, clk);
  dff _56284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _04068_, clk);
  dff _56285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _27105_, clk);
  dff _56286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _03673_, clk);
  dff _56287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _27098_, clk);
  dff _56288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _03671_, clk);
  dff _56289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _03507_, clk);
  dff _56290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _03695_, clk);
  dff _56291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _03718_, clk);
  dff _56292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _03498_, clk);
  dff _56293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _03726_, clk);
  dff _56294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _03921_, clk);
  dff _56295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _03948_, clk);
  dff _56296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _03560_, clk);
  dff _56297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _27097_, clk);
  dff _56298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _03969_, clk);
  dff _56299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _03989_, clk);
  dff _56300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _04007_, clk);
  dff _56301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _03456_, clk);
  dff _56302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _03477_, clk);
  dff _56303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _03848_, clk);
  dff _56304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _03475_, clk);
  dff _56305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _03854_, clk);
  dff _56306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _03627_, clk);
  dff _56307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _03864_, clk);
  dff _56308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _03918_, clk);
  dff _56309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _03467_, clk);
  dff _56310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _03761_, clk);
  dff _56311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _03486_, clk);
  dff _56312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _03768_, clk);
  dff _56313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _03573_, clk);
  dff _56314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _03780_, clk);
  dff _56315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _03800_, clk);
  dff _56316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _03817_, clk);
  dff _56317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _03483_, clk);
  dff _56318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _04968_, clk);
  dff _56319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _25245_, clk);
  dff _56320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _25087_, clk);
  dff _56321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _24958_, clk);
  dff _56322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _27095_, clk);
  dff _56323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _25282_, clk);
  dff _56324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _25273_, clk);
  dff _56325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _27096_, clk);
  dff _56326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _25437_, clk);
  dff _56327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _04960_, clk);
  dff _56328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _25324_, clk);
  dff _56329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _25337_, clk);
  dff _56330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _25326_, clk);
  dff _56331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _04972_, clk);
  dff _56332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _25373_, clk);
  dff _56333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _27094_, clk);
  dff _56334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _04883_, clk);
  dff _56335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _24135_, clk);
  dff _56336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _24128_, clk);
  dff _56337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _24103_, clk);
  dff _56338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _24316_, clk);
  dff _56339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _24282_, clk);
  dff _56340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _24242_, clk);
  dff _56341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _27093_, clk);
  dff _56342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _25871_, clk);
  dff _56343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _25853_, clk);
  dff _56344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _25906_, clk);
  dff _56345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _24329_, clk);
  dff _56346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _24344_, clk);
  dff _56347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _04906_, clk);
  dff _56348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _24359_, clk);
  dff _56349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _24370_, clk);
  dff _56350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _25471_, clk);
  dff _56351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _05154_, clk);
  dff _56352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _27091_, clk);
  dff _56353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _25525_, clk);
  dff _56354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _27092_, clk);
  dff _56355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _25733_, clk);
  dff _56356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _25725_, clk);
  dff _56357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _25717_, clk);
  dff _56358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _23180_, clk);
  dff _56359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _02770_, clk);
  dff _56360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _25562_, clk);
  dff _56361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _25555_, clk);
  dff _56362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _25676_, clk);
  dff _56363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _25671_, clk);
  dff _56364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _25641_, clk);
  dff _56365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _25476_, clk);
  dff _56366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _01070_, clk);
  dff _56367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _01307_, clk);
  dff _56368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _01379_, clk);
  dff _56369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _04473_, clk);
  dff _56370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _22684_, clk);
  dff _56371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _09347_, clk);
  dff _56372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _27089_, clk);
  dff _56373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _24235_, clk);
  dff _56374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _04445_, clk);
  dff _56375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _02165_, clk);
  dff _56376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _02081_, clk);
  dff _56377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _27088_, clk);
  dff _56378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _03766_, clk);
  dff _56379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _03648_, clk);
  dff _56380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _02773_, clk);
  dff _56381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _01196_, clk);
  dff _56382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _04432_, clk);
  dff _56383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _09686_, clk);
  dff _56384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _09103_, clk);
  dff _56385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _02781_, clk);
  dff _56386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _05027_, clk);
  dff _56387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _04850_, clk);
  dff _56388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _04776_, clk);
  dff _56389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _05648_, clk);
  dff _56390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _10154_, clk);
  dff _56391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _04417_, clk);
  dff _56392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _10622_, clk);
  dff _56393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _10668_, clk);
  dff _56394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _04408_, clk);
  dff _56395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _07449_, clk);
  dff _56396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _07100_, clk);
  dff _56397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _05935_, clk);
  dff _56398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _11916_, clk);
  dff _56399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _04369_, clk);
  dff _56400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _27085_, clk);
  dff _56401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _27086_, clk);
  dff _56402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _27087_, clk);
  dff _56403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _04398_, clk);
  dff _56404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _10886_, clk);
  dff _56405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _10891_, clk);
  dff _56406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _22627_, clk);
  dff _56407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _22665_, clk);
  dff _56408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _04354_, clk);
  dff _56409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _03116_, clk);
  dff _56410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _11133_, clk);
  dff _56411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _27084_, clk);
  dff _56412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _11076_, clk);
  dff _56413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _11925_, clk);
  dff _56414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _24363_, clk);
  dff _56415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _22720_, clk);
  dff _56416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _22714_, clk);
  dff _56417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _04346_, clk);
  dff _56418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _22680_, clk);
  dff _56419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _12416_, clk);
  dff _56420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _12353_, clk);
  dff _56421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _04359_, clk);
  dff _56422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _25379_, clk);
  dff _56423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _04321_, clk);
  dff _56424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _01500_, clk);
  dff _56425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _27083_, clk);
  dff _56426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _04318_, clk);
  dff _56427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _03117_, clk);
  dff _56428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _25095_, clk);
  dff _56429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _13109_, clk);
  dff _56430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _01925_, clk);
  dff _56431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _02151_, clk);
  dff _56432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _02042_, clk);
  dff _56433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _04313_, clk);
  dff _56434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _04490_, clk);
  dff _56435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _04422_, clk);
  dff _56436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _03609_, clk);
  dff _56437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _02797_, clk);
  dff _56438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _08865_, clk);
  dff _56439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _27081_, clk);
  dff _56440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _05217_, clk);
  dff _56441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _04870_, clk);
  dff _56442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _04307_, clk);
  dff _56443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _27082_, clk);
  dff _56444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _07123_, clk);
  dff _56445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _04299_, clk);
  dff _56446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _09096_, clk);
  dff _56447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _09317_, clk);
  dff _56448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _27078_, clk);
  dff _56449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _04269_, clk);
  dff _56450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _08782_, clk);
  dff _56451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _27079_, clk);
  dff _56452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _04294_, clk);
  dff _56453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _08873_, clk);
  dff _56454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _09416_, clk);
  dff _56455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _09402_, clk);
  dff _56456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _09391_, clk);
  dff _56457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _10048_, clk);
  dff _56458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _09743_, clk);
  dff _56459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _09544_, clk);
  dff _56460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _02808_, clk);
  dff _56461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _09270_, clk);
  dff _56462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _11927_, clk);
  dff _56463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _27076_, clk);
  dff _56464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _27077_, clk);
  dff _56465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _10736_, clk);
  dff _56466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _10630_, clk);
  dff _56467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _10918_, clk);
  dff _56468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _10925_, clk);
  dff _56469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _02828_, clk);
  dff _56470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _08767_, clk);
  dff _56471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _05290_, clk);
  dff _56472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _04218_, clk);
  dff _56473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _22687_, clk);
  dff _56474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _04205_, clk);
  dff _56475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _03130_, clk);
  dff _56476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _11614_, clk);
  dff _56477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _11596_, clk);
  dff _56478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _03268_, clk);
  dff _56479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _02052_, clk);
  dff _56480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _02261_, clk);
  dff _56481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _02128_, clk);
  dff _56482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _04200_, clk);
  dff _56483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _04515_, clk);
  dff _56484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _04731_, clk);
  dff _56485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _04600_, clk);
  dff _56486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _04177_, clk);
  dff _56487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _06555_, clk);
  dff _56488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _07427_, clk);
  dff _56489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _06604_, clk);
  dff _56490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _04191_, clk);
  dff _56491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _10844_, clk);
  dff _56492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _09613_, clk);
  dff _56493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _04187_, clk);
  dff _56494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _08667_, clk);
  dff _56495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _02864_, clk);
  dff _56496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _27074_, clk);
  dff _56497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _01799_, clk);
  dff _56498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _23384_, clk);
  dff _56499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _27075_, clk);
  dff _56500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _03079_, clk);
  dff _56501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _11528_, clk);
  dff _56502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _26771_, clk);
  dff _56503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _00044_, clk);
  dff _56504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _00079_, clk);
  dff _56505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _27073_, clk);
  dff _56506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _08738_, clk);
  dff _56507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _04168_, clk);
  dff _56508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _08650_, clk);
  dff _56509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _08655_, clk);
  dff _56510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _27070_, clk);
  dff _56511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _03932_, clk);
  dff _56512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _04198_, clk);
  dff _56513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _27071_, clk);
  dff _56514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _03160_, clk);
  dff _56515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _27072_, clk);
  dff _56516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _08597_, clk);
  dff _56517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _08602_, clk);
  dff _56518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _00172_, clk);
  dff _56519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _27067_, clk);
  dff _56520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _26774_, clk);
  dff _56521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _27068_, clk);
  dff _56522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _27069_, clk);
  dff _56523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _04107_, clk);
  dff _56524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _03426_, clk);
  dff _56525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _11001_, clk);
  dff _56526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _06349_, clk);
  dff _56527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _12202_, clk);
  dff _56528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _07226_, clk);
  dff _56529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _22659_, clk);
  dff _56530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _04097_, clk);
  dff _56531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _18267_, clk);
  dff _56532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _06239_, clk);
  dff _56533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _04089_, clk);
  dff _56534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _04072_, clk);
  dff _56535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _08817_, clk);
  dff _56536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _04050_, clk);
  dff _56537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _27063_, clk);
  dff _56538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _25114_, clk);
  dff _56539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _23315_, clk);
  dff _56540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _27064_, clk);
  dff _56541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _27065_, clk);
  dff _56542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _04026_, clk);
  dff _56543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _27057_, clk);
  dff _56544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _27058_, clk);
  dff _56545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _27059_, clk);
  dff _56546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _27060_, clk);
  dff _56547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _27061_, clk);
  dff _56548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _27062_, clk);
  dff _56549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _18155_, clk);
  dff _56550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _27056_, clk);
  dff _56551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _23993_, clk);
  dff _56552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _25749_, clk);
  dff _56553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _25595_, clk);
  dff _56554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _11326_, clk);
  dff _56555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _11496_, clk);
  dff _56556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _04037_, clk);
  dff _56557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _09147_, clk);
  dff _56558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _27053_, clk);
  dff _56559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _23200_, clk);
  dff _56560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _27054_, clk);
  dff _56561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _03099_, clk);
  dff _56562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _27055_, clk);
  dff _56563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _03753_, clk);
  dff _56564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _03741_, clk);
  dff _56565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _03240_, clk);
  dff _56566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _08023_, clk);
  dff _56567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _09950_, clk);
  dff _56568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _09966_, clk);
  dff _56569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _09974_, clk);
  dff _56570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _27285_, clk);
  dff _56571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _10008_, clk);
  dff _56572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _08020_, clk);
  dff _56573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _27286_, clk);
  dff _56574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _25624_, clk);
  dff _56575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _25474_, clk);
  dff _56576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _25419_, clk);
  dff _56577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _10968_, clk);
  dff _56578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _27284_, clk);
  dff _56579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _09886_, clk);
  dff _56580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _09908_, clk);
  dff _56581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _08238_, clk);
  dff _56582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _25843_, clk);
  dff _56583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _27280_, clk);
  dff _56584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _27281_, clk);
  dff _56585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _27282_, clk);
  dff _56586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _27283_, clk);
  dff _56587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _24901_, clk);
  dff _56588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _24796_, clk);
  dff _56589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _24683_, clk);
  dff _56590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _00972_, clk);
  dff _56591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _05091_, clk);
  dff _56592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _10950_, clk);
  dff _56593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _22622_, clk);
  dff _56594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _27278_, clk);
  dff _56595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _27279_, clk);
  dff _56596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _25824_, clk);
  dff _56597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _25943_, clk);
  dff _56598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _10948_, clk);
  dff _56599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _03395_, clk);
  dff _56600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _06732_, clk);
  dff _56601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _04137_, clk);
  dff _56602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _10938_, clk);
  dff _56603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _22614_, clk);
  dff _56604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _25847_, clk);
  dff _56605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _10955_, clk);
  dff _56606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _27274_, clk);
  dff _56607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _27275_, clk);
  dff _56608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _27276_, clk);
  dff _56609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _27277_, clk);
  dff _56610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _11036_, clk);
  dff _56611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _22689_, clk);
  dff _56612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _11173_, clk);
  dff _56613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _09287_, clk);
  dff _56614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _27268_, clk);
  dff _56615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _27269_, clk);
  dff _56616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _27270_, clk);
  dff _56617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _27271_, clk);
  dff _56618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _27272_, clk);
  dff _56619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _27273_, clk);
  dff _56620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _11048_, clk);
  dff _56621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _11017_, clk);
  dff _56622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _10838_, clk);
  dff _56623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _07338_, clk);
  dff _56624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _07626_, clk);
  dff _56625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _27263_, clk);
  dff _56626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _27264_, clk);
  dff _56627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _27265_, clk);
  dff _56628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _27266_, clk);
  dff _56629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _27267_, clk);
  dff _56630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _10901_, clk);
  dff _56631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _10999_, clk);
  dff _56632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _11014_, clk);
  dff _56633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _27261_, clk);
  dff _56634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _03548_, clk);
  dff _56635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _27262_, clk);
  dff _56636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _10820_, clk);
  dff _56637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _10866_, clk);
  dff _56638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _07346_, clk);
  dff _56639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _27257_, clk);
  dff _56640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _11071_, clk);
  dff _56641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _11156_, clk);
  dff _56642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _11144_, clk);
  dff _56643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _11124_, clk);
  dff _56644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _07344_, clk);
  dff _56645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _10897_, clk);
  dff _56646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _11752_, clk);
  dff _56647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _11694_, clk);
  dff _56648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _07353_, clk);
  dff _56649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _27256_, clk);
  dff _56650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _11242_, clk);
  dff _56651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _11220_, clk);
  dff _56652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _11369_, clk);
  dff _56653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _11303_, clk);
  dff _56654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _27253_, clk);
  dff _56655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _09331_, clk);
  dff _56656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _09427_, clk);
  dff _56657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _27254_, clk);
  dff _56658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _11601_, clk);
  dff _56659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _27255_, clk);
  dff _56660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _11452_, clk);
  dff _56661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _11425_, clk);
  dff _56662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _09666_, clk);
  dff _56663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _09662_, clk);
  dff _56664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _09649_, clk);
  dff _56665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _27251_, clk);
  dff _56666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _12148_, clk);
  dff _56667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _23365_, clk);
  dff _56668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _07355_, clk);
  dff _56669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _27252_, clk);
  dff _56670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _27249_, clk);
  dff _56671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _27250_, clk);
  dff _56672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _08400_, clk);
  dff _56673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _08408_, clk);
  dff _56674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _08949_, clk);
  dff _56675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _26817_, clk);
  dff _56676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _00022_, clk);
  dff _56677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _00082_, clk);
  dff _56678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _27248_, clk);
  dff _56679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _07360_, clk);
  dff _56680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _26728_, clk);
  dff _56681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _26685_, clk);
  dff _56682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _26725_, clk);
  dff _56683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _25076_, clk);
  dff _56684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _25082_, clk);
  dff _56685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _25747_, clk);
  dff _56686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _22623_, clk);
  dff _56687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _10090_, clk);
  dff _56688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _11550_, clk);
  dff _56689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _11594_, clk);
  dff _56690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _27217_, clk);
  dff _56691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _11658_, clk);
  dff _56692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _11902_, clk);
  dff _56693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _10111_, clk);
  dff _56694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _11213_, clk);
  dff _56695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _05882_, clk);
  dff _56696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _05940_, clk);
  dff _56697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _11167_, clk);
  dff _56698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _11234_, clk);
  dff _56699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _07386_, clk);
  dff _56700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _07614_, clk);
  dff _56701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _27195_, clk);
  dff _56702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _27214_, clk);
  dff _56703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _23135_, clk);
  dff _56704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _00674_, clk);
  dff _56705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _27215_, clk);
  dff _56706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _07565_, clk);
  dff _56707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _27216_, clk);
  dff _56708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _26078_, clk);
  dff _56709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _10097_, clk);
  dff _56710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _07199_, clk);
  dff _56711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _11126_, clk);
  dff _56712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _07223_, clk);
  dff _56713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _11200_, clk);
  dff _56714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _07276_, clk);
  dff _56715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _07366_, clk);
  dff _56716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _05608_, clk);
  dff _56717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _11172_, clk);
  dff _56718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _10059_, clk);
  dff _56719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _07580_, clk);
  dff _56720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _03443_, clk);
  dff _56721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _27212_, clk);
  dff _56722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _04814_, clk);
  dff _56723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _07462_, clk);
  dff _56724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _04780_, clk);
  dff _56725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _22645_, clk);
  dff _56726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _11204_, clk);
  dff _56727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _06772_, clk);
  dff _56728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _11135_, clk);
  dff _56729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _06814_, clk);
  dff _56730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _11202_, clk);
  dff _56731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _06894_, clk);
  dff _56732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _07047_, clk);
  dff _56733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _11128_, clk);
  dff _56734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _07898_, clk);
  dff _56735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _10818_, clk);
  dff _56736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _10928_, clk);
  dff _56737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _23110_, clk);
  dff _56738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _10043_, clk);
  dff _56739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _06806_, clk);
  dff _56740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _27211_, clk);
  dff _56741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _09412_, clk);
  dff _56742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _06304_, clk);
  dff _56743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _11146_, clk);
  dff _56744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _11232_, clk);
  dff _56745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _06382_, clk);
  dff _56746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _06622_, clk);
  dff _56747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _27193_, clk);
  dff _56748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _27194_, clk);
  dff _56749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _06722_, clk);
  dff _56750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _12422_, clk);
  dff _56751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _04624_, clk);
  dff _56752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _04621_, clk);
  dff _56753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _12424_, clk);
  dff _56754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _06025_, clk);
  dff _56755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _06076_, clk);
  dff _56756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _27192_, clk);
  dff _56757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _06235_, clk);
  dff _56758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _12399_, clk);
  dff _56759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _26661_, clk);
  dff _56760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _04365_, clk);
  dff _56761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _12274_, clk);
  dff _56762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _04371_, clk);
  dff _56763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _04588_, clk);
  dff _56764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _12332_, clk);
  dff _56765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _04591_, clk);
  dff _56766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _27190_, clk);
  dff _56767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _27191_, clk);
  dff _56768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _04655_, clk);
  dff _56769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _12397_, clk);
  dff _56770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _04728_, clk);
  dff _56771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _04720_, clk);
  dff _56772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _04713_, clk);
  dff _56773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _12357_, clk);
  dff _56774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _04857_, clk);
  dff _56775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _04788_, clk);
  dff _56776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _04784_, clk);
  dff _56777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _04771_, clk);
  dff _56778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _27188_, clk);
  dff _56779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _04836_, clk);
  dff _56780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _04834_, clk);
  dff _56781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _04822_, clk);
  dff _56782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _04296_, clk);
  dff _56783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _04284_, clk);
  dff _56784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _04415_, clk);
  dff _56785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _04411_, clk);
  dff _56786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _04391_, clk);
  dff _56787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _27186_, clk);
  dff _56788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _04351_, clk);
  dff _56789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _27187_, clk);
  dff _56790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _27185_, clk);
  dff _56791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _04453_, clk);
  dff _56792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _04457_, clk);
  dff _56793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _12293_, clk);
  dff _56794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _04509_, clk);
  dff _56795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _04546_, clk);
  dff _56796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _04511_, clk);
  dff _56797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _12280_, clk);
  dff _56798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _27182_, clk);
  dff _56799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _27183_, clk);
  dff _56800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _27184_, clk);
  dff _56801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _05143_, clk);
  dff _56802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _05206_, clk);
  dff _56803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _05187_, clk);
  dff _56804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _09513_, clk);
  dff _56805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _04618_, clk);
  dff _56806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _05064_, clk);
  dff _56807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _27179_, clk);
  dff _56808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _04922_, clk);
  dff _56809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _04919_, clk);
  dff _56810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _04911_, clk);
  dff _56811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _27180_, clk);
  dff _56812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _04963_, clk);
  dff _56813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _27181_, clk);
  dff _56814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _22658_, clk);
  dff _56815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _27019_, clk);
  dff _56816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _22674_, clk);
  dff _56817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _22673_, clk);
  dff _56818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _11285_, clk);
  dff _56819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _22651_, clk);
  dff _56820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _27020_, clk);
  dff _56821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _27021_, clk);
  dff _56822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _27099_, clk);
  dff _56823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _11759_, clk);
  dff _56824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _18441_, clk);
  dff _56825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _18950_, clk);
  dff _56826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _11757_, clk);
  dff _56827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _11375_, clk);
  dff _56828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _12748_, clk);
  dff _56829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _27100_, clk);
  dff _56830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _10953_, clk);
  dff _56831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _10942_, clk);
  dff _56832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _10984_, clk);
  dff _56833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _10995_, clk);
  dff _56834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _11005_, clk);
  dff _56835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _10976_, clk);
  dff _56836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _27310_, clk);
  dff _56837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _09884_, clk);
  dff _56838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _03123_, clk);
  dff _56839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _27023_, clk);
  dff _56840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _05607_, clk);
  dff _56841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _03125_, clk);
  dff _56842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _03154_, clk);
  dff _56843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _05189_, clk);
  dff _56844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _03163_, clk);
  dff _56845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _03179_, clk);
  dff _56846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _05466_, clk);
  dff _56847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _25452_, clk);
  dff _56848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _22879_, clk);
  dff _56849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _23021_, clk);
  dff _56850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _22959_, clk);
  dff _56851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _03095_, clk);
  dff _56852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _27024_, clk);
  dff _56853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _22798_, clk);
  dff _56854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _06948_, clk);
  dff _56855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _06955_, clk);
  dff _56856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _27008_, clk);
  dff _56857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _03418_, clk);
  dff _56858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _26029_, clk);
  dff _56859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _05445_, clk);
  dff _56860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _26033_, clk);
  dff _56861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _27009_, clk);
  dff _56862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _10923_, clk);
  dff _56863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _06340_, clk);
  dff _56864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _06086_, clk);
  dff _56865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _10431_, clk);
  dff _56866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _10434_, clk);
  dff _56867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _06346_, clk);
  dff _56868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _10739_, clk);
  dff _56869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _26959_, clk);
  dff _56870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _26960_, clk);
  dff _56871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _10151_, clk);
  dff _56872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _06350_, clk);
  dff _56873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _26961_, clk);
  dff _56874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _10194_, clk);
  dff _56875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _05917_, clk);
  dff _56876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06179_, clk);
  dff _56877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _12261_, clk);
  dff _56878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _11021_, clk);
  dff _56879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _06336_, clk);
  dff _56880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _26957_, clk);
  dff _56881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _05932_, clk);
  dff _56882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _10828_, clk);
  dff _56883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _10864_, clk);
  dff _56884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _10831_, clk);
  dff _56885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _26958_, clk);
  dff _56886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _26934_, clk);
  dff _56887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _10506_, clk);
  dff _56888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _07043_, clk);
  dff _56889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _10539_, clk);
  dff _56890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _07197_, clk);
  dff _56891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _10569_, clk);
  dff _56892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _26935_, clk);
  dff _56893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _07037_, clk);
  dff _56894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _07965_, clk);
  dff _56895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _08812_, clk);
  dff _56896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _11043_, clk);
  dff _56897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _27309_, clk);
  dff _56898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _11023_, clk);
  dff _56899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _11039_, clk);
  dff _56900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _11024_, clk);
  dff _56901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _10946_, clk);
  dff _56902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _10881_, clk);
  dff _56903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _27240_, clk);
  dff _56904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _10883_, clk);
  dff _56905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _07397_, clk);
  dff _56906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _10599_, clk);
  dff _56907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _10574_, clk);
  dff _56908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _10716_, clk);
  dff _56909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _10711_, clk);
  dff _56910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _27230_, clk);
  dff _56911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _25352_, clk);
  dff _56912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _06338_, clk);
  dff _56913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _03576_, clk);
  dff _56914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _14268_, clk);
  dff _56915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _27231_, clk);
  dff _56916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _08017_, clk);
  dff _56917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _04393_, clk);
  dff _56918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _01504_, clk);
  dff _56919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _01404_, clk);
  dff _56920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _23102_, clk);
  dff _56921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _22939_, clk);
  dff _56922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _10366_, clk);
  dff _56923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _25037_, clk);
  dff _56924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _25170_, clk);
  dff _56925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _27229_, clk);
  dff _56926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _27224_, clk);
  dff _56927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _09017_, clk);
  dff _56928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _09014_, clk);
  dff _56929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _10181_, clk);
  dff _56930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _07180_, clk);
  dff _56931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _27225_, clk);
  dff _56932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _10190_, clk);
  dff _56933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _07513_, clk);
  dff _56934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _02030_, clk);
  dff _56935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _10244_, clk);
  dff _56936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _02327_, clk);
  dff _56937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _03156_, clk);
  dff _56938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _10214_, clk);
  dff _56939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _26052_, clk);
  dff _56940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _00657_, clk);
  dff _56941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _00289_, clk);
  dff _56942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _27226_, clk);
  dff _56943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _04504_, clk);
  dff _56944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _04525_, clk);
  dff _56945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _04506_, clk);
  dff _56946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _05470_, clk);
  dff _56947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _05135_, clk);
  dff _56948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _10198_, clk);
  dff _56949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _27227_, clk);
  dff _56950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _23171_, clk);
  dff _56951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _27219_, clk);
  dff _56952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _24346_, clk);
  dff _56953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _25875_, clk);
  dff _56954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _25960_, clk);
  dff _56955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _09807_, clk);
  dff _56956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _27220_, clk);
  dff _56957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _09846_, clk);
  dff _56958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _27222_, clk);
  dff _56959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _09268_, clk);
  dff _56960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _09256_, clk);
  dff _56961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _10177_, clk);
  dff _56962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _27223_, clk);
  dff _56963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _09276_, clk);
  dff _56964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _07433_, clk);
  dff _56965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _08825_, clk);
  dff _56966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _06088_, clk);
  dff _56967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _06268_, clk);
  dff _56968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _01224_, clk);
  dff _56969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _07506_, clk);
  dff _56970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _07910_, clk);
  dff _56971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _09367_, clk);
  dff _56972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _09357_, clk);
  dff _56973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _27221_, clk);
  dff _56974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _10613_, clk);
  dff _56975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _10577_, clk);
  dff _56976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _10551_, clk);
  dff _56977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _09063_, clk);
  dff _56978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _09735_, clk);
  dff _56979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _09996_, clk);
  dff _56980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _09218_, clk);
  dff _56981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _06207_, clk);
  dff _56982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _18176_, clk);
  dff _56983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _07515_, clk);
  dff _56984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _10974_, clk);
  dff _56985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _12393_, clk);
  dff _56986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _09214_, clk);
  dff _56987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _01301_, clk);
  dff _56988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _09207_, clk);
  dff _56989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _07912_, clk);
  dff _56990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _19605_, clk);
  dff _56991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _27090_, clk);
  dff _56992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _19639_, clk);
  dff _56993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _21642_, clk);
  dff _56994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _21519_, clk);
  dff _56995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _21388_, clk);
  dff _56996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _11754_, clk);
  dff _56997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _17998_, clk);
  dff _56998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _11714_, clk);
  dff _56999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _22615_, clk);
  dff _57000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _22613_, clk);
  dff _57001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _22612_, clk);
  dff _57002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _22621_, clk);
  dff _57003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _22619_, clk);
  dff _57004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _22618_, clk);
  dff _57005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _11750_, clk);
  dff _57006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _22657_, clk);
  dff _57007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _22655_, clk);
  dff _57008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _11696_, clk);
  dff _57009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _27037_, clk);
  dff _57010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _22638_, clk);
  dff _57011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _22637_, clk);
  dff _57012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _27038_, clk);
  dff _57013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _22648_, clk);
  dff _57014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _22647_, clk);
  dff _57015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _11699_, clk);
  dff _57016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _11380_, clk);
  dff _57017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _11450_, clk);
  dff _57018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _27066_, clk);
  dff _57019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _22625_, clk);
  dff _57020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _22630_, clk);
  dff _57021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _22634_, clk);
  dff _57022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _27007_, clk);
  dff _57023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _11287_, clk);
  dff _57024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _11439_, clk);
  dff _57025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _22683_, clk);
  dff _57026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _22682_, clk);
  dff _57027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _11691_, clk);
  dff _57028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _22721_, clk);
  dff _57029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _22717_, clk);
  dff _57030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _03664_, clk);
  dff _57031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _03300_, clk);
  dff _57032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _03704_, clk);
  dff _57033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _23428_, clk);
  dff _57034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _03701_, clk);
  dff _57035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _23307_, clk);
  dff _57036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _27052_, clk);
  dff _57037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _23332_, clk);
  dff _57038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _26270_, clk);
  dff _57039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _26134_, clk);
  dff _57040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _27047_, clk);
  dff _57041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _27048_, clk);
  dff _57042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _27049_, clk);
  dff _57043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _04005_, clk);
  dff _57044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _03177_, clk);
  dff _57045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _23852_, clk);
  dff _57046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _23961_, clk);
  dff _57047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _03675_, clk);
  dff _57048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _27050_, clk);
  dff _57049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _27051_, clk);
  dff _57050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _03103_, clk);
  dff _57051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _24049_, clk);
  dff _57052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _24007_, clk);
  dff _57053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _24084_, clk);
  dff _57054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _27042_, clk);
  dff _57055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _03971_, clk);
  dff _57056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _27043_, clk);
  dff _57057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _27044_, clk);
  dff _57058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _03999_, clk);
  dff _57059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _27045_, clk);
  dff _57060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _27046_, clk);
  dff _57061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _03994_, clk);
  dff _57062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _27036_, clk);
  dff _57063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _12616_, clk);
  dff _57064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _12515_, clk);
  dff _57065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _03056_, clk);
  dff _57066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _10727_, clk);
  dff _57067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _10814_, clk);
  dff _57068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _11416_, clk);
  dff _57069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _03924_, clk);
  dff _57070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _27039_, clk);
  dff _57071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _03961_, clk);
  dff _57072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _06056_, clk);
  dff _57073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _06601_, clk);
  dff _57074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _03051_, clk);
  dff _57075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _27040_, clk);
  dff _57076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _27041_, clk);
  dff _57077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _03986_, clk);
  dff _57078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _07894_, clk);
  dff _57079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _08331_, clk);
  dff _57080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _08103_, clk);
  dff _57081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _10347_, clk);
  dff _57082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _10107_, clk);
  dff _57083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _10012_, clk);
  dff _57084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _03053_, clk);
  dff _57085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _05303_, clk);
  dff _57086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _27033_, clk);
  dff _57087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _03856_, clk);
  dff _57088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _03216_, clk);
  dff _57089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _15234_, clk);
  dff _57090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _15162_, clk);
  dff _57091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _03907_, clk);
  dff _57092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _27034_, clk);
  dff _57093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _27035_, clk);
  dff _57094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _03827_, clk);
  dff _57095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _22636_, clk);
  dff _57096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _03064_, clk);
  dff _57097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _27030_, clk);
  dff _57098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _27031_, clk);
  dff _57099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _22617_, clk);
  dff _57100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _27032_, clk);
  dff _57101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _19201_, clk);
  dff _57102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _03804_, clk);
  dff _57103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _22646_, clk);
  dff _57104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _27028_, clk);
  dff _57105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _27029_, clk);
  dff _57106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _22654_, clk);
  dff _57107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _22650_, clk);
  dff _57108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _03812_, clk);
  dff _57109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _22626_, clk);
  dff _57110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _05238_, clk);
  dff _57111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _03069_, clk);
  dff _57112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _05474_, clk);
  dff _57113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _05714_, clk);
  dff _57114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _03076_, clk);
  dff _57115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _27022_, clk);
  dff _57116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _05222_, clk);
  dff _57117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _03112_, clk);
  dff _57118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _03092_, clk);
  dff _57119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _27025_, clk);
  dff _57120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _22675_, clk);
  dff _57121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _27026_, clk);
  dff _57122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _22713_, clk);
  dff _57123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _27027_, clk);
  dff _57124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _22656_, clk);
  dff _57125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _22660_, clk);
  dff _57126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _27016_, clk);
  dff _57127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _02853_, clk);
  dff _57128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _02878_, clk);
  dff _57129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _27017_, clk);
  dff _57130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _05644_, clk);
  dff _57131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _27018_, clk);
  dff _57132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _05272_, clk);
  dff _57133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _02933_, clk);
  dff _57134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _03000_, clk);
  dff _57135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _05252_, clk);
  dff _57136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _03012_, clk);
  dff _57137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _05503_, clk);
  dff _57138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _03027_, clk);
  dff _57139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _05245_, clk);
  dff _57140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _03047_, clk);
  dff _57141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _05483_, clk);
  dff _57142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _01604_, clk);
  dff _57143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _27014_, clk);
  dff _57144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _01606_, clk);
  dff _57145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _27015_, clk);
  dff _57146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _05283_, clk);
  dff _57147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _05650_, clk);
  dff _57148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _02822_, clk);
  dff _57149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _02850_, clk);
  dff _57150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _00299_, clk);
  dff _57151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _05336_, clk);
  dff _57152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _00305_, clk);
  dff _57153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _05557_, clk);
  dff _57154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _00310_, clk);
  dff _57155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _00596_, clk);
  dff _57156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _05325_, clk);
  dff _57157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _01600_, clk);
  dff _57158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _27013_, clk);
  dff _57159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _00270_, clk);
  dff _57160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _05354_, clk);
  dff _57161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _00276_, clk);
  dff _57162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _05564_, clk);
  dff _57163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _00280_, clk);
  dff _57164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _00291_, clk);
  dff _57165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _05346_, clk);
  dff _57166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _05581_, clk);
  dff _57167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _00203_, clk);
  dff _57168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _05369_, clk);
  dff _57169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _00209_, clk);
  dff _57170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _05575_, clk);
  dff _57171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _00212_, clk);
  dff _57172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _00262_, clk);
  dff _57173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _05357_, clk);
  dff _57174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _05729_, clk);
  dff _57175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _25996_, clk);
  dff _57176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _26012_, clk);
  dff _57177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _05452_, clk);
  dff _57178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _26015_, clk);
  dff _57179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _26019_, clk);
  dff _57180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _05447_, clk);
  dff _57181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _05695_, clk);
  dff _57182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _27012_, clk);
  dff _57183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _05588_, clk);
  dff _57184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _26086_, clk);
  dff _57185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _05390_, clk);
  dff _57186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _26096_, clk);
  dff _57187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _05586_, clk);
  dff _57188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _26117_, clk);
  dff _57189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _00103_, clk);
  dff _57190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _03422_, clk);
  dff _57191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _03415_, clk);
  dff _57192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _06558_, clk);
  dff _57193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _03480_, clk);
  dff _57194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _03472_, clk);
  dff _57195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _05778_, clk);
  dff _57196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _27005_, clk);
  dff _57197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _27006_, clk);
  dff _57198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _05433_, clk);
  dff _57199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _27010_, clk);
  dff _57200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _27011_, clk);
  dff _57201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _26056_, clk);
  dff _57202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _05423_, clk);
  dff _57203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _26062_, clk);
  dff _57204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _05590_, clk);
  dff _57205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _26069_, clk);
  dff _57206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _03342_, clk);
  dff _57207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _03321_, clk);
  dff _57208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _25946_, clk);
  dff _57209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _25939_, clk);
  dff _57210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _06569_, clk);
  dff _57211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _03223_, clk);
  dff _57212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _03206_, clk);
  dff _57213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _06564_, clk);
  dff _57214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _03820_, clk);
  dff _57215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _05781_, clk);
  dff _57216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _03553_, clk);
  dff _57217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _27002_, clk);
  dff _57218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _03631_, clk);
  dff _57219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _27003_, clk);
  dff _57220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _27004_, clk);
  dff _57221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _03440_, clk);
  dff _57222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _04013_, clk);
  dff _57223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _27001_, clk);
  dff _57224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _03974_, clk);
  dff _57225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _05786_, clk);
  dff _57226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _03659_, clk);
  dff _57227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _03716_, clk);
  dff _57228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _03697_, clk);
  dff _57229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _03836_, clk);
  dff _57230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _04055_, clk);
  dff _57231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _04185_, clk);
  dff _57232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _04165_, clk);
  dff _57233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _04159_, clk);
  dff _57234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _06530_, clk);
  dff _57235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _27000_, clk);
  dff _57236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _03867_, clk);
  dff _57237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _03900_, clk);
  dff _57238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _04279_, clk);
  dff _57239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _04273_, clk);
  dff _57240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _26998_, clk);
  dff _57241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _26999_, clk);
  dff _57242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _04386_, clk);
  dff _57243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _06519_, clk);
  dff _57244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _04109_, clk);
  dff _57245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _04092_, clk);
  dff _57246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _07117_, clk);
  dff _57247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _07083_, clk);
  dff _57248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _01698_, clk);
  dff _57249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _27178_, clk);
  dff _57250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _01688_, clk);
  dff _57251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _06928_, clk);
  dff _57252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _06897_, clk);
  dff _57253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _01729_, clk);
  dff _57254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _26995_, clk);
  dff _57255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _04492_, clk);
  dff _57256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _04471_, clk);
  dff _57257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _26996_, clk);
  dff _57258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _04576_, clk);
  dff _57259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _04571_, clk);
  dff _57260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _26997_, clk);
  dff _57261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _06147_, clk);
  dff _57262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _06485_, clk);
  dff _57263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _26993_, clk);
  dff _57264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _26994_, clk);
  dff _57265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _04679_, clk);
  dff _57266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _04664_, clk);
  dff _57267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _04734_, clk);
  dff _57268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _04765_, clk);
  dff _57269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _04740_, clk);
  dff _57270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _05166_, clk);
  dff _57271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _06477_, clk);
  dff _57272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _05241_, clk);
  dff _57273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _05220_, clk);
  dff _57274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _05812_, clk);
  dff _57275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _06149_, clk);
  dff _57276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _26988_, clk);
  dff _57277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04966_, clk);
  dff _57278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _26989_, clk);
  dff _57279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _26990_, clk);
  dff _57280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _26991_, clk);
  dff _57281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _04817_, clk);
  dff _57282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _04845_, clk);
  dff _57283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _26992_, clk);
  dff _57284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _04927_, clk);
  dff _57285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _04917_, clk);
  dff _57286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _05740_, clk);
  dff _57287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _05718_, clk);
  dff _57288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _05320_, clk);
  dff _57289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _26987_, clk);
  dff _57290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _05794_, clk);
  dff _57291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _05788_, clk);
  dff _57292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _06467_, clk);
  dff _57293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _05172_, clk);
  dff _57294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _06457_, clk);
  dff _57295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _06059_, clk);
  dff _57296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _05820_, clk);
  dff _57297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _05840_, clk);
  dff _57298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _05833_, clk);
  dff _57299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _06462_, clk);
  dff _57300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _05928_, clk);
  dff _57301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _06459_, clk);
  dff _57302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _06123_, clk);
  dff _57303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _06107_, clk);
  dff _57304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _26984_, clk);
  dff _57305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _26985_, clk);
  dff _57306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _05825_, clk);
  dff _57307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _06151_, clk);
  dff _57308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _06021_, clk);
  dff _57309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _05998_, clk);
  dff _57310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _06434_, clk);
  dff _57311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _06380_, clk);
  dff _57312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _06408_, clk);
  dff _57313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _06396_, clk);
  dff _57314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _06444_, clk);
  dff _57315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _26982_, clk);
  dff _57316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _06465_, clk);
  dff _57317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _06439_, clk);
  dff _57318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _06280_, clk);
  dff _57319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _06266_, clk);
  dff _57320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _06248_, clk);
  dff _57321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _26983_, clk);
  dff _57322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _06333_, clk);
  dff _57323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _06327_, clk);
  dff _57324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _06314_, clk);
  dff _57325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _06445_, clk);
  dff _57326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _06428_, clk);
  dff _57327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _06068_, clk);
  dff _57328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _26980_, clk);
  dff _57329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _06547_, clk);
  dff _57330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _06541_, clk);
  dff _57331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _06436_, clk);
  dff _57332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _26981_, clk);
  dff _57333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _06627_, clk);
  dff _57334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _06886_, clk);
  dff _57335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _06881_, clk);
  dff _57336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _06420_, clk);
  dff _57337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _06667_, clk);
  dff _57338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _06707_, clk);
  dff _57339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _06744_, clk);
  dff _57340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _06760_, clk);
  dff _57341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _26979_, clk);
  dff _57342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _07010_, clk);
  dff _57343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _07049_, clk);
  dff _57344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _07039_, clk);
  dff _57345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _26976_, clk);
  dff _57346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _26977_, clk);
  dff _57347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _06823_, clk);
  dff _57348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _06817_, clk);
  dff _57349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _26978_, clk);
  dff _57350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _06401_, clk);
  dff _57351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _07270_, clk);
  dff _57352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _07266_, clk);
  dff _57353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _07251_, clk);
  dff _57354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _07349_, clk);
  dff _57355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _07341_, clk);
  dff _57356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _26974_, clk);
  dff _57357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _05859_, clk);
  dff _57358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _07125_, clk);
  dff _57359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _07115_, clk);
  dff _57360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _07089_, clk);
  dff _57361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _07204_, clk);
  dff _57362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _07185_, clk);
  dff _57363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _26975_, clk);
  dff _57364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _06964_, clk);
  dff _57365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _06960_, clk);
  dff _57366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _07607_, clk);
  dff _57367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _07586_, clk);
  dff _57368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _05866_, clk);
  dff _57369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _26973_, clk);
  dff _57370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _07407_, clk);
  dff _57371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _07394_, clk);
  dff _57372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _06403_, clk);
  dff _57373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _07471_, clk);
  dff _57374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _06169_, clk);
  dff _57375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _07648_, clk);
  dff _57376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _26969_, clk);
  dff _57377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _07908_, clk);
  dff _57378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _07902_, clk);
  dff _57379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _06390_, clk);
  dff _57380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07542_, clk);
  dff _57381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _07528_, clk);
  dff _57382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _09056_, clk);
  dff _57383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _09002_, clk);
  dff _57384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _05909_, clk);
  dff _57385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _08253_, clk);
  dff _57386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _08249_, clk);
  dff _57387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _08280_, clk);
  dff _57388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _08278_, clk);
  dff _57389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _06373_, clk);
  dff _57390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _06225_, clk);
  dff _57391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _06214_, clk);
  dff _57392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _26966_, clk);
  dff _57393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _26967_, clk);
  dff _57394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _10003_, clk);
  dff _57395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _10050_, clk);
  dff _57396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _26968_, clk);
  dff _57397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _05913_, clk);
  dff _57398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _09122_, clk);
  dff _57399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _09069_, clk);
  dff _57400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _09788_, clk);
  dff _57401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _09232_, clk);
  dff _57402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _09228_, clk);
  dff _57403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _06355_, clk);
  dff _57404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _08905_, clk);
  dff _57405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _08862_, clk);
  dff _57406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _01388_, clk);
  dff _57407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _26963_, clk);
  dff _57408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _04126_, clk);
  dff _57409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _26964_, clk);
  dff _57410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _26965_, clk);
  dff _57411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _00184_, clk);
  dff _57412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _25957_, clk);
  dff _57413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _02533_, clk);
  dff _57414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _26962_, clk);
  dff _57415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _06229_, clk);
  dff _57416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _10970_, clk);
  dff _57417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _11914_, clk);
  dff _57418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _06232_, clk);
  dff _57419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _06120_, clk);
  dff _57420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _06243_, clk);
  dff _57421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _10653_, clk);
  dff _57422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _26953_, clk);
  dff _57423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _26954_, clk);
  dff _57424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _26955_, clk);
  dff _57425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _11162_, clk);
  dff _57426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _11142_, clk);
  dff _57427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _11262_, clk);
  dff _57428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _11249_, clk);
  dff _57429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _26956_, clk);
  dff _57430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _11795_, clk);
  dff _57431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _11909_, clk);
  dff _57432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _05945_, clk);
  dff _57433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _11512_, clk);
  dff _57434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _06309_, clk);
  dff _57435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _11641_, clk);
  dff _57436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _26950_, clk);
  dff _57437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _11357_, clk);
  dff _57438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _12369_, clk);
  dff _57439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _12344_, clk);
  dff _57440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _05951_, clk);
  dff _57441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _11932_, clk);
  dff _57442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _26949_, clk);
  dff _57443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _12224_, clk);
  dff _57444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _06297_, clk);
  dff _57445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _06095_, clk);
  dff _57446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _11627_, clk);
  dff _57447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _06285_, clk);
  dff _57448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _26948_, clk);
  dff _57449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _06288_, clk);
  dff _57450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _10420_, clk);
  dff _57451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _05974_, clk);
  dff _57452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _10921_, clk);
  dff _57453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _10694_, clk);
  dff _57454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _08780_, clk);
  dff _57455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _24419_, clk);
  dff _57456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _05960_, clk);
  dff _57457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _12404_, clk);
  dff _57458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _24475_, clk);
  dff _57459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _05676_, clk);
  dff _57460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _05954_, clk);
  dff _57461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _12301_, clk);
  dff _57462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _05892_, clk);
  dff _57463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _06275_, clk);
  dff _57464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _05981_, clk);
  dff _57465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _11654_, clk);
  dff _57466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _06282_, clk);
  dff _57467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _06277_, clk);
  dff _57468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _26947_, clk);
  dff _57469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _11074_, clk);
  dff _57470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _26942_, clk);
  dff _57471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _26943_, clk);
  dff _57472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _06983_, clk);
  dff _57473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _26944_, clk);
  dff _57474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _06978_, clk);
  dff _57475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _26945_, clk);
  dff _57476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _26946_, clk);
  dff _57477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _10826_, clk);
  dff _57478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _07317_, clk);
  dff _57479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _10639_, clk);
  dff _57480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _07033_, clk);
  dff _57481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _26936_, clk);
  dff _57482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _07194_, clk);
  dff _57483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _10648_, clk);
  dff _57484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _10692_, clk);
  dff _57485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _26937_, clk);
  dff _57486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _10723_, clk);
  dff _57487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _10734_, clk);
  dff _57488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _26938_, clk);
  dff _57489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _07003_, clk);
  dff _57490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _26939_, clk);
  dff _57491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _07188_, clk);
  dff _57492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _26940_, clk);
  dff _57493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _26941_, clk);
  dff _57494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _09119_, clk);
  dff _57495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _07061_, clk);
  dff _57496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _09157_, clk);
  dff _57497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _07059_, clk);
  dff _57498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _09196_, clk);
  dff _57499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _07201_, clk);
  dff _57500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _09201_, clk);
  dff _57501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _09755_, clk);
  dff _57502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _07216_, clk);
  dff _57503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _07959_, clk);
  dff _57504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _08259_, clk);
  dff _57505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _07075_, clk);
  dff _57506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _07297_, clk);
  dff _57507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _08284_, clk);
  dff _57508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _08912_, clk);
  dff _57509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _26931_, clk);
  dff _57510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _07081_, clk);
  dff _57511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _07300_, clk);
  dff _57512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _05175_, clk);
  dff _57513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _26926_, clk);
  dff _57514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _07164_, clk);
  dff _57515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _05163_, clk);
  dff _57516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _26927_, clk);
  dff _57517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _05379_, clk);
  dff _57518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _26928_, clk);
  dff _57519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _26929_, clk);
  dff _57520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _26930_, clk);
  dff _57521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _05978_, clk);
  dff _57522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _07245_, clk);
  dff _57523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _07324_, clk);
  dff _57524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _07535_, clk);
  dff _57525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _07952_, clk);
  dff _57526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _07221_, clk);
  dff _57527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _07293_, clk);
  dff _57528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _07232_, clk);
  dff _57529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _07418_, clk);
  dff _57530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _07456_, clk);
  dff _57531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _07094_, clk);
  dff _57532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _07469_, clk);
  dff _57533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _07092_, clk);
  dff _57534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _07113_, clk);
  dff _57535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _07051_, clk);
  dff _57536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _26924_, clk);
  dff _57537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _07054_, clk);
  dff _57538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _26925_, clk);
  dff _57539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _07145_, clk);
  dff _57540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _07107_, clk);
  dff _57541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _07177_, clk);
  dff _57542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _06045_, clk);
  dff _57543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _07141_, clk);
  dff _57544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06054_, clk);
  dff _57545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _06065_, clk);
  dff _57546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _06414_, clk);
  dff _57547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _07130_, clk);
  dff _57548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _07309_, clk);
  dff _57549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _06416_, clk);
  dff _57550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _26918_, clk);
  dff _57551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _09057_, clk);
  dff _57552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _26919_, clk);
  dff _57553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _26920_, clk);
  dff _57554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _08887_, clk);
  dff _57555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _09139_, clk);
  dff _57556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _11042_, clk);
  dff _57557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _11050_, clk);
  dff _57558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _26911_, clk);
  dff _57559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _08896_, clk);
  dff _57560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _26912_, clk);
  dff _57561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _26913_, clk);
  dff _57562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _26914_, clk);
  dff _57563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _26915_, clk);
  dff _57564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _08892_, clk);
  dff _57565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _26916_, clk);
  dff _57566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _10645_, clk);
  dff _57567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _26906_, clk);
  dff _57568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _26907_, clk);
  dff _57569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _26908_, clk);
  dff _57570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _10696_, clk);
  dff _57571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _26909_, clk);
  dff _57572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _10747_, clk);
  dff _57573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _26910_, clk);
  dff _57574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _10093_, clk);
  dff _57575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _10113_, clk);
  dff _57576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _26897_, clk);
  dff _57577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _10144_, clk);
  dff _57578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _08995_, clk);
  dff _57579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _09216_, clk);
  dff _57580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _26898_, clk);
  dff _57581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _09209_, clk);
  dff _57582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _27218_, clk);
  dff _57583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _10853_, clk);
  dff _57584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _11170_, clk);
  dff _57585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _11305_, clk);
  dff _57586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _11197_, clk);
  dff _57587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _09977_, clk);
  dff _57588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _09664_, clk);
  dff _57589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _09630_, clk);
  dff _57590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _09108_, clk);
  dff _57591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _10572_, clk);
  dff _57592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _10601_, clk);
  dff _57593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _08925_, clk);
  dff _57594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _09177_, clk);
  dff _57595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _10618_, clk);
  dff _57596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _08923_, clk);
  dff _57597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _10624_, clk);
  dff _57598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _10018_, clk);
  dff _57599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _09034_, clk);
  dff _57600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _09188_, clk);
  dff _57601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _10045_, clk);
  dff _57602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _09009_, clk);
  dff _57603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _10055_, clk);
  dff _57604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _26896_, clk);
  dff _57605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _08999_, clk);
  dff _57606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _26895_, clk);
  dff _57607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _09939_, clk);
  dff _57608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _09953_, clk);
  dff _57609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _09042_, clk);
  dff _57610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _09961_, clk);
  dff _57611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _09972_, clk);
  dff _57612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _09038_, clk);
  dff _57613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _10006_, clk);
  dff _57614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _11068_, clk);
  dff _57615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _04666_, clk);
  dff _57616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _04746_, clk);
  dff _57617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _04805_, clk);
  dff _57618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _04717_, clk);
  dff _57619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _04460_, clk);
  dff _57620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _27313_[6], clk);
  dff _57621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _12348_, clk);
  dff _57622_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _57623_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _57624_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _57625_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _57626_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _57627_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _57628_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _57629_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _57630_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _57631_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _57632_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _57633_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _57634_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _57635_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _57636_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _57637_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _57638_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _57639_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _57640_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _57641_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _57642_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _57643_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _57644_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _57645_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _57646_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _57647_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _57648_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _57649_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _57650_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _57651_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _57652_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _57653_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _57654_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _27314_, clk);
  dff _57655_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _27315_[0], clk);
  dff _57656_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _27315_[1], clk);
  dff _57657_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _27315_[2], clk);
  dff _57658_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _27315_[3], clk);
  dff _57659_ (\oc8051_top_1.oc8051_sfr1.bit_out , _27316_, clk);
  dff _57660_ (\oc8051_top_1.oc8051_sfr1.wait_data , _27317_, clk);
  dff _57661_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _27318_[0], clk);
  dff _57662_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _27318_[1], clk);
  dff _57663_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _27318_[2], clk);
  dff _57664_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _27318_[3], clk);
  dff _57665_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _27318_[4], clk);
  dff _57666_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _27318_[5], clk);
  dff _57667_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _27318_[6], clk);
  dff _57668_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _27318_[7], clk);
  dff _57669_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10454_, clk);
  dff _57670_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10442_, clk);
  dff _57671_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10266_, clk);
  dff _57672_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10304_, clk);
  dff _57673_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10358_, clk);
  dff _57674_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10324_, clk);
  dff _57675_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10220_, clk);
  dff _57676_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10147_, clk);
  dff _57677_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _06501_, clk);
  dff _57678_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _06506_, clk);
  dff _57679_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _06504_, clk);
  dff _57680_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _06511_, clk);
  dff _57681_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _06517_, clk);
  dff _57682_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _06514_, clk);
  dff _57683_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _06526_, clk);
  dff _57684_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05463_, clk);
  dff _57685_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _09920_, clk);
  dff _57686_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _09918_, clk);
  dff _57687_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _09881_, clk);
  dff _57688_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _09875_, clk);
  dff _57689_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _09864_, clk);
  dff _57690_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _09741_, clk);
  dff _57691_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _09959_, clk);
  dff _57692_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _09766_, clk);
  dff _57693_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09776_, clk);
  dff _57694_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _09911_, clk);
  dff _57695_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _09837_, clk);
  dff _57696_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _09800_, clk);
  dff _57697_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _09916_, clk);
  dff _57698_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _09914_, clk);
  dff _57699_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _09835_, clk);
  dff _57700_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _09929_, clk);
  dff _57701_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _11411_, clk);
  dff _57702_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _22640_, clk);
  dff _57703_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _09539_, clk);
  dff _57704_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _09650_, clk);
  dff _57705_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _09621_, clk);
  dff _57706_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _09580_, clk);
  dff _57707_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _09560_, clk);
  dff _57708_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22639_, clk);
  dff _57709_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _11486_, clk);
  dff _57710_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _08845_, clk);
  dff _57711_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _11258_, clk);
  dff _57712_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _11366_, clk);
  dff _57713_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _08746_, clk);
  dff _57714_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _22642_, clk);
  dff _57715_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _11334_, clk);
  dff _57716_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _09118_, clk);
  dff _57717_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _22641_, clk);
  dff _57718_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _11328_, clk);
  dff _57719_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _08233_, clk);
  dff _57720_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08572_, clk);
  dff _57721_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _11352_, clk);
  dff _57722_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _11268_, clk);
  dff _57723_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _11347_, clk);
  dff _57724_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _11310_, clk);
  dff _57725_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _07742_, clk);
  dff _57726_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _07723_, clk);
  dff _57727_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _07703_, clk);
  dff _57728_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _11322_, clk);
  dff _57729_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _07156_, clk);
  dff _57730_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _06967_, clk);
  dff _57731_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _07135_, clk);
  dff _57732_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _07072_, clk);
  dff _57733_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _07024_, clk);
  dff _57734_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _22643_, clk);
  dff _57735_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _07479_, clk);
  dff _57736_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _11372_, clk);
  dff _57737_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _06560_, clk);
  dff _57738_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _06536_, clk);
  dff _57739_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _06510_, clk);
  dff _57740_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _06442_, clk);
  dff _57741_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _22644_, clk);
  dff _57742_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _06793_, clk);
  dff _57743_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _06752_, clk);
  dff _57744_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _11355_, clk);
  dff _57745_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _11669_, clk);
  dff _57746_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _11644_, clk);
  dff _57747_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _11618_, clk);
  dff _57748_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _05791_, clk);
  dff _57749_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _11994_, clk);
  dff _57750_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _11891_, clk);
  dff _57751_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _11973_, clk);
  dff _57752_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _10870_, clk);
  dff _57753_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _11035_, clk);
  dff _57754_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _10987_, clk);
  dff _57755_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _10960_, clk);
  dff _57756_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _10934_, clk);
  dff _57757_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _05805_, clk);
  dff _57758_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _11356_, clk);
  dff _57759_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _11255_, clk);
  dff _57760_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _10857_, clk);
  dff _57761_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _10592_, clk);
  dff _57762_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _10460_, clk);
  dff _57763_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _10565_, clk);
  dff _57764_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _10541_, clk);
  dff _57765_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _10516_, clk);
  dff _57766_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _10482_, clk);
  dff _57767_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _05816_, clk);
  dff _57768_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _10753_, clk);
  dff _57769_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _09922_, clk);
  dff _57770_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _09894_, clk);
  dff _57771_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _09868_, clk);
  dff _57772_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _09786_, clk);
  dff _57773_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _05843_, clk);
  dff _57774_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _10293_, clk);
  dff _57775_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _10136_, clk);
  dff _57776_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _10842_, clk);
  dff _57777_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10161_, clk);
  dff _57778_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10130_, clk);
  dff _57779_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10118_, clk);
  dff _57780_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10102_, clk);
  dff _57781_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10120_, clk);
  dff _57782_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10132_, clk);
  dff _57783_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _09826_, clk);
  dff _57784_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _06681_, clk);
  dff _57785_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _06980_, clk);
  dff _57786_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _06974_, clk);
  dff _57787_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _06992_, clk);
  dff _57788_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _06988_, clk);
  dff _57789_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _06990_, clk);
  dff _57790_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _06999_, clk);
  dff _57791_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _06997_, clk);
  dff _57792_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _06701_, clk);
  dff _57793_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _22716_, clk);
  dff _57794_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _03359_, clk);
  dff _57795_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _04010_, clk);
  dff _57796_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _05666_, clk);
  dff _57797_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _05602_, clk);
  dff _57798_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _04002_, clk);
  dff _57799_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _01093_, clk);
  dff _57800_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _11027_, clk);
  dff _57801_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _10620_, clk);
  dff _57802_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _22697_, clk);
  dff _57803_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _04015_, clk);
  dff _57804_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _05476_, clk);
  dff _57805_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _05019_, clk);
  dff _57806_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _09955_, clk);
  dff _57807_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _08662_, clk);
  dff _57808_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _06161_, clk);
  dff _57809_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _22670_, clk);
  dff _57810_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _09079_, clk);
  dff _57811_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _22652_, clk);
  dff _57812_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _09462_, clk);
  dff _57813_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12417_, clk);
  dff _57814_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12413_, clk);
  dff _57815_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12412_, clk);
  dff _57816_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _04044_, clk);
  dff _57817_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12432_, clk);
  dff _57818_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _07109_, clk);
  dff _57819_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _02667_, clk);
  dff _57820_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _22649_, clk);
  dff _57821_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12355_, clk);
  dff _57822_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12351_, clk);
  dff _57823_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _04046_, clk);
  dff _57824_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _12391_, clk);
  dff _57825_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _12390_, clk);
  dff _57826_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _12387_, clk);
  dff _57827_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _12384_, clk);
  dff _57828_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _22653_, clk);
  dff _57829_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _22624_, clk);
  dff _57830_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12325_, clk);
  dff _57831_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12316_, clk);
  dff _57832_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _04077_, clk);
  dff _57833_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _05477_, clk);
  dff _57834_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _26179_, clk);
  dff _57835_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _09136_, clk);
  dff _57836_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _24427_, clk);
  dff _57837_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _02924_, clk);
  dff _57838_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _18134_, clk);
  dff _57839_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _18119_, clk);
  dff _57840_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _18105_, clk);
  dff _57841_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _17956_, clk);
  dff _57842_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _08907_, clk);
  dff _57843_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02719_, clk);
  dff _57844_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _07409_, clk);
  dff _57845_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _08711_, clk);
  dff _57846_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _08701_, clk);
  dff _57847_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _08288_, clk);
  dff _57848_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02751_, clk);
  dff _57849_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _17942_, clk);
  dff _57850_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02766_, clk);
  dff _57851_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _08270_, clk);
  dff _57852_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _08268_, clk);
  dff _57853_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _08266_, clk);
  dff _57854_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02763_, clk);
  dff _57855_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _08242_, clk);
  dff _57856_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _08237_, clk);
  dff _57857_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _17922_, clk);
  dff _57858_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _17853_, clk);
  dff _57859_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _07896_, clk);
  dff _57860_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _07891_, clk);
  dff _57861_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _07889_, clk);
  dff _57862_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02788_, clk);
  dff _57863_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _07917_, clk);
  dff _57864_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _07905_, clk);
  dff _57865_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _07914_, clk);
  dff _57866_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _17818_, clk);
  dff _57867_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _07875_, clk);
  dff _57868_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _07884_, clk);
  dff _57869_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _07881_, clk);
  dff _57870_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _07879_, clk);
  dff _57871_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _07877_, clk);
  dff _57872_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02791_, clk);
  dff _57873_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _07624_, clk);
  dff _57874_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _17768_, clk);
  dff _57875_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _17752_, clk);
  dff _57876_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _07639_, clk);
  dff _57877_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02805_, clk);
  dff _57878_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _07577_, clk);
  dff _57879_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _07562_, clk);
  dff _57880_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _07558_, clk);
  dff _57881_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02843_, clk);
  dff _57882_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _07603_, clk);
  dff _57883_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _17618_, clk);
  dff _57884_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _22883_, clk);
  dff _57885_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _22895_, clk);
  dff _57886_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _22892_, clk);
  dff _57887_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _22889_, clk);
  dff _57888_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _22722_, clk);
  dff _57889_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _22765_, clk);
  dff _57890_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _22715_, clk);
  dff _57891_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _22718_, clk);
  dff _57892_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _22719_, clk);
  dff _57893_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _22725_, clk);
  dff _57894_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22727_, clk);
  dff _57895_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01368_, clk);
  dff _57896_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _01336_, clk);
  dff _57897_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _25690_, clk);
  dff _57898_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _25688_, clk);
  dff _57899_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _01421_, clk);
  dff _57900_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _25708_, clk);
  dff _57901_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _25706_, clk);
  dff _57902_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _22748_, clk);
  dff _57903_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _01409_, clk);
  dff _57904_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _22726_, clk);
  dff _57905_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _22728_, clk);
  dff _57906_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _22807_, clk);
  dff _57907_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _01334_, clk);
  dff _57908_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _22632_, clk);
  dff _57909_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _22633_, clk);
  dff _57910_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _22842_, clk);
  dff _57911_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _22631_, clk);
  dff _57912_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _22870_, clk);
  dff _57913_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _22819_, clk);
  dff _57914_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _22848_, clk);
  dff _57915_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _01355_, clk);
  dff _57916_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _25655_, clk);
  dff _57917_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _25638_, clk);
  dff _57918_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _25646_, clk);
  dff _57919_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _01426_, clk);
  dff _57920_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _22730_, clk);
  dff _57921_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _22754_, clk);
  dff _57922_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _22756_, clk);
  dff _57923_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _25680_, clk);
  dff _57924_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _22712_, clk);
  dff _57925_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _22711_, clk);
  dff _57926_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _22710_, clk);
  dff _57927_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _22709_, clk);
  dff _57928_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _22708_, clk);
  dff _57929_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _22707_, clk);
  dff _57930_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _22706_, clk);
  dff _57931_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _22705_, clk);
  dff _57932_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22704_, clk);
  dff _57933_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22703_, clk);
  dff _57934_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _25678_, clk);
  dff _57935_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _22702_, clk);
  dff _57936_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _22701_, clk);
  dff _57937_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _22629_, clk);
  dff _57938_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _22700_, clk);
  dff _57939_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _26109_, clk);
  dff _57940_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _22699_, clk);
  dff _57941_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _22698_, clk);
  dff _57942_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01423_, clk);
  dff _57943_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _22696_, clk);
  dff _57944_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _22695_, clk);
  dff _57945_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _22694_, clk);
  dff _57946_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _22693_, clk);
  dff _57947_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _22692_, clk);
  dff _57948_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _22691_, clk);
  dff _57949_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _22690_, clk);
  dff _57950_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01332_, clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
